library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package angrypkg is
    type angry2D is array(0 to 23, 0 to 25) of integer range 0 to 9;
end package;

use work.angrypkg.all;

entity angryBird is
      Port (bird: out angry2D );
end angryBird;

architecture Behavioral of angryBird is

begin

bird(0, 0) <= 0; bird(0, 1) <= 0; bird(0, 2) <= 0; bird(0, 3) <= 0; bird(0, 4) <= 0; bird(0, 5) <= 0; bird(0, 6) <= 0; bird(0, 7) <= 0; bird(0, 8) <= 0; bird(0, 9) <= 0; bird(0, 10) <= 0; bird(0, 11) <= 0; bird(0, 12) <= 5; bird(0, 13) <= 5; bird(0, 14) <= 5; bird(0, 15) <= 0; bird(0, 16) <= 0; bird(0, 17) <= 0; bird(0, 18) <= 0; bird(0, 19) <= 0; bird(0, 20) <= 0; bird(0, 21) <= 0; bird(0, 22) <= 0; bird(0, 23) <= 0; bird(0, 24) <= 0; bird(1, 0) <= 0; 
bird(1, 1) <= 0; bird(1, 2) <= 0; bird(1, 3) <= 0; bird(1, 4) <= 0; bird(1, 5) <= 0; bird(1, 6) <= 0; bird(1, 7) <= 0; 
bird(1, 8) <= 0; bird(1, 9) <= 0; bird(1, 10) <= 0; bird(1, 11) <= 5; bird(1, 12) <= 4; bird(1, 13) <= 4; bird(1, 14) <= 4; 
bird(1, 15) <= 5; bird(1, 16) <= 0; bird(1, 17) <= 0; bird(1, 18) <= 0; bird(1, 19) <= 0; bird(1, 20) <= 0; bird(1, 21) <= 0; 
bird(1, 22) <= 0; bird(1, 23) <= 0; bird(1, 24) <= 0; bird(2, 0) <= 0; 
bird(2, 1) <= 0; bird(2, 2) <= 0; bird(2, 3) <= 0; bird(2, 4) <= 0; bird(2, 5) <= 0; bird(2, 6) <= 0; bird(2, 7) <= 0; 
bird(2, 8) <= 5; bird(2, 9) <= 5; bird(2, 10) <= 5; bird(2, 11) <= 5; bird(2, 12) <= 4; bird(2, 13) <= 4; bird(2, 14) <= 4; 
bird(2, 15) <= 4; bird(2, 16) <= 5; bird(2, 17) <= 0; bird(2, 18) <= 0; bird(2, 19) <= 0; bird(2, 20) <= 0; bird(2, 21) <= 0; 
bird(2, 22) <= 0; bird(2, 23) <= 0; bird(2, 24) <= 0; bird(3, 0) <= 0; 
bird(3, 1) <= 0; bird(3, 2) <= 0; bird(3, 3) <= 0; bird(3, 4) <= 0; bird(3, 5) <= 0; bird(3, 6) <= 0; bird(3, 7) <= 5; 
bird(3, 8) <= 4; bird(3, 9) <= 4; bird(3, 10) <= 4; bird(3, 11) <= 4; bird(3, 12) <= 4; bird(3, 13) <= 4; bird(3, 14) <= 4; 
bird(3, 15) <= 4; bird(3, 16) <= 4; bird(3, 17) <= 5; bird(3, 18) <= 0; bird(3, 19) <= 0; bird(3, 20) <= 0; bird(3, 21) <= 0; 
bird(3, 22) <= 0; bird(3, 23) <= 0; bird(3, 24) <= 0; bird(4, 0) <= 0; 
bird(4, 1) <= 0; bird(4, 2) <= 0; bird(4, 3) <= 0; bird(4, 4) <= 0; bird(4, 5) <= 0; bird(4, 6) <= 0; bird(4, 7) <= 5; 
bird(4, 8) <= 4; bird(4, 9) <= 4; bird(4, 10) <= 4; bird(4, 11) <= 4; bird(4, 12) <= 4; bird(4, 13) <= 4; bird(4, 14) <= 4; 
bird(4, 15) <= 4; bird(4, 16) <= 4; bird(4, 17) <= 4; bird(4, 18) <= 5; bird(4, 19) <= 0; bird(4, 20) <= 0; bird(4, 21) <= 0; 
bird(4, 22) <= 0; bird(4, 23) <= 0; bird(4, 24) <= 0; bird(5, 0) <= 0; 
bird(5, 1) <= 0; bird(5, 2) <= 0; bird(5, 3) <= 0; bird(5, 4) <= 0; bird(5, 5) <= 0; bird(5, 6) <= 0; bird(5, 7) <= 0; 
bird(5, 8) <= 5; bird(5, 9) <= 5; bird(5, 10) <= 5; bird(5, 11) <= 4; bird(5, 12) <= 4; bird(5, 13) <= 4; bird(5, 14) <= 4; 
bird(5, 15) <= 4; bird(5, 16) <= 4; bird(5, 17) <= 4; bird(5, 18) <= 4; bird(5, 19) <= 5; bird(5, 20) <= 0; bird(5, 21) <= 0; 
bird(5, 22) <= 0; bird(5, 23) <= 0; bird(5, 24) <= 0; bird(6, 0) <= 0; 
bird(6, 1) <= 0; bird(6, 2) <= 0; bird(6, 3) <= 0; bird(6, 4) <= 0; bird(6, 5) <= 0; bird(6, 6) <= 0; bird(6, 7) <= 5; 
bird(6, 8) <= 4; bird(6, 9) <= 4; bird(6, 10) <= 4; bird(6, 11) <= 4; bird(6, 12) <= 4; bird(6, 13) <= 4; bird(6, 14) <= 4; 
bird(6, 15) <= 4; bird(6, 16) <= 4; bird(6, 17) <= 4; bird(6, 18) <= 4; bird(6, 19) <= 4; bird(6, 20) <= 5; bird(6, 21) <= 0; 
bird(6, 22) <= 0; bird(6, 23) <= 0; bird(6, 24) <= 0; bird(7, 0) <= 0; 
bird(7, 1) <= 0; bird(7, 2) <= 0; bird(7, 3) <= 0; bird(7, 4) <= 0; bird(7, 5) <= 0; bird(7, 6) <= 5; bird(7, 7) <= 4; 
bird(7, 8) <= 4; bird(7, 9) <= 4; bird(7, 10) <= 4; bird(7, 11) <= 4; bird(7, 12) <= 4; bird(7, 13) <= 4; bird(7, 14) <= 4; 
bird(7, 15) <= 4; bird(7, 16) <= 4; bird(7, 17) <= 4; bird(7, 18) <= 4; bird(7, 19) <= 4; bird(7, 20) <= 4; bird(7, 21) <= 5; 
bird(7, 22) <= 0; bird(7, 23) <= 0; bird(7, 24) <= 0; bird(8, 0) <= 0; 
bird(8, 1) <= 0; bird(8, 2) <= 0; bird(8, 3) <= 0; bird(8, 4) <= 0; bird(8, 5) <= 0; bird(8, 6) <= 5; bird(8, 7) <= 4; 
bird(8, 8) <= 4; bird(8, 9) <= 4; bird(8, 10) <= 4; bird(8, 11) <= 4; bird(8, 12) <= 4; bird(8, 13) <= 4; bird(8, 14) <= 4; 
bird(8, 15) <= 4; bird(8, 16) <= 4; bird(8, 17) <= 4; bird(8, 18) <= 4; bird(8, 19) <= 4; bird(8, 20) <= 4; bird(8, 21) <= 4; 
bird(8, 22) <= 5; bird(8, 23) <= 0; bird(8, 24) <= 0; bird(9, 0) <= 0; 
bird(9, 1) <= 0; bird(9, 2) <= 0; bird(9, 3) <= 0; bird(9, 4) <= 0; bird(9, 5) <= 0; bird(9, 6) <= 5; bird(9, 7) <= 4; 
bird(9, 8) <= 4; bird(9, 9) <= 4; bird(9, 10) <= 4; bird(9, 11) <= 4; bird(9, 12) <= 4; bird(9, 13) <= 4; bird(9, 14) <= 4; 
bird(9, 15) <= 4; bird(9, 16) <= 4; bird(9, 17) <= 4; bird(9, 18) <= 4; bird(9, 19) <= 4; bird(9, 20) <= 4; bird(9, 21) <= 4; 
bird(9, 22) <= 4; bird(9, 23) <= 5; bird(9, 24) <= 0; bird(10, 0) <= 0; 
bird(10, 1) <= 0; bird(10, 2) <= 0; bird(10, 3) <= 0; bird(10, 4) <= 0; bird(10, 5) <= 5; bird(10, 6) <= 4; bird(10, 7) <= 4; 
bird(10, 8) <= 4; bird(10, 9) <= 4; bird(10, 10) <= 4; bird(10, 11) <= 4; bird(10, 12) <= 5; bird(10, 13) <= 5; bird(10, 14) <= 5; 
bird(10, 15) <= 5; bird(10, 16) <= 4; bird(10, 17) <= 4; bird(10, 18) <= 4; bird(10, 19) <= 4; bird(10, 20) <= 4; bird(10, 21) <= 5; 
bird(10, 22) <= 5; bird(10, 23) <= 5; bird(10, 24) <= 0; bird(11, 0) <= 5; 
bird(11, 1) <= 5; bird(11, 2) <= 5; bird(11, 3) <= 0; bird(11, 4) <= 5; bird(11, 5) <= 4; bird(11, 6) <= 4; bird(11, 7) <= 4; 
bird(11, 8) <= 4; bird(11, 9) <= 4; bird(11, 10) <= 4; bird(11, 11) <= 4; bird(11, 12) <= 4; bird(11, 13) <= 5; bird(11, 14) <= 5; 
bird(11, 15) <= 5; bird(11, 16) <= 5; bird(11, 17) <= 5; bird(11, 18) <= 4; bird(11, 19) <= 4; bird(11, 20) <= 5; bird(11, 21) <= 5; 
bird(11, 22) <= 5; bird(11, 23) <= 5; bird(11, 24) <= 5; bird(12, 0) <= 0; 
bird(12, 1) <= 5; bird(12, 2) <= 5; bird(12, 3) <= 5; bird(12, 4) <= 5; bird(12, 5) <= 4; bird(12, 6) <= 4; bird(12, 7) <= 4; 
bird(12, 8) <= 4; bird(12, 9) <= 4; bird(12, 10) <= 4; bird(12, 11) <= 4; bird(12, 12) <= 4; bird(12, 13) <= 5; bird(12, 14) <= 2; 
bird(12, 15) <= 2; bird(12, 16) <= 5; bird(12, 17) <= 5; bird(12, 18) <= 5; bird(12, 19) <= 5; bird(12, 20) <= 5; bird(12, 21) <= 5; 
bird(12, 22) <= 5; bird(12, 23) <= 4; bird(12, 24) <= 5; bird(13, 0) <= 0; 
bird(13, 1) <= 5; bird(13, 2) <= 5; bird(13, 3) <= 5; bird(13, 4) <= 5; bird(13, 5) <= 4; bird(13, 6) <= 4; bird(13, 7) <= 4; 
bird(13, 8) <= 4; bird(13, 9) <= 4; bird(13, 10) <= 4; bird(13, 11) <= 4; bird(13, 12) <= 4; bird(13, 13) <= 5; bird(13, 14) <= 2; 
bird(13, 15) <= 2; bird(13, 16) <= 2; bird(13, 17) <= 5; bird(13, 18) <= 2; bird(13, 19) <= 2; bird(13, 20) <= 5; bird(13, 21) <= 2; 
bird(13, 22) <= 5; bird(13, 23) <= 4; bird(13, 24) <= 5; bird(14, 0) <= 0; 
bird(14, 1) <= 5; bird(14, 2) <= 5; bird(14, 3) <= 5; bird(14, 4) <= 5; bird(14, 5) <= 4; bird(14, 6) <= 4; bird(14, 7) <= 4; 
bird(14, 8) <= 4; bird(14, 9) <= 4; bird(14, 10) <= 4; bird(14, 11) <= 4; bird(14, 12) <= 4; bird(14, 13) <= 4; bird(14, 14) <= 5; 
bird(14, 15) <= 2; bird(14, 16) <= 2; bird(14, 17) <= 2; bird(14, 18) <= 5; bird(14, 19) <= 5; bird(14, 20) <= 2; bird(14, 21) <= 2; 
bird(14, 22) <= 5; bird(14, 23) <= 4; bird(14, 24) <= 5; bird(15, 0) <= 0; 
bird(15, 1) <= 0; bird(15, 2) <= 0; bird(15, 3) <= 5; bird(15, 4) <= 5; bird(15, 5) <= 4; bird(15, 6) <= 4; bird(15, 7) <= 4; 
bird(15, 8) <= 4; bird(15, 9) <= 4; bird(15, 10) <= 4; bird(15, 11) <= 4; bird(15, 12) <= 4; bird(15, 13) <= 4; bird(15, 14) <= 4; 
bird(15, 15) <= 5; bird(15, 16) <= 5; bird(15, 17) <= 3; bird(15, 18) <= 3; bird(15, 19) <= 3; bird(15, 20) <= 5; bird(15, 21) <= 5; 
bird(15, 22) <= 4; bird(15, 23) <= 4; bird(15, 24) <= 5; bird(16, 0) <= 0; 
bird(16, 1) <= 5; bird(16, 2) <= 5; bird(16, 3) <= 0; bird(16, 4) <= 4; bird(16, 5) <= 4; bird(16, 6) <= 4; bird(16, 7) <= 4; 
bird(16, 8) <= 4; bird(16, 9) <= 4; bird(16, 10) <= 4; bird(16, 11) <= 4; bird(16, 12) <= 4; bird(16, 13) <= 4; bird(16, 14) <= 4; 
bird(16, 15) <= 5; bird(16, 16) <= 3; bird(16, 17) <= 3; bird(16, 18) <= 3; bird(16, 19) <= 3; bird(16, 20) <= 3; bird(16, 21) <= 3; 
bird(16, 22) <= 5; bird(16, 23) <= 4; bird(16, 24) <= 5; bird(17, 0) <= 0; 
bird(17, 1) <= 0; bird(17, 2) <= 0; bird(17, 3) <= 0; bird(17, 4) <= 5; bird(17, 5) <= 4; bird(17, 6) <= 4; bird(17, 7) <= 4; 
bird(17, 8) <= 4; bird(17, 9) <= 4; bird(17, 10) <= 4; bird(17, 11) <= 2; bird(17, 12) <= 2; bird(17, 13) <= 2; bird(17, 14) <= 2; 
bird(17, 15) <= 5; bird(17, 16) <= 3; bird(17, 17) <= 5; bird(17, 18) <= 5; bird(17, 19) <= 3; bird(17, 20) <= 3; bird(17, 21) <= 3; 
bird(17, 22) <= 3; bird(17, 23) <= 5; bird(17, 24) <= 5; bird(18, 0) <= 0; 
bird(18, 1) <= 0; bird(18, 2) <= 0; bird(18, 3) <= 0; bird(18, 4) <= 0; bird(18, 5) <= 5; bird(18, 6) <= 4; bird(18, 7) <= 4; 
bird(18, 8) <= 4; bird(18, 9) <= 4; bird(18, 10) <= 2; bird(18, 11) <= 2; bird(18, 12) <= 2; bird(18, 13) <= 2; bird(18, 14) <= 2; 
bird(18, 15) <= 2; bird(18, 16) <= 5; bird(18, 17) <= 3; bird(18, 18) <= 3; bird(18, 19) <= 5; bird(18, 20) <= 5; bird(18, 21) <= 5; 
bird(18, 22) <= 5; bird(18, 23) <= 4; bird(18, 24) <= 5; bird(19, 0) <= 0; 
bird(19, 1) <= 0; bird(19, 2) <= 0; bird(19, 3) <= 0; bird(19, 4) <= 0; bird(19, 5) <= 0; bird(19, 6) <= 5; bird(19, 7) <= 4; 
bird(19, 8) <= 4; bird(19, 9) <= 2; bird(19, 10) <= 2; bird(19, 11) <= 2; bird(19, 12) <= 2; bird(19, 13) <= 2; bird(19, 14) <= 2; 
bird(19, 15) <= 2; bird(19, 16) <= 2; bird(19, 17) <= 5; bird(19, 18) <= 5; bird(19, 19) <= 5; bird(19, 20) <= 2; bird(19, 21) <= 2; 
bird(19, 22) <= 4; bird(19, 23) <= 5; bird(19, 24) <= 0; bird(20, 0) <= 0; 
bird(20, 1) <= 0; bird(20, 2) <= 0; bird(20, 3) <= 0; bird(20, 4) <= 0; bird(20, 5) <= 0; bird(20, 6) <= 0; bird(20, 7) <= 5; 
bird(20, 8) <= 2; bird(20, 9) <= 2; bird(20, 10) <= 2; bird(20, 11) <= 2; bird(20, 12) <= 2; bird(20, 13) <= 2; bird(20, 14) <= 2; 
bird(20, 15) <= 2; bird(20, 16) <= 2; bird(20, 17) <= 2; bird(20, 18) <= 2; bird(20, 19) <= 2; bird(20, 20) <= 2; bird(20, 21) <= 2; 
bird(20, 22) <= 5; bird(20, 23) <= 0; bird(20, 24) <= 0; bird(21, 0) <= 0; 
bird(21, 1) <= 0; bird(21, 2) <= 0; bird(21, 3) <= 0; bird(21, 4) <= 0; bird(21, 5) <= 0; bird(21, 6) <= 0; bird(21, 7) <= 0; 
bird(21, 8) <= 5; bird(21, 9) <= 5; bird(21, 10) <= 2; bird(21, 11) <= 2; bird(21, 12) <= 2; bird(21, 13) <= 2; bird(21, 14) <= 2; 
bird(21, 15) <= 2; bird(21, 16) <= 2; bird(21, 17) <= 2; bird(21, 18) <= 2; bird(21, 19) <= 2; bird(21, 20) <= 2; bird(21, 21) <= 5; 
bird(21, 22) <= 0; bird(21, 23) <= 0; bird(21, 24) <= 0; bird(22, 0) <= 0; 
bird(22, 1) <= 0; bird(22, 2) <= 0; bird(22, 3) <= 0; bird(22, 4) <= 0; bird(22, 5) <= 0; bird(22, 6) <= 0; bird(22, 7) <= 0; 
bird(22, 8) <= 0; bird(22, 9) <= 0; bird(22, 10) <= 5; bird(22, 11) <= 5; bird(22, 12) <= 5; bird(22, 13) <= 5; bird(22, 14) <= 5; 
bird(22, 15) <= 5; bird(22, 16) <= 5; bird(22, 17) <= 5; bird(22, 18) <= 5; bird(22, 19) <= 5; bird(22, 20) <= 5; bird(22, 21) <= 0; 
bird(22, 22) <= 0; bird(22, 23) <= 0; bird(22, 24) <= 0; bird(23, 0) <= 0; 
bird(23, 1) <= 0; bird(23, 2) <= 0; bird(23, 3) <= 0; bird(23, 4) <= 0; bird(23, 5) <= 0; bird(23, 6) <= 0; bird(23, 7) <= 0; 
bird(23, 8) <= 0; bird(23, 9) <= 0; bird(23, 10) <= 0; bird(23, 11) <= 0; bird(23, 12) <= 0; bird(23, 13) <= 0; bird(23, 14) <= 0; 
bird(23, 15) <= 0; bird(23, 16) <= 0; bird(23, 17) <= 0; bird(23, 18) <= 0; bird(23, 19) <= 0; bird(23, 20) <= 0; bird(23, 21) <= 0; 
bird(23, 22) <= 0; bird(23, 23) <= 0; bird(23, 24) <= 0; 

end Behavioral;
