library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package papkg is
    type playAgain2D is array(0 to 19, 0 to 287) of integer;
end package;

use work.papkg.all;

entity playAgain is
    Port (playAgain_W: out playAgain2D );
end playAgain;

architecture Behavioral of playAgain is

begin

playAgain_W(0, 0) <= 1; playAgain_W(0, 1) <= 1; playAgain_W(0, 2) <= 1; playAgain_W(0, 3) <= 1; playAgain_W(0, 4) <= 1; playAgain_W(0, 5) <= 1; playAgain_W(0, 6) <= 1; playAgain_W(0, 7) <= 1; playAgain_W(0, 8) <= 1; playAgain_W(0, 9) <= 1; playAgain_W(0, 10) <= 1; playAgain_W(0, 11) <= 1; playAgain_W(0, 12) <= 0; playAgain_W(0, 13) <= 0; playAgain_W(0, 14) <= 0; playAgain_W(0, 15) <= 0; playAgain_W(0, 16) <= 0; playAgain_W(0, 17) <= 0; playAgain_W(0, 18) <= 1; playAgain_W(0, 19) <= 1; playAgain_W(0, 20) <= 1; playAgain_W(0, 21) <= 1; playAgain_W(0, 22) <= 1; playAgain_W(0, 23) <= 1; playAgain_W(0, 24) <= 1; playAgain_W(0, 25) <= 1; playAgain_W(0, 26) <= 0; playAgain_W(0, 27) <= 0; playAgain_W(0, 28) <= 0; playAgain_W(0, 29) <= 0; playAgain_W(0, 30) <= 0; playAgain_W(0, 31) <= 0; playAgain_W(0, 32) <= 0; playAgain_W(0, 33) <= 0; playAgain_W(0, 34) <= 0; playAgain_W(0, 35) <= 0; playAgain_W(0, 36) <= 0; playAgain_W(0, 37) <= 0; playAgain_W(0, 38) <= 0; playAgain_W(0, 39) <= 0; playAgain_W(0, 40) <= 0; playAgain_W(0, 41) <= 0; playAgain_W(0, 42) <= 1; playAgain_W(0, 43) <= 1; playAgain_W(0, 44) <= 0; playAgain_W(0, 45) <= 0; playAgain_W(0, 46) <= 0; playAgain_W(0, 47) <= 0; playAgain_W(0, 48) <= 0; playAgain_W(0, 49) <= 0; playAgain_W(0, 50) <= 0; playAgain_W(0, 51) <= 0; playAgain_W(0, 52) <= 0; playAgain_W(0, 53) <= 0; playAgain_W(0, 54) <= 1; playAgain_W(0, 55) <= 1; playAgain_W(0, 56) <= 1; playAgain_W(0, 57) <= 1; playAgain_W(0, 58) <= 0; playAgain_W(0, 59) <= 0; playAgain_W(0, 60) <= 0; playAgain_W(0, 61) <= 0; playAgain_W(0, 62) <= 0; playAgain_W(0, 63) <= 0; playAgain_W(0, 64) <= 0; playAgain_W(0, 65) <= 0; playAgain_W(0, 66) <= 1; playAgain_W(0, 67) <= 1; playAgain_W(0, 68) <= 1; playAgain_W(0, 69) <= 1; playAgain_W(0, 70) <= 0; playAgain_W(0, 71) <= 0; playAgain_W(0, 72) <= 0; playAgain_W(0, 73) <= 0; playAgain_W(0, 74) <= 0; playAgain_W(0, 75) <= 0; playAgain_W(0, 76) <= 0; playAgain_W(0, 77) <= 0; playAgain_W(0, 78) <= 0; playAgain_W(0, 79) <= 0; playAgain_W(0, 80) <= 0; playAgain_W(0, 81) <= 0; playAgain_W(0, 82) <= 0; playAgain_W(0, 83) <= 0; playAgain_W(0, 84) <= 0; playAgain_W(0, 85) <= 0; playAgain_W(0, 86) <= 0; playAgain_W(0, 87) <= 0; playAgain_W(0, 88) <= 0; playAgain_W(0, 89) <= 0; playAgain_W(0, 90) <= 0; playAgain_W(0, 91) <= 0; playAgain_W(0, 92) <= 0; playAgain_W(0, 93) <= 0; playAgain_W(0, 94) <= 0; playAgain_W(0, 95) <= 0; playAgain_W(0, 96) <= 1; playAgain_W(0, 97) <= 1; playAgain_W(0, 98) <= 0; playAgain_W(0, 99) <= 0; playAgain_W(0, 100) <= 0; playAgain_W(0, 101) <= 0; playAgain_W(0, 102) <= 0; playAgain_W(0, 103) <= 0; playAgain_W(0, 104) <= 0; playAgain_W(0, 105) <= 0; playAgain_W(0, 106) <= 0; playAgain_W(0, 107) <= 0; playAgain_W(0, 108) <= 0; playAgain_W(0, 109) <= 0; playAgain_W(0, 110) <= 0; playAgain_W(0, 111) <= 0; playAgain_W(0, 112) <= 1; playAgain_W(0, 113) <= 1; playAgain_W(0, 114) <= 1; playAgain_W(0, 115) <= 1; playAgain_W(0, 116) <= 1; playAgain_W(0, 117) <= 1; playAgain_W(0, 118) <= 1; playAgain_W(0, 119) <= 1; playAgain_W(0, 120) <= 0; playAgain_W(0, 121) <= 0; playAgain_W(0, 122) <= 0; playAgain_W(0, 123) <= 0; playAgain_W(0, 124) <= 0; playAgain_W(0, 125) <= 0; playAgain_W(0, 126) <= 0; playAgain_W(0, 127) <= 0; playAgain_W(0, 128) <= 0; playAgain_W(0, 129) <= 0; playAgain_W(0, 130) <= 0; playAgain_W(0, 131) <= 0; playAgain_W(0, 132) <= 1; playAgain_W(0, 133) <= 1; playAgain_W(0, 134) <= 0; playAgain_W(0, 135) <= 0; playAgain_W(0, 136) <= 0; playAgain_W(0, 137) <= 0; playAgain_W(0, 138) <= 0; playAgain_W(0, 139) <= 0; playAgain_W(0, 140) <= 0; playAgain_W(0, 141) <= 0; playAgain_W(0, 142) <= 0; playAgain_W(0, 143) <= 0; playAgain_W(0, 144) <= 0; playAgain_W(0, 145) <= 0; playAgain_W(0, 146) <= 0; playAgain_W(0, 147) <= 0; playAgain_W(0, 148) <= 1; playAgain_W(0, 149) <= 1; playAgain_W(0, 150) <= 1; playAgain_W(0, 151) <= 1; playAgain_W(0, 152) <= 1; playAgain_W(0, 153) <= 1; playAgain_W(0, 154) <= 1; playAgain_W(0, 155) <= 1; playAgain_W(0, 156) <= 0; playAgain_W(0, 157) <= 0; playAgain_W(0, 158) <= 0; playAgain_W(0, 159) <= 0; playAgain_W(0, 160) <= 0; playAgain_W(0, 161) <= 0; playAgain_W(0, 162) <= 1; playAgain_W(0, 163) <= 1; playAgain_W(0, 164) <= 1; playAgain_W(0, 165) <= 1; playAgain_W(0, 166) <= 0; playAgain_W(0, 167) <= 0; playAgain_W(0, 168) <= 0; playAgain_W(0, 169) <= 0; playAgain_W(0, 170) <= 0; playAgain_W(0, 171) <= 0; playAgain_W(0, 172) <= 1; playAgain_W(0, 173) <= 1; playAgain_W(0, 174) <= 1; playAgain_W(0, 175) <= 1; playAgain_W(0, 176) <= 0; playAgain_W(0, 177) <= 0; playAgain_W(0, 178) <= 0; playAgain_W(0, 179) <= 0; playAgain_W(0, 180) <= 0; playAgain_W(0, 181) <= 0; playAgain_W(0, 182) <= 0; playAgain_W(0, 183) <= 0; playAgain_W(0, 184) <= 0; playAgain_W(0, 185) <= 0; playAgain_W(0, 186) <= 0; playAgain_W(0, 187) <= 0; playAgain_W(0, 188) <= 0; playAgain_W(0, 189) <= 0; playAgain_W(0, 190) <= 0; playAgain_W(0, 191) <= 0; playAgain_W(0, 192) <= 0; playAgain_W(0, 193) <= 0; playAgain_W(0, 194) <= 0; playAgain_W(0, 195) <= 0; playAgain_W(0, 196) <= 0; playAgain_W(0, 197) <= 0; playAgain_W(0, 198) <= 0; playAgain_W(0, 199) <= 0; playAgain_W(0, 200) <= 0; playAgain_W(0, 201) <= 0; playAgain_W(0, 202) <= 0; playAgain_W(0, 203) <= 0; playAgain_W(0, 204) <= 0; playAgain_W(0, 205) <= 0; playAgain_W(0, 206) <= 0; playAgain_W(0, 207) <= 0; playAgain_W(0, 208) <= 0; playAgain_W(0, 209) <= 0; playAgain_W(0, 210) <= 0; playAgain_W(0, 211) <= 0; playAgain_W(0, 212) <= 0; playAgain_W(0, 213) <= 0; playAgain_W(0, 214) <= 0; playAgain_W(0, 215) <= 0; playAgain_W(0, 216) <= 1; playAgain_W(0, 217) <= 1; playAgain_W(0, 218) <= 1; playAgain_W(0, 219) <= 1; playAgain_W(0, 220) <= 1; playAgain_W(0, 221) <= 1; playAgain_W(0, 222) <= 1; playAgain_W(0, 223) <= 1; playAgain_W(0, 224) <= 1; playAgain_W(0, 225) <= 1; playAgain_W(0, 226) <= 1; playAgain_W(0, 227) <= 1; playAgain_W(0, 228) <= 0; playAgain_W(0, 229) <= 0; playAgain_W(0, 230) <= 0; playAgain_W(0, 231) <= 0; playAgain_W(0, 232) <= 0; playAgain_W(0, 233) <= 0; playAgain_W(0, 234) <= 1; playAgain_W(0, 235) <= 1; playAgain_W(0, 236) <= 1; playAgain_W(0, 237) <= 1; playAgain_W(0, 238) <= 1; playAgain_W(0, 239) <= 1; playAgain_W(0, 240) <= 1; playAgain_W(0, 241) <= 1; playAgain_W(0, 242) <= 1; playAgain_W(0, 243) <= 1; playAgain_W(0, 244) <= 1; playAgain_W(0, 245) <= 1; playAgain_W(0, 246) <= 1; playAgain_W(0, 247) <= 1; playAgain_W(0, 248) <= 1; playAgain_W(0, 249) <= 1; playAgain_W(0, 250) <= 0; playAgain_W(0, 251) <= 0; playAgain_W(0, 252) <= 1; playAgain_W(0, 253) <= 1; playAgain_W(0, 254) <= 1; playAgain_W(0, 255) <= 1; playAgain_W(0, 256) <= 0; playAgain_W(0, 257) <= 0; playAgain_W(0, 258) <= 0; playAgain_W(0, 259) <= 0; playAgain_W(0, 260) <= 0; playAgain_W(0, 261) <= 0; playAgain_W(0, 262) <= 1; playAgain_W(0, 263) <= 1; playAgain_W(0, 264) <= 1; playAgain_W(0, 265) <= 1; playAgain_W(0, 266) <= 0; playAgain_W(0, 267) <= 0; playAgain_W(0, 268) <= 0; playAgain_W(0, 269) <= 0; playAgain_W(0, 270) <= 1; playAgain_W(0, 271) <= 1; playAgain_W(0, 272) <= 1; playAgain_W(0, 273) <= 1; playAgain_W(0, 274) <= 1; playAgain_W(0, 275) <= 1; playAgain_W(0, 276) <= 1; playAgain_W(0, 277) <= 1; playAgain_W(0, 278) <= 1; playAgain_W(0, 279) <= 1; playAgain_W(0, 280) <= 0; playAgain_W(0, 281) <= 0; playAgain_W(0, 282) <= 0; playAgain_W(0, 283) <= 0; playAgain_W(0, 284) <= 0; playAgain_W(0, 285) <= 0; playAgain_W(0, 286) <= 0; playAgain_W(0, 287) <= 0; 
playAgain_W(1, 0) <= 1; playAgain_W(1, 1) <= 1; playAgain_W(1, 2) <= 1; playAgain_W(1, 3) <= 1; playAgain_W(1, 4) <= 1; playAgain_W(1, 5) <= 1; playAgain_W(1, 6) <= 1; playAgain_W(1, 7) <= 1; playAgain_W(1, 8) <= 1; playAgain_W(1, 9) <= 1; playAgain_W(1, 10) <= 1; playAgain_W(1, 11) <= 1; playAgain_W(1, 12) <= 0; playAgain_W(1, 13) <= 0; playAgain_W(1, 14) <= 0; playAgain_W(1, 15) <= 0; playAgain_W(1, 16) <= 0; playAgain_W(1, 17) <= 0; playAgain_W(1, 18) <= 1; playAgain_W(1, 19) <= 1; playAgain_W(1, 20) <= 1; playAgain_W(1, 21) <= 1; playAgain_W(1, 22) <= 1; playAgain_W(1, 23) <= 1; playAgain_W(1, 24) <= 1; playAgain_W(1, 25) <= 1; playAgain_W(1, 26) <= 0; playAgain_W(1, 27) <= 0; playAgain_W(1, 28) <= 0; playAgain_W(1, 29) <= 0; playAgain_W(1, 30) <= 0; playAgain_W(1, 31) <= 0; playAgain_W(1, 32) <= 0; playAgain_W(1, 33) <= 0; playAgain_W(1, 34) <= 0; playAgain_W(1, 35) <= 0; playAgain_W(1, 36) <= 0; playAgain_W(1, 37) <= 0; playAgain_W(1, 38) <= 0; playAgain_W(1, 39) <= 0; playAgain_W(1, 40) <= 0; playAgain_W(1, 41) <= 0; playAgain_W(1, 42) <= 1; playAgain_W(1, 43) <= 1; playAgain_W(1, 44) <= 0; playAgain_W(1, 45) <= 0; playAgain_W(1, 46) <= 0; playAgain_W(1, 47) <= 0; playAgain_W(1, 48) <= 0; playAgain_W(1, 49) <= 0; playAgain_W(1, 50) <= 0; playAgain_W(1, 51) <= 0; playAgain_W(1, 52) <= 0; playAgain_W(1, 53) <= 0; playAgain_W(1, 54) <= 1; playAgain_W(1, 55) <= 1; playAgain_W(1, 56) <= 1; playAgain_W(1, 57) <= 1; playAgain_W(1, 58) <= 0; playAgain_W(1, 59) <= 0; playAgain_W(1, 60) <= 0; playAgain_W(1, 61) <= 0; playAgain_W(1, 62) <= 0; playAgain_W(1, 63) <= 0; playAgain_W(1, 64) <= 0; playAgain_W(1, 65) <= 0; playAgain_W(1, 66) <= 1; playAgain_W(1, 67) <= 1; playAgain_W(1, 68) <= 1; playAgain_W(1, 69) <= 1; playAgain_W(1, 70) <= 0; playAgain_W(1, 71) <= 0; playAgain_W(1, 72) <= 0; playAgain_W(1, 73) <= 0; playAgain_W(1, 74) <= 0; playAgain_W(1, 75) <= 0; playAgain_W(1, 76) <= 0; playAgain_W(1, 77) <= 0; playAgain_W(1, 78) <= 0; playAgain_W(1, 79) <= 0; playAgain_W(1, 80) <= 0; playAgain_W(1, 81) <= 0; playAgain_W(1, 82) <= 0; playAgain_W(1, 83) <= 0; playAgain_W(1, 84) <= 0; playAgain_W(1, 85) <= 0; playAgain_W(1, 86) <= 0; playAgain_W(1, 87) <= 0; playAgain_W(1, 88) <= 0; playAgain_W(1, 89) <= 0; playAgain_W(1, 90) <= 0; playAgain_W(1, 91) <= 0; playAgain_W(1, 92) <= 0; playAgain_W(1, 93) <= 0; playAgain_W(1, 94) <= 0; playAgain_W(1, 95) <= 0; playAgain_W(1, 96) <= 1; playAgain_W(1, 97) <= 1; playAgain_W(1, 98) <= 0; playAgain_W(1, 99) <= 0; playAgain_W(1, 100) <= 0; playAgain_W(1, 101) <= 0; playAgain_W(1, 102) <= 0; playAgain_W(1, 103) <= 0; playAgain_W(1, 104) <= 0; playAgain_W(1, 105) <= 0; playAgain_W(1, 106) <= 0; playAgain_W(1, 107) <= 0; playAgain_W(1, 108) <= 0; playAgain_W(1, 109) <= 0; playAgain_W(1, 110) <= 0; playAgain_W(1, 111) <= 0; playAgain_W(1, 112) <= 1; playAgain_W(1, 113) <= 1; playAgain_W(1, 114) <= 1; playAgain_W(1, 115) <= 1; playAgain_W(1, 116) <= 1; playAgain_W(1, 117) <= 1; playAgain_W(1, 118) <= 1; playAgain_W(1, 119) <= 1; playAgain_W(1, 120) <= 0; playAgain_W(1, 121) <= 0; playAgain_W(1, 122) <= 0; playAgain_W(1, 123) <= 0; playAgain_W(1, 124) <= 0; playAgain_W(1, 125) <= 0; playAgain_W(1, 126) <= 0; playAgain_W(1, 127) <= 0; playAgain_W(1, 128) <= 0; playAgain_W(1, 129) <= 0; playAgain_W(1, 130) <= 0; playAgain_W(1, 131) <= 0; playAgain_W(1, 132) <= 1; playAgain_W(1, 133) <= 1; playAgain_W(1, 134) <= 0; playAgain_W(1, 135) <= 0; playAgain_W(1, 136) <= 0; playAgain_W(1, 137) <= 0; playAgain_W(1, 138) <= 0; playAgain_W(1, 139) <= 0; playAgain_W(1, 140) <= 0; playAgain_W(1, 141) <= 0; playAgain_W(1, 142) <= 0; playAgain_W(1, 143) <= 0; playAgain_W(1, 144) <= 0; playAgain_W(1, 145) <= 0; playAgain_W(1, 146) <= 0; playAgain_W(1, 147) <= 0; playAgain_W(1, 148) <= 1; playAgain_W(1, 149) <= 1; playAgain_W(1, 150) <= 1; playAgain_W(1, 151) <= 1; playAgain_W(1, 152) <= 1; playAgain_W(1, 153) <= 1; playAgain_W(1, 154) <= 1; playAgain_W(1, 155) <= 1; playAgain_W(1, 156) <= 0; playAgain_W(1, 157) <= 0; playAgain_W(1, 158) <= 0; playAgain_W(1, 159) <= 0; playAgain_W(1, 160) <= 0; playAgain_W(1, 161) <= 0; playAgain_W(1, 162) <= 1; playAgain_W(1, 163) <= 1; playAgain_W(1, 164) <= 1; playAgain_W(1, 165) <= 1; playAgain_W(1, 166) <= 0; playAgain_W(1, 167) <= 0; playAgain_W(1, 168) <= 0; playAgain_W(1, 169) <= 0; playAgain_W(1, 170) <= 0; playAgain_W(1, 171) <= 0; playAgain_W(1, 172) <= 1; playAgain_W(1, 173) <= 1; playAgain_W(1, 174) <= 1; playAgain_W(1, 175) <= 1; playAgain_W(1, 176) <= 0; playAgain_W(1, 177) <= 0; playAgain_W(1, 178) <= 0; playAgain_W(1, 179) <= 0; playAgain_W(1, 180) <= 0; playAgain_W(1, 181) <= 0; playAgain_W(1, 182) <= 0; playAgain_W(1, 183) <= 0; playAgain_W(1, 184) <= 0; playAgain_W(1, 185) <= 0; playAgain_W(1, 186) <= 0; playAgain_W(1, 187) <= 0; playAgain_W(1, 188) <= 0; playAgain_W(1, 189) <= 0; playAgain_W(1, 190) <= 0; playAgain_W(1, 191) <= 0; playAgain_W(1, 192) <= 0; playAgain_W(1, 193) <= 0; playAgain_W(1, 194) <= 0; playAgain_W(1, 195) <= 0; playAgain_W(1, 196) <= 0; playAgain_W(1, 197) <= 0; playAgain_W(1, 198) <= 0; playAgain_W(1, 199) <= 0; playAgain_W(1, 200) <= 0; playAgain_W(1, 201) <= 0; playAgain_W(1, 202) <= 0; playAgain_W(1, 203) <= 0; playAgain_W(1, 204) <= 0; playAgain_W(1, 205) <= 0; playAgain_W(1, 206) <= 0; playAgain_W(1, 207) <= 0; playAgain_W(1, 208) <= 0; playAgain_W(1, 209) <= 0; playAgain_W(1, 210) <= 0; playAgain_W(1, 211) <= 0; playAgain_W(1, 212) <= 0; playAgain_W(1, 213) <= 0; playAgain_W(1, 214) <= 0; playAgain_W(1, 215) <= 0; playAgain_W(1, 216) <= 1; playAgain_W(1, 217) <= 1; playAgain_W(1, 218) <= 1; playAgain_W(1, 219) <= 1; playAgain_W(1, 220) <= 1; playAgain_W(1, 221) <= 1; playAgain_W(1, 222) <= 1; playAgain_W(1, 223) <= 1; playAgain_W(1, 224) <= 1; playAgain_W(1, 225) <= 1; playAgain_W(1, 226) <= 1; playAgain_W(1, 227) <= 1; playAgain_W(1, 228) <= 0; playAgain_W(1, 229) <= 0; playAgain_W(1, 230) <= 0; playAgain_W(1, 231) <= 0; playAgain_W(1, 232) <= 0; playAgain_W(1, 233) <= 0; playAgain_W(1, 234) <= 1; playAgain_W(1, 235) <= 1; playAgain_W(1, 236) <= 1; playAgain_W(1, 237) <= 1; playAgain_W(1, 238) <= 1; playAgain_W(1, 239) <= 1; playAgain_W(1, 240) <= 1; playAgain_W(1, 241) <= 1; playAgain_W(1, 242) <= 1; playAgain_W(1, 243) <= 1; playAgain_W(1, 244) <= 1; playAgain_W(1, 245) <= 1; playAgain_W(1, 246) <= 1; playAgain_W(1, 247) <= 1; playAgain_W(1, 248) <= 1; playAgain_W(1, 249) <= 1; playAgain_W(1, 250) <= 0; playAgain_W(1, 251) <= 0; playAgain_W(1, 252) <= 1; playAgain_W(1, 253) <= 1; playAgain_W(1, 254) <= 1; playAgain_W(1, 255) <= 1; playAgain_W(1, 256) <= 0; playAgain_W(1, 257) <= 0; playAgain_W(1, 258) <= 0; playAgain_W(1, 259) <= 0; playAgain_W(1, 260) <= 0; playAgain_W(1, 261) <= 0; playAgain_W(1, 262) <= 1; playAgain_W(1, 263) <= 1; playAgain_W(1, 264) <= 1; playAgain_W(1, 265) <= 1; playAgain_W(1, 266) <= 0; playAgain_W(1, 267) <= 0; playAgain_W(1, 268) <= 0; playAgain_W(1, 269) <= 0; playAgain_W(1, 270) <= 1; playAgain_W(1, 271) <= 1; playAgain_W(1, 272) <= 1; playAgain_W(1, 273) <= 1; playAgain_W(1, 274) <= 1; playAgain_W(1, 275) <= 1; playAgain_W(1, 276) <= 1; playAgain_W(1, 277) <= 1; playAgain_W(1, 278) <= 1; playAgain_W(1, 279) <= 1; playAgain_W(1, 280) <= 0; playAgain_W(1, 281) <= 0; playAgain_W(1, 282) <= 0; playAgain_W(1, 283) <= 0; playAgain_W(1, 284) <= 0; playAgain_W(1, 285) <= 0; playAgain_W(1, 286) <= 0; playAgain_W(1, 287) <= 0; 
playAgain_W(2, 0) <= 0; playAgain_W(2, 1) <= 0; playAgain_W(2, 2) <= 1; playAgain_W(2, 3) <= 1; playAgain_W(2, 4) <= 1; playAgain_W(2, 5) <= 1; playAgain_W(2, 6) <= 0; playAgain_W(2, 7) <= 0; playAgain_W(2, 8) <= 0; playAgain_W(2, 9) <= 0; playAgain_W(2, 10) <= 1; playAgain_W(2, 11) <= 1; playAgain_W(2, 12) <= 1; playAgain_W(2, 13) <= 1; playAgain_W(2, 14) <= 0; playAgain_W(2, 15) <= 0; playAgain_W(2, 16) <= 0; playAgain_W(2, 17) <= 0; playAgain_W(2, 18) <= 0; playAgain_W(2, 19) <= 0; playAgain_W(2, 20) <= 1; playAgain_W(2, 21) <= 1; playAgain_W(2, 22) <= 1; playAgain_W(2, 23) <= 1; playAgain_W(2, 24) <= 0; playAgain_W(2, 25) <= 0; playAgain_W(2, 26) <= 0; playAgain_W(2, 27) <= 0; playAgain_W(2, 28) <= 0; playAgain_W(2, 29) <= 0; playAgain_W(2, 30) <= 0; playAgain_W(2, 31) <= 0; playAgain_W(2, 32) <= 0; playAgain_W(2, 33) <= 0; playAgain_W(2, 34) <= 0; playAgain_W(2, 35) <= 0; playAgain_W(2, 36) <= 0; playAgain_W(2, 37) <= 0; playAgain_W(2, 38) <= 0; playAgain_W(2, 39) <= 0; playAgain_W(2, 40) <= 1; playAgain_W(2, 41) <= 1; playAgain_W(2, 42) <= 1; playAgain_W(2, 43) <= 1; playAgain_W(2, 44) <= 1; playAgain_W(2, 45) <= 1; playAgain_W(2, 46) <= 0; playAgain_W(2, 47) <= 0; playAgain_W(2, 48) <= 0; playAgain_W(2, 49) <= 0; playAgain_W(2, 50) <= 0; playAgain_W(2, 51) <= 0; playAgain_W(2, 52) <= 0; playAgain_W(2, 53) <= 0; playAgain_W(2, 54) <= 1; playAgain_W(2, 55) <= 1; playAgain_W(2, 56) <= 1; playAgain_W(2, 57) <= 1; playAgain_W(2, 58) <= 0; playAgain_W(2, 59) <= 0; playAgain_W(2, 60) <= 0; playAgain_W(2, 61) <= 0; playAgain_W(2, 62) <= 0; playAgain_W(2, 63) <= 0; playAgain_W(2, 64) <= 0; playAgain_W(2, 65) <= 0; playAgain_W(2, 66) <= 1; playAgain_W(2, 67) <= 1; playAgain_W(2, 68) <= 1; playAgain_W(2, 69) <= 1; playAgain_W(2, 70) <= 0; playAgain_W(2, 71) <= 0; playAgain_W(2, 72) <= 0; playAgain_W(2, 73) <= 0; playAgain_W(2, 74) <= 0; playAgain_W(2, 75) <= 0; playAgain_W(2, 76) <= 0; playAgain_W(2, 77) <= 0; playAgain_W(2, 78) <= 0; playAgain_W(2, 79) <= 0; playAgain_W(2, 80) <= 0; playAgain_W(2, 81) <= 0; playAgain_W(2, 82) <= 0; playAgain_W(2, 83) <= 0; playAgain_W(2, 84) <= 0; playAgain_W(2, 85) <= 0; playAgain_W(2, 86) <= 0; playAgain_W(2, 87) <= 0; playAgain_W(2, 88) <= 0; playAgain_W(2, 89) <= 0; playAgain_W(2, 90) <= 0; playAgain_W(2, 91) <= 0; playAgain_W(2, 92) <= 0; playAgain_W(2, 93) <= 0; playAgain_W(2, 94) <= 1; playAgain_W(2, 95) <= 1; playAgain_W(2, 96) <= 1; playAgain_W(2, 97) <= 1; playAgain_W(2, 98) <= 1; playAgain_W(2, 99) <= 1; playAgain_W(2, 100) <= 0; playAgain_W(2, 101) <= 0; playAgain_W(2, 102) <= 0; playAgain_W(2, 103) <= 0; playAgain_W(2, 104) <= 0; playAgain_W(2, 105) <= 0; playAgain_W(2, 106) <= 0; playAgain_W(2, 107) <= 0; playAgain_W(2, 108) <= 0; playAgain_W(2, 109) <= 0; playAgain_W(2, 110) <= 1; playAgain_W(2, 111) <= 1; playAgain_W(2, 112) <= 1; playAgain_W(2, 113) <= 1; playAgain_W(2, 114) <= 0; playAgain_W(2, 115) <= 0; playAgain_W(2, 116) <= 0; playAgain_W(2, 117) <= 0; playAgain_W(2, 118) <= 1; playAgain_W(2, 119) <= 1; playAgain_W(2, 120) <= 1; playAgain_W(2, 121) <= 1; playAgain_W(2, 122) <= 0; playAgain_W(2, 123) <= 0; playAgain_W(2, 124) <= 0; playAgain_W(2, 125) <= 0; playAgain_W(2, 126) <= 0; playAgain_W(2, 127) <= 0; playAgain_W(2, 128) <= 0; playAgain_W(2, 129) <= 0; playAgain_W(2, 130) <= 1; playAgain_W(2, 131) <= 1; playAgain_W(2, 132) <= 1; playAgain_W(2, 133) <= 1; playAgain_W(2, 134) <= 1; playAgain_W(2, 135) <= 1; playAgain_W(2, 136) <= 0; playAgain_W(2, 137) <= 0; playAgain_W(2, 138) <= 0; playAgain_W(2, 139) <= 0; playAgain_W(2, 140) <= 0; playAgain_W(2, 141) <= 0; playAgain_W(2, 142) <= 0; playAgain_W(2, 143) <= 0; playAgain_W(2, 144) <= 0; playAgain_W(2, 145) <= 0; playAgain_W(2, 146) <= 0; playAgain_W(2, 147) <= 0; playAgain_W(2, 148) <= 0; playAgain_W(2, 149) <= 0; playAgain_W(2, 150) <= 1; playAgain_W(2, 151) <= 1; playAgain_W(2, 152) <= 1; playAgain_W(2, 153) <= 1; playAgain_W(2, 154) <= 0; playAgain_W(2, 155) <= 0; playAgain_W(2, 156) <= 0; playAgain_W(2, 157) <= 0; playAgain_W(2, 158) <= 0; playAgain_W(2, 159) <= 0; playAgain_W(2, 160) <= 0; playAgain_W(2, 161) <= 0; playAgain_W(2, 162) <= 1; playAgain_W(2, 163) <= 1; playAgain_W(2, 164) <= 1; playAgain_W(2, 165) <= 1; playAgain_W(2, 166) <= 1; playAgain_W(2, 167) <= 1; playAgain_W(2, 168) <= 0; playAgain_W(2, 169) <= 0; playAgain_W(2, 170) <= 0; playAgain_W(2, 171) <= 0; playAgain_W(2, 172) <= 1; playAgain_W(2, 173) <= 1; playAgain_W(2, 174) <= 1; playAgain_W(2, 175) <= 1; playAgain_W(2, 176) <= 0; playAgain_W(2, 177) <= 0; playAgain_W(2, 178) <= 0; playAgain_W(2, 179) <= 0; playAgain_W(2, 180) <= 0; playAgain_W(2, 181) <= 0; playAgain_W(2, 182) <= 0; playAgain_W(2, 183) <= 0; playAgain_W(2, 184) <= 0; playAgain_W(2, 185) <= 0; playAgain_W(2, 186) <= 0; playAgain_W(2, 187) <= 0; playAgain_W(2, 188) <= 0; playAgain_W(2, 189) <= 0; playAgain_W(2, 190) <= 0; playAgain_W(2, 191) <= 0; playAgain_W(2, 192) <= 0; playAgain_W(2, 193) <= 0; playAgain_W(2, 194) <= 0; playAgain_W(2, 195) <= 0; playAgain_W(2, 196) <= 0; playAgain_W(2, 197) <= 0; playAgain_W(2, 198) <= 0; playAgain_W(2, 199) <= 0; playAgain_W(2, 200) <= 0; playAgain_W(2, 201) <= 0; playAgain_W(2, 202) <= 0; playAgain_W(2, 203) <= 0; playAgain_W(2, 204) <= 0; playAgain_W(2, 205) <= 0; playAgain_W(2, 206) <= 0; playAgain_W(2, 207) <= 0; playAgain_W(2, 208) <= 0; playAgain_W(2, 209) <= 0; playAgain_W(2, 210) <= 0; playAgain_W(2, 211) <= 0; playAgain_W(2, 212) <= 0; playAgain_W(2, 213) <= 0; playAgain_W(2, 214) <= 0; playAgain_W(2, 215) <= 0; playAgain_W(2, 216) <= 0; playAgain_W(2, 217) <= 0; playAgain_W(2, 218) <= 1; playAgain_W(2, 219) <= 1; playAgain_W(2, 220) <= 1; playAgain_W(2, 221) <= 1; playAgain_W(2, 222) <= 0; playAgain_W(2, 223) <= 0; playAgain_W(2, 224) <= 0; playAgain_W(2, 225) <= 0; playAgain_W(2, 226) <= 1; playAgain_W(2, 227) <= 1; playAgain_W(2, 228) <= 1; playAgain_W(2, 229) <= 1; playAgain_W(2, 230) <= 0; playAgain_W(2, 231) <= 0; playAgain_W(2, 232) <= 0; playAgain_W(2, 233) <= 0; playAgain_W(2, 234) <= 1; playAgain_W(2, 235) <= 1; playAgain_W(2, 236) <= 1; playAgain_W(2, 237) <= 1; playAgain_W(2, 238) <= 0; playAgain_W(2, 239) <= 0; playAgain_W(2, 240) <= 1; playAgain_W(2, 241) <= 1; playAgain_W(2, 242) <= 1; playAgain_W(2, 243) <= 1; playAgain_W(2, 244) <= 0; playAgain_W(2, 245) <= 0; playAgain_W(2, 246) <= 1; playAgain_W(2, 247) <= 1; playAgain_W(2, 248) <= 1; playAgain_W(2, 249) <= 1; playAgain_W(2, 250) <= 0; playAgain_W(2, 251) <= 0; playAgain_W(2, 252) <= 1; playAgain_W(2, 253) <= 1; playAgain_W(2, 254) <= 1; playAgain_W(2, 255) <= 1; playAgain_W(2, 256) <= 1; playAgain_W(2, 257) <= 1; playAgain_W(2, 258) <= 0; playAgain_W(2, 259) <= 0; playAgain_W(2, 260) <= 0; playAgain_W(2, 261) <= 0; playAgain_W(2, 262) <= 1; playAgain_W(2, 263) <= 1; playAgain_W(2, 264) <= 1; playAgain_W(2, 265) <= 1; playAgain_W(2, 266) <= 0; playAgain_W(2, 267) <= 0; playAgain_W(2, 268) <= 0; playAgain_W(2, 269) <= 0; playAgain_W(2, 270) <= 0; playAgain_W(2, 271) <= 0; playAgain_W(2, 272) <= 1; playAgain_W(2, 273) <= 1; playAgain_W(2, 274) <= 1; playAgain_W(2, 275) <= 1; playAgain_W(2, 276) <= 0; playAgain_W(2, 277) <= 0; playAgain_W(2, 278) <= 1; playAgain_W(2, 279) <= 1; playAgain_W(2, 280) <= 1; playAgain_W(2, 281) <= 1; playAgain_W(2, 282) <= 0; playAgain_W(2, 283) <= 0; playAgain_W(2, 284) <= 0; playAgain_W(2, 285) <= 0; playAgain_W(2, 286) <= 0; playAgain_W(2, 287) <= 0; 
playAgain_W(3, 0) <= 0; playAgain_W(3, 1) <= 0; playAgain_W(3, 2) <= 1; playAgain_W(3, 3) <= 1; playAgain_W(3, 4) <= 1; playAgain_W(3, 5) <= 1; playAgain_W(3, 6) <= 0; playAgain_W(3, 7) <= 0; playAgain_W(3, 8) <= 0; playAgain_W(3, 9) <= 0; playAgain_W(3, 10) <= 1; playAgain_W(3, 11) <= 1; playAgain_W(3, 12) <= 1; playAgain_W(3, 13) <= 1; playAgain_W(3, 14) <= 0; playAgain_W(3, 15) <= 0; playAgain_W(3, 16) <= 0; playAgain_W(3, 17) <= 0; playAgain_W(3, 18) <= 0; playAgain_W(3, 19) <= 0; playAgain_W(3, 20) <= 1; playAgain_W(3, 21) <= 1; playAgain_W(3, 22) <= 1; playAgain_W(3, 23) <= 1; playAgain_W(3, 24) <= 0; playAgain_W(3, 25) <= 0; playAgain_W(3, 26) <= 0; playAgain_W(3, 27) <= 0; playAgain_W(3, 28) <= 0; playAgain_W(3, 29) <= 0; playAgain_W(3, 30) <= 0; playAgain_W(3, 31) <= 0; playAgain_W(3, 32) <= 0; playAgain_W(3, 33) <= 0; playAgain_W(3, 34) <= 0; playAgain_W(3, 35) <= 0; playAgain_W(3, 36) <= 0; playAgain_W(3, 37) <= 0; playAgain_W(3, 38) <= 0; playAgain_W(3, 39) <= 0; playAgain_W(3, 40) <= 1; playAgain_W(3, 41) <= 1; playAgain_W(3, 42) <= 1; playAgain_W(3, 43) <= 1; playAgain_W(3, 44) <= 1; playAgain_W(3, 45) <= 1; playAgain_W(3, 46) <= 0; playAgain_W(3, 47) <= 0; playAgain_W(3, 48) <= 0; playAgain_W(3, 49) <= 0; playAgain_W(3, 50) <= 0; playAgain_W(3, 51) <= 0; playAgain_W(3, 52) <= 0; playAgain_W(3, 53) <= 0; playAgain_W(3, 54) <= 1; playAgain_W(3, 55) <= 1; playAgain_W(3, 56) <= 1; playAgain_W(3, 57) <= 1; playAgain_W(3, 58) <= 0; playAgain_W(3, 59) <= 0; playAgain_W(3, 60) <= 0; playAgain_W(3, 61) <= 0; playAgain_W(3, 62) <= 0; playAgain_W(3, 63) <= 0; playAgain_W(3, 64) <= 0; playAgain_W(3, 65) <= 0; playAgain_W(3, 66) <= 1; playAgain_W(3, 67) <= 1; playAgain_W(3, 68) <= 1; playAgain_W(3, 69) <= 1; playAgain_W(3, 70) <= 0; playAgain_W(3, 71) <= 0; playAgain_W(3, 72) <= 0; playAgain_W(3, 73) <= 0; playAgain_W(3, 74) <= 0; playAgain_W(3, 75) <= 0; playAgain_W(3, 76) <= 0; playAgain_W(3, 77) <= 0; playAgain_W(3, 78) <= 0; playAgain_W(3, 79) <= 0; playAgain_W(3, 80) <= 0; playAgain_W(3, 81) <= 0; playAgain_W(3, 82) <= 0; playAgain_W(3, 83) <= 0; playAgain_W(3, 84) <= 0; playAgain_W(3, 85) <= 0; playAgain_W(3, 86) <= 0; playAgain_W(3, 87) <= 0; playAgain_W(3, 88) <= 0; playAgain_W(3, 89) <= 0; playAgain_W(3, 90) <= 0; playAgain_W(3, 91) <= 0; playAgain_W(3, 92) <= 0; playAgain_W(3, 93) <= 0; playAgain_W(3, 94) <= 1; playAgain_W(3, 95) <= 1; playAgain_W(3, 96) <= 1; playAgain_W(3, 97) <= 1; playAgain_W(3, 98) <= 1; playAgain_W(3, 99) <= 1; playAgain_W(3, 100) <= 0; playAgain_W(3, 101) <= 0; playAgain_W(3, 102) <= 0; playAgain_W(3, 103) <= 0; playAgain_W(3, 104) <= 0; playAgain_W(3, 105) <= 0; playAgain_W(3, 106) <= 0; playAgain_W(3, 107) <= 0; playAgain_W(3, 108) <= 0; playAgain_W(3, 109) <= 0; playAgain_W(3, 110) <= 1; playAgain_W(3, 111) <= 1; playAgain_W(3, 112) <= 1; playAgain_W(3, 113) <= 1; playAgain_W(3, 114) <= 0; playAgain_W(3, 115) <= 0; playAgain_W(3, 116) <= 0; playAgain_W(3, 117) <= 0; playAgain_W(3, 118) <= 1; playAgain_W(3, 119) <= 1; playAgain_W(3, 120) <= 1; playAgain_W(3, 121) <= 1; playAgain_W(3, 122) <= 0; playAgain_W(3, 123) <= 0; playAgain_W(3, 124) <= 0; playAgain_W(3, 125) <= 0; playAgain_W(3, 126) <= 0; playAgain_W(3, 127) <= 0; playAgain_W(3, 128) <= 0; playAgain_W(3, 129) <= 0; playAgain_W(3, 130) <= 1; playAgain_W(3, 131) <= 1; playAgain_W(3, 132) <= 1; playAgain_W(3, 133) <= 1; playAgain_W(3, 134) <= 1; playAgain_W(3, 135) <= 1; playAgain_W(3, 136) <= 0; playAgain_W(3, 137) <= 0; playAgain_W(3, 138) <= 0; playAgain_W(3, 139) <= 0; playAgain_W(3, 140) <= 0; playAgain_W(3, 141) <= 0; playAgain_W(3, 142) <= 0; playAgain_W(3, 143) <= 0; playAgain_W(3, 144) <= 0; playAgain_W(3, 145) <= 0; playAgain_W(3, 146) <= 0; playAgain_W(3, 147) <= 0; playAgain_W(3, 148) <= 0; playAgain_W(3, 149) <= 0; playAgain_W(3, 150) <= 1; playAgain_W(3, 151) <= 1; playAgain_W(3, 152) <= 1; playAgain_W(3, 153) <= 1; playAgain_W(3, 154) <= 0; playAgain_W(3, 155) <= 0; playAgain_W(3, 156) <= 0; playAgain_W(3, 157) <= 0; playAgain_W(3, 158) <= 0; playAgain_W(3, 159) <= 0; playAgain_W(3, 160) <= 0; playAgain_W(3, 161) <= 0; playAgain_W(3, 162) <= 1; playAgain_W(3, 163) <= 1; playAgain_W(3, 164) <= 1; playAgain_W(3, 165) <= 1; playAgain_W(3, 166) <= 1; playAgain_W(3, 167) <= 1; playAgain_W(3, 168) <= 0; playAgain_W(3, 169) <= 0; playAgain_W(3, 170) <= 0; playAgain_W(3, 171) <= 0; playAgain_W(3, 172) <= 1; playAgain_W(3, 173) <= 1; playAgain_W(3, 174) <= 1; playAgain_W(3, 175) <= 1; playAgain_W(3, 176) <= 0; playAgain_W(3, 177) <= 0; playAgain_W(3, 178) <= 0; playAgain_W(3, 179) <= 0; playAgain_W(3, 180) <= 0; playAgain_W(3, 181) <= 0; playAgain_W(3, 182) <= 0; playAgain_W(3, 183) <= 0; playAgain_W(3, 184) <= 0; playAgain_W(3, 185) <= 0; playAgain_W(3, 186) <= 0; playAgain_W(3, 187) <= 0; playAgain_W(3, 188) <= 0; playAgain_W(3, 189) <= 0; playAgain_W(3, 190) <= 0; playAgain_W(3, 191) <= 0; playAgain_W(3, 192) <= 0; playAgain_W(3, 193) <= 0; playAgain_W(3, 194) <= 0; playAgain_W(3, 195) <= 0; playAgain_W(3, 196) <= 0; playAgain_W(3, 197) <= 0; playAgain_W(3, 198) <= 0; playAgain_W(3, 199) <= 0; playAgain_W(3, 200) <= 0; playAgain_W(3, 201) <= 0; playAgain_W(3, 202) <= 0; playAgain_W(3, 203) <= 0; playAgain_W(3, 204) <= 0; playAgain_W(3, 205) <= 0; playAgain_W(3, 206) <= 0; playAgain_W(3, 207) <= 0; playAgain_W(3, 208) <= 0; playAgain_W(3, 209) <= 0; playAgain_W(3, 210) <= 0; playAgain_W(3, 211) <= 0; playAgain_W(3, 212) <= 0; playAgain_W(3, 213) <= 0; playAgain_W(3, 214) <= 0; playAgain_W(3, 215) <= 0; playAgain_W(3, 216) <= 0; playAgain_W(3, 217) <= 0; playAgain_W(3, 218) <= 1; playAgain_W(3, 219) <= 1; playAgain_W(3, 220) <= 1; playAgain_W(3, 221) <= 1; playAgain_W(3, 222) <= 0; playAgain_W(3, 223) <= 0; playAgain_W(3, 224) <= 0; playAgain_W(3, 225) <= 0; playAgain_W(3, 226) <= 1; playAgain_W(3, 227) <= 1; playAgain_W(3, 228) <= 1; playAgain_W(3, 229) <= 1; playAgain_W(3, 230) <= 0; playAgain_W(3, 231) <= 0; playAgain_W(3, 232) <= 0; playAgain_W(3, 233) <= 0; playAgain_W(3, 234) <= 1; playAgain_W(3, 235) <= 1; playAgain_W(3, 236) <= 1; playAgain_W(3, 237) <= 1; playAgain_W(3, 238) <= 0; playAgain_W(3, 239) <= 0; playAgain_W(3, 240) <= 1; playAgain_W(3, 241) <= 1; playAgain_W(3, 242) <= 1; playAgain_W(3, 243) <= 1; playAgain_W(3, 244) <= 0; playAgain_W(3, 245) <= 0; playAgain_W(3, 246) <= 1; playAgain_W(3, 247) <= 1; playAgain_W(3, 248) <= 1; playAgain_W(3, 249) <= 1; playAgain_W(3, 250) <= 0; playAgain_W(3, 251) <= 0; playAgain_W(3, 252) <= 1; playAgain_W(3, 253) <= 1; playAgain_W(3, 254) <= 1; playAgain_W(3, 255) <= 1; playAgain_W(3, 256) <= 1; playAgain_W(3, 257) <= 1; playAgain_W(3, 258) <= 0; playAgain_W(3, 259) <= 0; playAgain_W(3, 260) <= 0; playAgain_W(3, 261) <= 0; playAgain_W(3, 262) <= 1; playAgain_W(3, 263) <= 1; playAgain_W(3, 264) <= 1; playAgain_W(3, 265) <= 1; playAgain_W(3, 266) <= 0; playAgain_W(3, 267) <= 0; playAgain_W(3, 268) <= 0; playAgain_W(3, 269) <= 0; playAgain_W(3, 270) <= 0; playAgain_W(3, 271) <= 0; playAgain_W(3, 272) <= 1; playAgain_W(3, 273) <= 1; playAgain_W(3, 274) <= 1; playAgain_W(3, 275) <= 1; playAgain_W(3, 276) <= 0; playAgain_W(3, 277) <= 0; playAgain_W(3, 278) <= 1; playAgain_W(3, 279) <= 1; playAgain_W(3, 280) <= 1; playAgain_W(3, 281) <= 1; playAgain_W(3, 282) <= 0; playAgain_W(3, 283) <= 0; playAgain_W(3, 284) <= 0; playAgain_W(3, 285) <= 0; playAgain_W(3, 286) <= 0; playAgain_W(3, 287) <= 0; 
playAgain_W(4, 0) <= 0; playAgain_W(4, 1) <= 0; playAgain_W(4, 2) <= 1; playAgain_W(4, 3) <= 1; playAgain_W(4, 4) <= 1; playAgain_W(4, 5) <= 1; playAgain_W(4, 6) <= 0; playAgain_W(4, 7) <= 0; playAgain_W(4, 8) <= 0; playAgain_W(4, 9) <= 0; playAgain_W(4, 10) <= 1; playAgain_W(4, 11) <= 1; playAgain_W(4, 12) <= 1; playAgain_W(4, 13) <= 1; playAgain_W(4, 14) <= 0; playAgain_W(4, 15) <= 0; playAgain_W(4, 16) <= 0; playAgain_W(4, 17) <= 0; playAgain_W(4, 18) <= 0; playAgain_W(4, 19) <= 0; playAgain_W(4, 20) <= 1; playAgain_W(4, 21) <= 1; playAgain_W(4, 22) <= 1; playAgain_W(4, 23) <= 1; playAgain_W(4, 24) <= 0; playAgain_W(4, 25) <= 0; playAgain_W(4, 26) <= 0; playAgain_W(4, 27) <= 0; playAgain_W(4, 28) <= 0; playAgain_W(4, 29) <= 0; playAgain_W(4, 30) <= 0; playAgain_W(4, 31) <= 0; playAgain_W(4, 32) <= 0; playAgain_W(4, 33) <= 0; playAgain_W(4, 34) <= 0; playAgain_W(4, 35) <= 0; playAgain_W(4, 36) <= 0; playAgain_W(4, 37) <= 0; playAgain_W(4, 38) <= 1; playAgain_W(4, 39) <= 1; playAgain_W(4, 40) <= 1; playAgain_W(4, 41) <= 1; playAgain_W(4, 42) <= 0; playAgain_W(4, 43) <= 0; playAgain_W(4, 44) <= 1; playAgain_W(4, 45) <= 1; playAgain_W(4, 46) <= 1; playAgain_W(4, 47) <= 1; playAgain_W(4, 48) <= 0; playAgain_W(4, 49) <= 0; playAgain_W(4, 50) <= 0; playAgain_W(4, 51) <= 0; playAgain_W(4, 52) <= 0; playAgain_W(4, 53) <= 0; playAgain_W(4, 54) <= 1; playAgain_W(4, 55) <= 1; playAgain_W(4, 56) <= 1; playAgain_W(4, 57) <= 1; playAgain_W(4, 58) <= 0; playAgain_W(4, 59) <= 0; playAgain_W(4, 60) <= 0; playAgain_W(4, 61) <= 0; playAgain_W(4, 62) <= 0; playAgain_W(4, 63) <= 0; playAgain_W(4, 64) <= 0; playAgain_W(4, 65) <= 0; playAgain_W(4, 66) <= 1; playAgain_W(4, 67) <= 1; playAgain_W(4, 68) <= 1; playAgain_W(4, 69) <= 1; playAgain_W(4, 70) <= 0; playAgain_W(4, 71) <= 0; playAgain_W(4, 72) <= 0; playAgain_W(4, 73) <= 0; playAgain_W(4, 74) <= 0; playAgain_W(4, 75) <= 0; playAgain_W(4, 76) <= 0; playAgain_W(4, 77) <= 0; playAgain_W(4, 78) <= 0; playAgain_W(4, 79) <= 0; playAgain_W(4, 80) <= 0; playAgain_W(4, 81) <= 0; playAgain_W(4, 82) <= 0; playAgain_W(4, 83) <= 0; playAgain_W(4, 84) <= 0; playAgain_W(4, 85) <= 0; playAgain_W(4, 86) <= 0; playAgain_W(4, 87) <= 0; playAgain_W(4, 88) <= 0; playAgain_W(4, 89) <= 0; playAgain_W(4, 90) <= 0; playAgain_W(4, 91) <= 0; playAgain_W(4, 92) <= 1; playAgain_W(4, 93) <= 1; playAgain_W(4, 94) <= 1; playAgain_W(4, 95) <= 1; playAgain_W(4, 96) <= 0; playAgain_W(4, 97) <= 0; playAgain_W(4, 98) <= 1; playAgain_W(4, 99) <= 1; playAgain_W(4, 100) <= 1; playAgain_W(4, 101) <= 1; playAgain_W(4, 102) <= 0; playAgain_W(4, 103) <= 0; playAgain_W(4, 104) <= 0; playAgain_W(4, 105) <= 0; playAgain_W(4, 106) <= 0; playAgain_W(4, 107) <= 0; playAgain_W(4, 108) <= 1; playAgain_W(4, 109) <= 1; playAgain_W(4, 110) <= 1; playAgain_W(4, 111) <= 1; playAgain_W(4, 112) <= 0; playAgain_W(4, 113) <= 0; playAgain_W(4, 114) <= 0; playAgain_W(4, 115) <= 0; playAgain_W(4, 116) <= 0; playAgain_W(4, 117) <= 0; playAgain_W(4, 118) <= 0; playAgain_W(4, 119) <= 0; playAgain_W(4, 120) <= 1; playAgain_W(4, 121) <= 1; playAgain_W(4, 122) <= 0; playAgain_W(4, 123) <= 0; playAgain_W(4, 124) <= 0; playAgain_W(4, 125) <= 0; playAgain_W(4, 126) <= 0; playAgain_W(4, 127) <= 0; playAgain_W(4, 128) <= 1; playAgain_W(4, 129) <= 1; playAgain_W(4, 130) <= 1; playAgain_W(4, 131) <= 1; playAgain_W(4, 132) <= 0; playAgain_W(4, 133) <= 0; playAgain_W(4, 134) <= 1; playAgain_W(4, 135) <= 1; playAgain_W(4, 136) <= 1; playAgain_W(4, 137) <= 1; playAgain_W(4, 138) <= 0; playAgain_W(4, 139) <= 0; playAgain_W(4, 140) <= 0; playAgain_W(4, 141) <= 0; playAgain_W(4, 142) <= 0; playAgain_W(4, 143) <= 0; playAgain_W(4, 144) <= 0; playAgain_W(4, 145) <= 0; playAgain_W(4, 146) <= 0; playAgain_W(4, 147) <= 0; playAgain_W(4, 148) <= 0; playAgain_W(4, 149) <= 0; playAgain_W(4, 150) <= 1; playAgain_W(4, 151) <= 1; playAgain_W(4, 152) <= 1; playAgain_W(4, 153) <= 1; playAgain_W(4, 154) <= 0; playAgain_W(4, 155) <= 0; playAgain_W(4, 156) <= 0; playAgain_W(4, 157) <= 0; playAgain_W(4, 158) <= 0; playAgain_W(4, 159) <= 0; playAgain_W(4, 160) <= 0; playAgain_W(4, 161) <= 0; playAgain_W(4, 162) <= 1; playAgain_W(4, 163) <= 1; playAgain_W(4, 164) <= 1; playAgain_W(4, 165) <= 1; playAgain_W(4, 166) <= 1; playAgain_W(4, 167) <= 1; playAgain_W(4, 168) <= 1; playAgain_W(4, 169) <= 1; playAgain_W(4, 170) <= 0; playAgain_W(4, 171) <= 0; playAgain_W(4, 172) <= 1; playAgain_W(4, 173) <= 1; playAgain_W(4, 174) <= 1; playAgain_W(4, 175) <= 1; playAgain_W(4, 176) <= 0; playAgain_W(4, 177) <= 0; playAgain_W(4, 178) <= 0; playAgain_W(4, 179) <= 0; playAgain_W(4, 180) <= 0; playAgain_W(4, 181) <= 0; playAgain_W(4, 182) <= 0; playAgain_W(4, 183) <= 0; playAgain_W(4, 184) <= 0; playAgain_W(4, 185) <= 0; playAgain_W(4, 186) <= 1; playAgain_W(4, 187) <= 1; playAgain_W(4, 188) <= 1; playAgain_W(4, 189) <= 1; playAgain_W(4, 190) <= 0; playAgain_W(4, 191) <= 0; playAgain_W(4, 192) <= 0; playAgain_W(4, 193) <= 0; playAgain_W(4, 194) <= 0; playAgain_W(4, 195) <= 0; playAgain_W(4, 196) <= 0; playAgain_W(4, 197) <= 0; playAgain_W(4, 198) <= 0; playAgain_W(4, 199) <= 0; playAgain_W(4, 200) <= 0; playAgain_W(4, 201) <= 0; playAgain_W(4, 202) <= 0; playAgain_W(4, 203) <= 0; playAgain_W(4, 204) <= 0; playAgain_W(4, 205) <= 0; playAgain_W(4, 206) <= 0; playAgain_W(4, 207) <= 0; playAgain_W(4, 208) <= 0; playAgain_W(4, 209) <= 0; playAgain_W(4, 210) <= 0; playAgain_W(4, 211) <= 0; playAgain_W(4, 212) <= 0; playAgain_W(4, 213) <= 0; playAgain_W(4, 214) <= 0; playAgain_W(4, 215) <= 0; playAgain_W(4, 216) <= 0; playAgain_W(4, 217) <= 0; playAgain_W(4, 218) <= 1; playAgain_W(4, 219) <= 1; playAgain_W(4, 220) <= 1; playAgain_W(4, 221) <= 1; playAgain_W(4, 222) <= 0; playAgain_W(4, 223) <= 0; playAgain_W(4, 224) <= 0; playAgain_W(4, 225) <= 0; playAgain_W(4, 226) <= 1; playAgain_W(4, 227) <= 1; playAgain_W(4, 228) <= 1; playAgain_W(4, 229) <= 1; playAgain_W(4, 230) <= 0; playAgain_W(4, 231) <= 0; playAgain_W(4, 232) <= 0; playAgain_W(4, 233) <= 0; playAgain_W(4, 234) <= 1; playAgain_W(4, 235) <= 1; playAgain_W(4, 236) <= 0; playAgain_W(4, 237) <= 0; playAgain_W(4, 238) <= 0; playAgain_W(4, 239) <= 0; playAgain_W(4, 240) <= 1; playAgain_W(4, 241) <= 1; playAgain_W(4, 242) <= 1; playAgain_W(4, 243) <= 1; playAgain_W(4, 244) <= 0; playAgain_W(4, 245) <= 0; playAgain_W(4, 246) <= 0; playAgain_W(4, 247) <= 0; playAgain_W(4, 248) <= 1; playAgain_W(4, 249) <= 1; playAgain_W(4, 250) <= 0; playAgain_W(4, 251) <= 0; playAgain_W(4, 252) <= 1; playAgain_W(4, 253) <= 1; playAgain_W(4, 254) <= 1; playAgain_W(4, 255) <= 1; playAgain_W(4, 256) <= 1; playAgain_W(4, 257) <= 1; playAgain_W(4, 258) <= 1; playAgain_W(4, 259) <= 1; playAgain_W(4, 260) <= 0; playAgain_W(4, 261) <= 0; playAgain_W(4, 262) <= 1; playAgain_W(4, 263) <= 1; playAgain_W(4, 264) <= 1; playAgain_W(4, 265) <= 1; playAgain_W(4, 266) <= 0; playAgain_W(4, 267) <= 0; playAgain_W(4, 268) <= 0; playAgain_W(4, 269) <= 0; playAgain_W(4, 270) <= 0; playAgain_W(4, 271) <= 0; playAgain_W(4, 272) <= 1; playAgain_W(4, 273) <= 1; playAgain_W(4, 274) <= 1; playAgain_W(4, 275) <= 1; playAgain_W(4, 276) <= 0; playAgain_W(4, 277) <= 0; playAgain_W(4, 278) <= 0; playAgain_W(4, 279) <= 0; playAgain_W(4, 280) <= 1; playAgain_W(4, 281) <= 1; playAgain_W(4, 282) <= 1; playAgain_W(4, 283) <= 1; playAgain_W(4, 284) <= 0; playAgain_W(4, 285) <= 0; playAgain_W(4, 286) <= 0; playAgain_W(4, 287) <= 0; 
playAgain_W(5, 0) <= 0; playAgain_W(5, 1) <= 0; playAgain_W(5, 2) <= 1; playAgain_W(5, 3) <= 1; playAgain_W(5, 4) <= 1; playAgain_W(5, 5) <= 1; playAgain_W(5, 6) <= 0; playAgain_W(5, 7) <= 0; playAgain_W(5, 8) <= 0; playAgain_W(5, 9) <= 0; playAgain_W(5, 10) <= 1; playAgain_W(5, 11) <= 1; playAgain_W(5, 12) <= 1; playAgain_W(5, 13) <= 1; playAgain_W(5, 14) <= 0; playAgain_W(5, 15) <= 0; playAgain_W(5, 16) <= 0; playAgain_W(5, 17) <= 0; playAgain_W(5, 18) <= 0; playAgain_W(5, 19) <= 0; playAgain_W(5, 20) <= 1; playAgain_W(5, 21) <= 1; playAgain_W(5, 22) <= 1; playAgain_W(5, 23) <= 1; playAgain_W(5, 24) <= 0; playAgain_W(5, 25) <= 0; playAgain_W(5, 26) <= 0; playAgain_W(5, 27) <= 0; playAgain_W(5, 28) <= 0; playAgain_W(5, 29) <= 0; playAgain_W(5, 30) <= 0; playAgain_W(5, 31) <= 0; playAgain_W(5, 32) <= 0; playAgain_W(5, 33) <= 0; playAgain_W(5, 34) <= 0; playAgain_W(5, 35) <= 0; playAgain_W(5, 36) <= 0; playAgain_W(5, 37) <= 0; playAgain_W(5, 38) <= 1; playAgain_W(5, 39) <= 1; playAgain_W(5, 40) <= 1; playAgain_W(5, 41) <= 1; playAgain_W(5, 42) <= 0; playAgain_W(5, 43) <= 0; playAgain_W(5, 44) <= 1; playAgain_W(5, 45) <= 1; playAgain_W(5, 46) <= 1; playAgain_W(5, 47) <= 1; playAgain_W(5, 48) <= 0; playAgain_W(5, 49) <= 0; playAgain_W(5, 50) <= 0; playAgain_W(5, 51) <= 0; playAgain_W(5, 52) <= 0; playAgain_W(5, 53) <= 0; playAgain_W(5, 54) <= 1; playAgain_W(5, 55) <= 1; playAgain_W(5, 56) <= 1; playAgain_W(5, 57) <= 1; playAgain_W(5, 58) <= 0; playAgain_W(5, 59) <= 0; playAgain_W(5, 60) <= 0; playAgain_W(5, 61) <= 0; playAgain_W(5, 62) <= 0; playAgain_W(5, 63) <= 0; playAgain_W(5, 64) <= 0; playAgain_W(5, 65) <= 0; playAgain_W(5, 66) <= 1; playAgain_W(5, 67) <= 1; playAgain_W(5, 68) <= 1; playAgain_W(5, 69) <= 1; playAgain_W(5, 70) <= 0; playAgain_W(5, 71) <= 0; playAgain_W(5, 72) <= 0; playAgain_W(5, 73) <= 0; playAgain_W(5, 74) <= 0; playAgain_W(5, 75) <= 0; playAgain_W(5, 76) <= 0; playAgain_W(5, 77) <= 0; playAgain_W(5, 78) <= 0; playAgain_W(5, 79) <= 0; playAgain_W(5, 80) <= 0; playAgain_W(5, 81) <= 0; playAgain_W(5, 82) <= 0; playAgain_W(5, 83) <= 0; playAgain_W(5, 84) <= 0; playAgain_W(5, 85) <= 0; playAgain_W(5, 86) <= 0; playAgain_W(5, 87) <= 0; playAgain_W(5, 88) <= 0; playAgain_W(5, 89) <= 0; playAgain_W(5, 90) <= 0; playAgain_W(5, 91) <= 0; playAgain_W(5, 92) <= 1; playAgain_W(5, 93) <= 1; playAgain_W(5, 94) <= 1; playAgain_W(5, 95) <= 1; playAgain_W(5, 96) <= 0; playAgain_W(5, 97) <= 0; playAgain_W(5, 98) <= 1; playAgain_W(5, 99) <= 1; playAgain_W(5, 100) <= 1; playAgain_W(5, 101) <= 1; playAgain_W(5, 102) <= 0; playAgain_W(5, 103) <= 0; playAgain_W(5, 104) <= 0; playAgain_W(5, 105) <= 0; playAgain_W(5, 106) <= 0; playAgain_W(5, 107) <= 0; playAgain_W(5, 108) <= 1; playAgain_W(5, 109) <= 1; playAgain_W(5, 110) <= 1; playAgain_W(5, 111) <= 1; playAgain_W(5, 112) <= 0; playAgain_W(5, 113) <= 0; playAgain_W(5, 114) <= 0; playAgain_W(5, 115) <= 0; playAgain_W(5, 116) <= 0; playAgain_W(5, 117) <= 0; playAgain_W(5, 118) <= 0; playAgain_W(5, 119) <= 0; playAgain_W(5, 120) <= 1; playAgain_W(5, 121) <= 1; playAgain_W(5, 122) <= 0; playAgain_W(5, 123) <= 0; playAgain_W(5, 124) <= 0; playAgain_W(5, 125) <= 0; playAgain_W(5, 126) <= 0; playAgain_W(5, 127) <= 0; playAgain_W(5, 128) <= 1; playAgain_W(5, 129) <= 1; playAgain_W(5, 130) <= 1; playAgain_W(5, 131) <= 1; playAgain_W(5, 132) <= 0; playAgain_W(5, 133) <= 0; playAgain_W(5, 134) <= 1; playAgain_W(5, 135) <= 1; playAgain_W(5, 136) <= 1; playAgain_W(5, 137) <= 1; playAgain_W(5, 138) <= 0; playAgain_W(5, 139) <= 0; playAgain_W(5, 140) <= 0; playAgain_W(5, 141) <= 0; playAgain_W(5, 142) <= 0; playAgain_W(5, 143) <= 0; playAgain_W(5, 144) <= 0; playAgain_W(5, 145) <= 0; playAgain_W(5, 146) <= 0; playAgain_W(5, 147) <= 0; playAgain_W(5, 148) <= 0; playAgain_W(5, 149) <= 0; playAgain_W(5, 150) <= 1; playAgain_W(5, 151) <= 1; playAgain_W(5, 152) <= 1; playAgain_W(5, 153) <= 1; playAgain_W(5, 154) <= 0; playAgain_W(5, 155) <= 0; playAgain_W(5, 156) <= 0; playAgain_W(5, 157) <= 0; playAgain_W(5, 158) <= 0; playAgain_W(5, 159) <= 0; playAgain_W(5, 160) <= 0; playAgain_W(5, 161) <= 0; playAgain_W(5, 162) <= 1; playAgain_W(5, 163) <= 1; playAgain_W(5, 164) <= 1; playAgain_W(5, 165) <= 1; playAgain_W(5, 166) <= 1; playAgain_W(5, 167) <= 1; playAgain_W(5, 168) <= 1; playAgain_W(5, 169) <= 1; playAgain_W(5, 170) <= 0; playAgain_W(5, 171) <= 0; playAgain_W(5, 172) <= 1; playAgain_W(5, 173) <= 1; playAgain_W(5, 174) <= 1; playAgain_W(5, 175) <= 1; playAgain_W(5, 176) <= 0; playAgain_W(5, 177) <= 0; playAgain_W(5, 178) <= 0; playAgain_W(5, 179) <= 0; playAgain_W(5, 180) <= 0; playAgain_W(5, 181) <= 0; playAgain_W(5, 182) <= 0; playAgain_W(5, 183) <= 0; playAgain_W(5, 184) <= 0; playAgain_W(5, 185) <= 0; playAgain_W(5, 186) <= 1; playAgain_W(5, 187) <= 1; playAgain_W(5, 188) <= 1; playAgain_W(5, 189) <= 1; playAgain_W(5, 190) <= 0; playAgain_W(5, 191) <= 0; playAgain_W(5, 192) <= 0; playAgain_W(5, 193) <= 0; playAgain_W(5, 194) <= 0; playAgain_W(5, 195) <= 0; playAgain_W(5, 196) <= 0; playAgain_W(5, 197) <= 0; playAgain_W(5, 198) <= 0; playAgain_W(5, 199) <= 0; playAgain_W(5, 200) <= 0; playAgain_W(5, 201) <= 0; playAgain_W(5, 202) <= 0; playAgain_W(5, 203) <= 0; playAgain_W(5, 204) <= 0; playAgain_W(5, 205) <= 0; playAgain_W(5, 206) <= 0; playAgain_W(5, 207) <= 0; playAgain_W(5, 208) <= 0; playAgain_W(5, 209) <= 0; playAgain_W(5, 210) <= 0; playAgain_W(5, 211) <= 0; playAgain_W(5, 212) <= 0; playAgain_W(5, 213) <= 0; playAgain_W(5, 214) <= 0; playAgain_W(5, 215) <= 0; playAgain_W(5, 216) <= 0; playAgain_W(5, 217) <= 0; playAgain_W(5, 218) <= 1; playAgain_W(5, 219) <= 1; playAgain_W(5, 220) <= 1; playAgain_W(5, 221) <= 1; playAgain_W(5, 222) <= 0; playAgain_W(5, 223) <= 0; playAgain_W(5, 224) <= 0; playAgain_W(5, 225) <= 0; playAgain_W(5, 226) <= 1; playAgain_W(5, 227) <= 1; playAgain_W(5, 228) <= 1; playAgain_W(5, 229) <= 1; playAgain_W(5, 230) <= 0; playAgain_W(5, 231) <= 0; playAgain_W(5, 232) <= 0; playAgain_W(5, 233) <= 0; playAgain_W(5, 234) <= 1; playAgain_W(5, 235) <= 1; playAgain_W(5, 236) <= 0; playAgain_W(5, 237) <= 0; playAgain_W(5, 238) <= 0; playAgain_W(5, 239) <= 0; playAgain_W(5, 240) <= 1; playAgain_W(5, 241) <= 1; playAgain_W(5, 242) <= 1; playAgain_W(5, 243) <= 1; playAgain_W(5, 244) <= 0; playAgain_W(5, 245) <= 0; playAgain_W(5, 246) <= 0; playAgain_W(5, 247) <= 0; playAgain_W(5, 248) <= 1; playAgain_W(5, 249) <= 1; playAgain_W(5, 250) <= 0; playAgain_W(5, 251) <= 0; playAgain_W(5, 252) <= 1; playAgain_W(5, 253) <= 1; playAgain_W(5, 254) <= 1; playAgain_W(5, 255) <= 1; playAgain_W(5, 256) <= 1; playAgain_W(5, 257) <= 1; playAgain_W(5, 258) <= 1; playAgain_W(5, 259) <= 1; playAgain_W(5, 260) <= 0; playAgain_W(5, 261) <= 0; playAgain_W(5, 262) <= 1; playAgain_W(5, 263) <= 1; playAgain_W(5, 264) <= 1; playAgain_W(5, 265) <= 1; playAgain_W(5, 266) <= 0; playAgain_W(5, 267) <= 0; playAgain_W(5, 268) <= 0; playAgain_W(5, 269) <= 0; playAgain_W(5, 270) <= 0; playAgain_W(5, 271) <= 0; playAgain_W(5, 272) <= 1; playAgain_W(5, 273) <= 1; playAgain_W(5, 274) <= 1; playAgain_W(5, 275) <= 1; playAgain_W(5, 276) <= 0; playAgain_W(5, 277) <= 0; playAgain_W(5, 278) <= 0; playAgain_W(5, 279) <= 0; playAgain_W(5, 280) <= 1; playAgain_W(5, 281) <= 1; playAgain_W(5, 282) <= 1; playAgain_W(5, 283) <= 1; playAgain_W(5, 284) <= 0; playAgain_W(5, 285) <= 0; playAgain_W(5, 286) <= 0; playAgain_W(5, 287) <= 0; 
playAgain_W(6, 0) <= 0; playAgain_W(6, 1) <= 0; playAgain_W(6, 2) <= 1; playAgain_W(6, 3) <= 1; playAgain_W(6, 4) <= 1; playAgain_W(6, 5) <= 1; playAgain_W(6, 6) <= 0; playAgain_W(6, 7) <= 0; playAgain_W(6, 8) <= 0; playAgain_W(6, 9) <= 0; playAgain_W(6, 10) <= 1; playAgain_W(6, 11) <= 1; playAgain_W(6, 12) <= 1; playAgain_W(6, 13) <= 1; playAgain_W(6, 14) <= 0; playAgain_W(6, 15) <= 0; playAgain_W(6, 16) <= 0; playAgain_W(6, 17) <= 0; playAgain_W(6, 18) <= 0; playAgain_W(6, 19) <= 0; playAgain_W(6, 20) <= 1; playAgain_W(6, 21) <= 1; playAgain_W(6, 22) <= 1; playAgain_W(6, 23) <= 1; playAgain_W(6, 24) <= 0; playAgain_W(6, 25) <= 0; playAgain_W(6, 26) <= 0; playAgain_W(6, 27) <= 0; playAgain_W(6, 28) <= 0; playAgain_W(6, 29) <= 0; playAgain_W(6, 30) <= 0; playAgain_W(6, 31) <= 0; playAgain_W(6, 32) <= 0; playAgain_W(6, 33) <= 0; playAgain_W(6, 34) <= 0; playAgain_W(6, 35) <= 0; playAgain_W(6, 36) <= 1; playAgain_W(6, 37) <= 1; playAgain_W(6, 38) <= 1; playAgain_W(6, 39) <= 1; playAgain_W(6, 40) <= 0; playAgain_W(6, 41) <= 0; playAgain_W(6, 42) <= 0; playAgain_W(6, 43) <= 0; playAgain_W(6, 44) <= 0; playAgain_W(6, 45) <= 0; playAgain_W(6, 46) <= 1; playAgain_W(6, 47) <= 1; playAgain_W(6, 48) <= 1; playAgain_W(6, 49) <= 1; playAgain_W(6, 50) <= 0; playAgain_W(6, 51) <= 0; playAgain_W(6, 52) <= 0; playAgain_W(6, 53) <= 0; playAgain_W(6, 54) <= 0; playAgain_W(6, 55) <= 0; playAgain_W(6, 56) <= 1; playAgain_W(6, 57) <= 1; playAgain_W(6, 58) <= 1; playAgain_W(6, 59) <= 1; playAgain_W(6, 60) <= 0; playAgain_W(6, 61) <= 0; playAgain_W(6, 62) <= 0; playAgain_W(6, 63) <= 0; playAgain_W(6, 64) <= 1; playAgain_W(6, 65) <= 1; playAgain_W(6, 66) <= 1; playAgain_W(6, 67) <= 1; playAgain_W(6, 68) <= 0; playAgain_W(6, 69) <= 0; playAgain_W(6, 70) <= 0; playAgain_W(6, 71) <= 0; playAgain_W(6, 72) <= 0; playAgain_W(6, 73) <= 0; playAgain_W(6, 74) <= 0; playAgain_W(6, 75) <= 0; playAgain_W(6, 76) <= 0; playAgain_W(6, 77) <= 0; playAgain_W(6, 78) <= 0; playAgain_W(6, 79) <= 0; playAgain_W(6, 80) <= 0; playAgain_W(6, 81) <= 0; playAgain_W(6, 82) <= 0; playAgain_W(6, 83) <= 0; playAgain_W(6, 84) <= 0; playAgain_W(6, 85) <= 0; playAgain_W(6, 86) <= 0; playAgain_W(6, 87) <= 0; playAgain_W(6, 88) <= 0; playAgain_W(6, 89) <= 0; playAgain_W(6, 90) <= 1; playAgain_W(6, 91) <= 1; playAgain_W(6, 92) <= 1; playAgain_W(6, 93) <= 1; playAgain_W(6, 94) <= 0; playAgain_W(6, 95) <= 0; playAgain_W(6, 96) <= 0; playAgain_W(6, 97) <= 0; playAgain_W(6, 98) <= 0; playAgain_W(6, 99) <= 0; playAgain_W(6, 100) <= 1; playAgain_W(6, 101) <= 1; playAgain_W(6, 102) <= 1; playAgain_W(6, 103) <= 1; playAgain_W(6, 104) <= 0; playAgain_W(6, 105) <= 0; playAgain_W(6, 106) <= 0; playAgain_W(6, 107) <= 0; playAgain_W(6, 108) <= 1; playAgain_W(6, 109) <= 1; playAgain_W(6, 110) <= 1; playAgain_W(6, 111) <= 1; playAgain_W(6, 112) <= 0; playAgain_W(6, 113) <= 0; playAgain_W(6, 114) <= 0; playAgain_W(6, 115) <= 0; playAgain_W(6, 116) <= 0; playAgain_W(6, 117) <= 0; playAgain_W(6, 118) <= 0; playAgain_W(6, 119) <= 0; playAgain_W(6, 120) <= 0; playAgain_W(6, 121) <= 0; playAgain_W(6, 122) <= 0; playAgain_W(6, 123) <= 0; playAgain_W(6, 124) <= 0; playAgain_W(6, 125) <= 0; playAgain_W(6, 126) <= 1; playAgain_W(6, 127) <= 1; playAgain_W(6, 128) <= 1; playAgain_W(6, 129) <= 1; playAgain_W(6, 130) <= 0; playAgain_W(6, 131) <= 0; playAgain_W(6, 132) <= 0; playAgain_W(6, 133) <= 0; playAgain_W(6, 134) <= 0; playAgain_W(6, 135) <= 0; playAgain_W(6, 136) <= 1; playAgain_W(6, 137) <= 1; playAgain_W(6, 138) <= 1; playAgain_W(6, 139) <= 1; playAgain_W(6, 140) <= 0; playAgain_W(6, 141) <= 0; playAgain_W(6, 142) <= 0; playAgain_W(6, 143) <= 0; playAgain_W(6, 144) <= 0; playAgain_W(6, 145) <= 0; playAgain_W(6, 146) <= 0; playAgain_W(6, 147) <= 0; playAgain_W(6, 148) <= 0; playAgain_W(6, 149) <= 0; playAgain_W(6, 150) <= 1; playAgain_W(6, 151) <= 1; playAgain_W(6, 152) <= 1; playAgain_W(6, 153) <= 1; playAgain_W(6, 154) <= 0; playAgain_W(6, 155) <= 0; playAgain_W(6, 156) <= 0; playAgain_W(6, 157) <= 0; playAgain_W(6, 158) <= 0; playAgain_W(6, 159) <= 0; playAgain_W(6, 160) <= 0; playAgain_W(6, 161) <= 0; playAgain_W(6, 162) <= 1; playAgain_W(6, 163) <= 1; playAgain_W(6, 164) <= 1; playAgain_W(6, 165) <= 1; playAgain_W(6, 166) <= 1; playAgain_W(6, 167) <= 1; playAgain_W(6, 168) <= 1; playAgain_W(6, 169) <= 1; playAgain_W(6, 170) <= 1; playAgain_W(6, 171) <= 1; playAgain_W(6, 172) <= 1; playAgain_W(6, 173) <= 1; playAgain_W(6, 174) <= 1; playAgain_W(6, 175) <= 1; playAgain_W(6, 176) <= 0; playAgain_W(6, 177) <= 0; playAgain_W(6, 178) <= 0; playAgain_W(6, 179) <= 0; playAgain_W(6, 180) <= 0; playAgain_W(6, 181) <= 0; playAgain_W(6, 182) <= 0; playAgain_W(6, 183) <= 0; playAgain_W(6, 184) <= 0; playAgain_W(6, 185) <= 0; playAgain_W(6, 186) <= 1; playAgain_W(6, 187) <= 1; playAgain_W(6, 188) <= 1; playAgain_W(6, 189) <= 1; playAgain_W(6, 190) <= 0; playAgain_W(6, 191) <= 0; playAgain_W(6, 192) <= 0; playAgain_W(6, 193) <= 0; playAgain_W(6, 194) <= 0; playAgain_W(6, 195) <= 0; playAgain_W(6, 196) <= 0; playAgain_W(6, 197) <= 0; playAgain_W(6, 198) <= 0; playAgain_W(6, 199) <= 0; playAgain_W(6, 200) <= 0; playAgain_W(6, 201) <= 0; playAgain_W(6, 202) <= 0; playAgain_W(6, 203) <= 0; playAgain_W(6, 204) <= 0; playAgain_W(6, 205) <= 0; playAgain_W(6, 206) <= 0; playAgain_W(6, 207) <= 0; playAgain_W(6, 208) <= 0; playAgain_W(6, 209) <= 0; playAgain_W(6, 210) <= 0; playAgain_W(6, 211) <= 0; playAgain_W(6, 212) <= 0; playAgain_W(6, 213) <= 0; playAgain_W(6, 214) <= 0; playAgain_W(6, 215) <= 0; playAgain_W(6, 216) <= 0; playAgain_W(6, 217) <= 0; playAgain_W(6, 218) <= 1; playAgain_W(6, 219) <= 1; playAgain_W(6, 220) <= 1; playAgain_W(6, 221) <= 1; playAgain_W(6, 222) <= 0; playAgain_W(6, 223) <= 0; playAgain_W(6, 224) <= 0; playAgain_W(6, 225) <= 0; playAgain_W(6, 226) <= 1; playAgain_W(6, 227) <= 1; playAgain_W(6, 228) <= 1; playAgain_W(6, 229) <= 1; playAgain_W(6, 230) <= 0; playAgain_W(6, 231) <= 0; playAgain_W(6, 232) <= 0; playAgain_W(6, 233) <= 0; playAgain_W(6, 234) <= 0; playAgain_W(6, 235) <= 0; playAgain_W(6, 236) <= 0; playAgain_W(6, 237) <= 0; playAgain_W(6, 238) <= 0; playAgain_W(6, 239) <= 0; playAgain_W(6, 240) <= 1; playAgain_W(6, 241) <= 1; playAgain_W(6, 242) <= 1; playAgain_W(6, 243) <= 1; playAgain_W(6, 244) <= 0; playAgain_W(6, 245) <= 0; playAgain_W(6, 246) <= 0; playAgain_W(6, 247) <= 0; playAgain_W(6, 248) <= 0; playAgain_W(6, 249) <= 0; playAgain_W(6, 250) <= 0; playAgain_W(6, 251) <= 0; playAgain_W(6, 252) <= 1; playAgain_W(6, 253) <= 1; playAgain_W(6, 254) <= 1; playAgain_W(6, 255) <= 1; playAgain_W(6, 256) <= 1; playAgain_W(6, 257) <= 1; playAgain_W(6, 258) <= 1; playAgain_W(6, 259) <= 1; playAgain_W(6, 260) <= 1; playAgain_W(6, 261) <= 1; playAgain_W(6, 262) <= 1; playAgain_W(6, 263) <= 1; playAgain_W(6, 264) <= 1; playAgain_W(6, 265) <= 1; playAgain_W(6, 266) <= 0; playAgain_W(6, 267) <= 0; playAgain_W(6, 268) <= 0; playAgain_W(6, 269) <= 0; playAgain_W(6, 270) <= 0; playAgain_W(6, 271) <= 0; playAgain_W(6, 272) <= 1; playAgain_W(6, 273) <= 1; playAgain_W(6, 274) <= 1; playAgain_W(6, 275) <= 1; playAgain_W(6, 276) <= 0; playAgain_W(6, 277) <= 0; playAgain_W(6, 278) <= 0; playAgain_W(6, 279) <= 0; playAgain_W(6, 280) <= 1; playAgain_W(6, 281) <= 1; playAgain_W(6, 282) <= 1; playAgain_W(6, 283) <= 1; playAgain_W(6, 284) <= 0; playAgain_W(6, 285) <= 0; playAgain_W(6, 286) <= 0; playAgain_W(6, 287) <= 0; 
playAgain_W(7, 0) <= 0; playAgain_W(7, 1) <= 0; playAgain_W(7, 2) <= 1; playAgain_W(7, 3) <= 1; playAgain_W(7, 4) <= 1; playAgain_W(7, 5) <= 1; playAgain_W(7, 6) <= 0; playAgain_W(7, 7) <= 0; playAgain_W(7, 8) <= 0; playAgain_W(7, 9) <= 0; playAgain_W(7, 10) <= 1; playAgain_W(7, 11) <= 1; playAgain_W(7, 12) <= 1; playAgain_W(7, 13) <= 1; playAgain_W(7, 14) <= 0; playAgain_W(7, 15) <= 0; playAgain_W(7, 16) <= 0; playAgain_W(7, 17) <= 0; playAgain_W(7, 18) <= 0; playAgain_W(7, 19) <= 0; playAgain_W(7, 20) <= 1; playAgain_W(7, 21) <= 1; playAgain_W(7, 22) <= 1; playAgain_W(7, 23) <= 1; playAgain_W(7, 24) <= 0; playAgain_W(7, 25) <= 0; playAgain_W(7, 26) <= 0; playAgain_W(7, 27) <= 0; playAgain_W(7, 28) <= 0; playAgain_W(7, 29) <= 0; playAgain_W(7, 30) <= 0; playAgain_W(7, 31) <= 0; playAgain_W(7, 32) <= 0; playAgain_W(7, 33) <= 0; playAgain_W(7, 34) <= 0; playAgain_W(7, 35) <= 0; playAgain_W(7, 36) <= 1; playAgain_W(7, 37) <= 1; playAgain_W(7, 38) <= 1; playAgain_W(7, 39) <= 1; playAgain_W(7, 40) <= 0; playAgain_W(7, 41) <= 0; playAgain_W(7, 42) <= 0; playAgain_W(7, 43) <= 0; playAgain_W(7, 44) <= 0; playAgain_W(7, 45) <= 0; playAgain_W(7, 46) <= 1; playAgain_W(7, 47) <= 1; playAgain_W(7, 48) <= 1; playAgain_W(7, 49) <= 1; playAgain_W(7, 50) <= 0; playAgain_W(7, 51) <= 0; playAgain_W(7, 52) <= 0; playAgain_W(7, 53) <= 0; playAgain_W(7, 54) <= 0; playAgain_W(7, 55) <= 0; playAgain_W(7, 56) <= 1; playAgain_W(7, 57) <= 1; playAgain_W(7, 58) <= 1; playAgain_W(7, 59) <= 1; playAgain_W(7, 60) <= 0; playAgain_W(7, 61) <= 0; playAgain_W(7, 62) <= 0; playAgain_W(7, 63) <= 0; playAgain_W(7, 64) <= 1; playAgain_W(7, 65) <= 1; playAgain_W(7, 66) <= 1; playAgain_W(7, 67) <= 1; playAgain_W(7, 68) <= 0; playAgain_W(7, 69) <= 0; playAgain_W(7, 70) <= 0; playAgain_W(7, 71) <= 0; playAgain_W(7, 72) <= 0; playAgain_W(7, 73) <= 0; playAgain_W(7, 74) <= 0; playAgain_W(7, 75) <= 0; playAgain_W(7, 76) <= 0; playAgain_W(7, 77) <= 0; playAgain_W(7, 78) <= 0; playAgain_W(7, 79) <= 0; playAgain_W(7, 80) <= 0; playAgain_W(7, 81) <= 0; playAgain_W(7, 82) <= 0; playAgain_W(7, 83) <= 0; playAgain_W(7, 84) <= 0; playAgain_W(7, 85) <= 0; playAgain_W(7, 86) <= 0; playAgain_W(7, 87) <= 0; playAgain_W(7, 88) <= 0; playAgain_W(7, 89) <= 0; playAgain_W(7, 90) <= 1; playAgain_W(7, 91) <= 1; playAgain_W(7, 92) <= 1; playAgain_W(7, 93) <= 1; playAgain_W(7, 94) <= 0; playAgain_W(7, 95) <= 0; playAgain_W(7, 96) <= 0; playAgain_W(7, 97) <= 0; playAgain_W(7, 98) <= 0; playAgain_W(7, 99) <= 0; playAgain_W(7, 100) <= 1; playAgain_W(7, 101) <= 1; playAgain_W(7, 102) <= 1; playAgain_W(7, 103) <= 1; playAgain_W(7, 104) <= 0; playAgain_W(7, 105) <= 0; playAgain_W(7, 106) <= 0; playAgain_W(7, 107) <= 0; playAgain_W(7, 108) <= 1; playAgain_W(7, 109) <= 1; playAgain_W(7, 110) <= 1; playAgain_W(7, 111) <= 1; playAgain_W(7, 112) <= 0; playAgain_W(7, 113) <= 0; playAgain_W(7, 114) <= 0; playAgain_W(7, 115) <= 0; playAgain_W(7, 116) <= 0; playAgain_W(7, 117) <= 0; playAgain_W(7, 118) <= 0; playAgain_W(7, 119) <= 0; playAgain_W(7, 120) <= 0; playAgain_W(7, 121) <= 0; playAgain_W(7, 122) <= 0; playAgain_W(7, 123) <= 0; playAgain_W(7, 124) <= 0; playAgain_W(7, 125) <= 0; playAgain_W(7, 126) <= 1; playAgain_W(7, 127) <= 1; playAgain_W(7, 128) <= 1; playAgain_W(7, 129) <= 1; playAgain_W(7, 130) <= 0; playAgain_W(7, 131) <= 0; playAgain_W(7, 132) <= 0; playAgain_W(7, 133) <= 0; playAgain_W(7, 134) <= 0; playAgain_W(7, 135) <= 0; playAgain_W(7, 136) <= 1; playAgain_W(7, 137) <= 1; playAgain_W(7, 138) <= 1; playAgain_W(7, 139) <= 1; playAgain_W(7, 140) <= 0; playAgain_W(7, 141) <= 0; playAgain_W(7, 142) <= 0; playAgain_W(7, 143) <= 0; playAgain_W(7, 144) <= 0; playAgain_W(7, 145) <= 0; playAgain_W(7, 146) <= 0; playAgain_W(7, 147) <= 0; playAgain_W(7, 148) <= 0; playAgain_W(7, 149) <= 0; playAgain_W(7, 150) <= 1; playAgain_W(7, 151) <= 1; playAgain_W(7, 152) <= 1; playAgain_W(7, 153) <= 1; playAgain_W(7, 154) <= 0; playAgain_W(7, 155) <= 0; playAgain_W(7, 156) <= 0; playAgain_W(7, 157) <= 0; playAgain_W(7, 158) <= 0; playAgain_W(7, 159) <= 0; playAgain_W(7, 160) <= 0; playAgain_W(7, 161) <= 0; playAgain_W(7, 162) <= 1; playAgain_W(7, 163) <= 1; playAgain_W(7, 164) <= 1; playAgain_W(7, 165) <= 1; playAgain_W(7, 166) <= 1; playAgain_W(7, 167) <= 1; playAgain_W(7, 168) <= 1; playAgain_W(7, 169) <= 1; playAgain_W(7, 170) <= 1; playAgain_W(7, 171) <= 1; playAgain_W(7, 172) <= 1; playAgain_W(7, 173) <= 1; playAgain_W(7, 174) <= 1; playAgain_W(7, 175) <= 1; playAgain_W(7, 176) <= 0; playAgain_W(7, 177) <= 0; playAgain_W(7, 178) <= 0; playAgain_W(7, 179) <= 0; playAgain_W(7, 180) <= 0; playAgain_W(7, 181) <= 0; playAgain_W(7, 182) <= 0; playAgain_W(7, 183) <= 0; playAgain_W(7, 184) <= 0; playAgain_W(7, 185) <= 0; playAgain_W(7, 186) <= 1; playAgain_W(7, 187) <= 1; playAgain_W(7, 188) <= 1; playAgain_W(7, 189) <= 1; playAgain_W(7, 190) <= 0; playAgain_W(7, 191) <= 0; playAgain_W(7, 192) <= 0; playAgain_W(7, 193) <= 0; playAgain_W(7, 194) <= 0; playAgain_W(7, 195) <= 0; playAgain_W(7, 196) <= 0; playAgain_W(7, 197) <= 0; playAgain_W(7, 198) <= 0; playAgain_W(7, 199) <= 0; playAgain_W(7, 200) <= 0; playAgain_W(7, 201) <= 0; playAgain_W(7, 202) <= 0; playAgain_W(7, 203) <= 0; playAgain_W(7, 204) <= 0; playAgain_W(7, 205) <= 0; playAgain_W(7, 206) <= 0; playAgain_W(7, 207) <= 0; playAgain_W(7, 208) <= 0; playAgain_W(7, 209) <= 0; playAgain_W(7, 210) <= 0; playAgain_W(7, 211) <= 0; playAgain_W(7, 212) <= 0; playAgain_W(7, 213) <= 0; playAgain_W(7, 214) <= 0; playAgain_W(7, 215) <= 0; playAgain_W(7, 216) <= 0; playAgain_W(7, 217) <= 0; playAgain_W(7, 218) <= 1; playAgain_W(7, 219) <= 1; playAgain_W(7, 220) <= 1; playAgain_W(7, 221) <= 1; playAgain_W(7, 222) <= 0; playAgain_W(7, 223) <= 0; playAgain_W(7, 224) <= 0; playAgain_W(7, 225) <= 0; playAgain_W(7, 226) <= 1; playAgain_W(7, 227) <= 1; playAgain_W(7, 228) <= 1; playAgain_W(7, 229) <= 1; playAgain_W(7, 230) <= 0; playAgain_W(7, 231) <= 0; playAgain_W(7, 232) <= 0; playAgain_W(7, 233) <= 0; playAgain_W(7, 234) <= 0; playAgain_W(7, 235) <= 0; playAgain_W(7, 236) <= 0; playAgain_W(7, 237) <= 0; playAgain_W(7, 238) <= 0; playAgain_W(7, 239) <= 0; playAgain_W(7, 240) <= 1; playAgain_W(7, 241) <= 1; playAgain_W(7, 242) <= 1; playAgain_W(7, 243) <= 1; playAgain_W(7, 244) <= 0; playAgain_W(7, 245) <= 0; playAgain_W(7, 246) <= 0; playAgain_W(7, 247) <= 0; playAgain_W(7, 248) <= 0; playAgain_W(7, 249) <= 0; playAgain_W(7, 250) <= 0; playAgain_W(7, 251) <= 0; playAgain_W(7, 252) <= 1; playAgain_W(7, 253) <= 1; playAgain_W(7, 254) <= 1; playAgain_W(7, 255) <= 1; playAgain_W(7, 256) <= 1; playAgain_W(7, 257) <= 1; playAgain_W(7, 258) <= 1; playAgain_W(7, 259) <= 1; playAgain_W(7, 260) <= 1; playAgain_W(7, 261) <= 1; playAgain_W(7, 262) <= 1; playAgain_W(7, 263) <= 1; playAgain_W(7, 264) <= 1; playAgain_W(7, 265) <= 1; playAgain_W(7, 266) <= 0; playAgain_W(7, 267) <= 0; playAgain_W(7, 268) <= 0; playAgain_W(7, 269) <= 0; playAgain_W(7, 270) <= 0; playAgain_W(7, 271) <= 0; playAgain_W(7, 272) <= 1; playAgain_W(7, 273) <= 1; playAgain_W(7, 274) <= 1; playAgain_W(7, 275) <= 1; playAgain_W(7, 276) <= 0; playAgain_W(7, 277) <= 0; playAgain_W(7, 278) <= 0; playAgain_W(7, 279) <= 0; playAgain_W(7, 280) <= 1; playAgain_W(7, 281) <= 1; playAgain_W(7, 282) <= 1; playAgain_W(7, 283) <= 1; playAgain_W(7, 284) <= 0; playAgain_W(7, 285) <= 0; playAgain_W(7, 286) <= 0; playAgain_W(7, 287) <= 0; 
playAgain_W(8, 0) <= 0; playAgain_W(8, 1) <= 0; playAgain_W(8, 2) <= 1; playAgain_W(8, 3) <= 1; playAgain_W(8, 4) <= 1; playAgain_W(8, 5) <= 1; playAgain_W(8, 6) <= 1; playAgain_W(8, 7) <= 1; playAgain_W(8, 8) <= 1; playAgain_W(8, 9) <= 1; playAgain_W(8, 10) <= 1; playAgain_W(8, 11) <= 1; playAgain_W(8, 12) <= 0; playAgain_W(8, 13) <= 0; playAgain_W(8, 14) <= 0; playAgain_W(8, 15) <= 0; playAgain_W(8, 16) <= 0; playAgain_W(8, 17) <= 0; playAgain_W(8, 18) <= 0; playAgain_W(8, 19) <= 0; playAgain_W(8, 20) <= 1; playAgain_W(8, 21) <= 1; playAgain_W(8, 22) <= 1; playAgain_W(8, 23) <= 1; playAgain_W(8, 24) <= 0; playAgain_W(8, 25) <= 0; playAgain_W(8, 26) <= 0; playAgain_W(8, 27) <= 0; playAgain_W(8, 28) <= 0; playAgain_W(8, 29) <= 0; playAgain_W(8, 30) <= 0; playAgain_W(8, 31) <= 0; playAgain_W(8, 32) <= 0; playAgain_W(8, 33) <= 0; playAgain_W(8, 34) <= 0; playAgain_W(8, 35) <= 0; playAgain_W(8, 36) <= 1; playAgain_W(8, 37) <= 1; playAgain_W(8, 38) <= 1; playAgain_W(8, 39) <= 1; playAgain_W(8, 40) <= 0; playAgain_W(8, 41) <= 0; playAgain_W(8, 42) <= 0; playAgain_W(8, 43) <= 0; playAgain_W(8, 44) <= 0; playAgain_W(8, 45) <= 0; playAgain_W(8, 46) <= 1; playAgain_W(8, 47) <= 1; playAgain_W(8, 48) <= 1; playAgain_W(8, 49) <= 1; playAgain_W(8, 50) <= 0; playAgain_W(8, 51) <= 0; playAgain_W(8, 52) <= 0; playAgain_W(8, 53) <= 0; playAgain_W(8, 54) <= 0; playAgain_W(8, 55) <= 0; playAgain_W(8, 56) <= 0; playAgain_W(8, 57) <= 0; playAgain_W(8, 58) <= 1; playAgain_W(8, 59) <= 1; playAgain_W(8, 60) <= 1; playAgain_W(8, 61) <= 1; playAgain_W(8, 62) <= 1; playAgain_W(8, 63) <= 1; playAgain_W(8, 64) <= 1; playAgain_W(8, 65) <= 1; playAgain_W(8, 66) <= 0; playAgain_W(8, 67) <= 0; playAgain_W(8, 68) <= 0; playAgain_W(8, 69) <= 0; playAgain_W(8, 70) <= 0; playAgain_W(8, 71) <= 0; playAgain_W(8, 72) <= 0; playAgain_W(8, 73) <= 0; playAgain_W(8, 74) <= 0; playAgain_W(8, 75) <= 0; playAgain_W(8, 76) <= 0; playAgain_W(8, 77) <= 0; playAgain_W(8, 78) <= 0; playAgain_W(8, 79) <= 0; playAgain_W(8, 80) <= 0; playAgain_W(8, 81) <= 0; playAgain_W(8, 82) <= 0; playAgain_W(8, 83) <= 0; playAgain_W(8, 84) <= 0; playAgain_W(8, 85) <= 0; playAgain_W(8, 86) <= 0; playAgain_W(8, 87) <= 0; playAgain_W(8, 88) <= 0; playAgain_W(8, 89) <= 0; playAgain_W(8, 90) <= 1; playAgain_W(8, 91) <= 1; playAgain_W(8, 92) <= 1; playAgain_W(8, 93) <= 1; playAgain_W(8, 94) <= 0; playAgain_W(8, 95) <= 0; playAgain_W(8, 96) <= 0; playAgain_W(8, 97) <= 0; playAgain_W(8, 98) <= 0; playAgain_W(8, 99) <= 0; playAgain_W(8, 100) <= 1; playAgain_W(8, 101) <= 1; playAgain_W(8, 102) <= 1; playAgain_W(8, 103) <= 1; playAgain_W(8, 104) <= 0; playAgain_W(8, 105) <= 0; playAgain_W(8, 106) <= 0; playAgain_W(8, 107) <= 0; playAgain_W(8, 108) <= 1; playAgain_W(8, 109) <= 1; playAgain_W(8, 110) <= 1; playAgain_W(8, 111) <= 1; playAgain_W(8, 112) <= 0; playAgain_W(8, 113) <= 0; playAgain_W(8, 114) <= 0; playAgain_W(8, 115) <= 0; playAgain_W(8, 116) <= 0; playAgain_W(8, 117) <= 0; playAgain_W(8, 118) <= 0; playAgain_W(8, 119) <= 0; playAgain_W(8, 120) <= 0; playAgain_W(8, 121) <= 0; playAgain_W(8, 122) <= 0; playAgain_W(8, 123) <= 0; playAgain_W(8, 124) <= 0; playAgain_W(8, 125) <= 0; playAgain_W(8, 126) <= 1; playAgain_W(8, 127) <= 1; playAgain_W(8, 128) <= 1; playAgain_W(8, 129) <= 1; playAgain_W(8, 130) <= 0; playAgain_W(8, 131) <= 0; playAgain_W(8, 132) <= 0; playAgain_W(8, 133) <= 0; playAgain_W(8, 134) <= 0; playAgain_W(8, 135) <= 0; playAgain_W(8, 136) <= 1; playAgain_W(8, 137) <= 1; playAgain_W(8, 138) <= 1; playAgain_W(8, 139) <= 1; playAgain_W(8, 140) <= 0; playAgain_W(8, 141) <= 0; playAgain_W(8, 142) <= 0; playAgain_W(8, 143) <= 0; playAgain_W(8, 144) <= 0; playAgain_W(8, 145) <= 0; playAgain_W(8, 146) <= 0; playAgain_W(8, 147) <= 0; playAgain_W(8, 148) <= 0; playAgain_W(8, 149) <= 0; playAgain_W(8, 150) <= 1; playAgain_W(8, 151) <= 1; playAgain_W(8, 152) <= 1; playAgain_W(8, 153) <= 1; playAgain_W(8, 154) <= 0; playAgain_W(8, 155) <= 0; playAgain_W(8, 156) <= 0; playAgain_W(8, 157) <= 0; playAgain_W(8, 158) <= 0; playAgain_W(8, 159) <= 0; playAgain_W(8, 160) <= 0; playAgain_W(8, 161) <= 0; playAgain_W(8, 162) <= 1; playAgain_W(8, 163) <= 1; playAgain_W(8, 164) <= 1; playAgain_W(8, 165) <= 1; playAgain_W(8, 166) <= 0; playAgain_W(8, 167) <= 0; playAgain_W(8, 168) <= 1; playAgain_W(8, 169) <= 1; playAgain_W(8, 170) <= 1; playAgain_W(8, 171) <= 1; playAgain_W(8, 172) <= 1; playAgain_W(8, 173) <= 1; playAgain_W(8, 174) <= 1; playAgain_W(8, 175) <= 1; playAgain_W(8, 176) <= 0; playAgain_W(8, 177) <= 0; playAgain_W(8, 178) <= 0; playAgain_W(8, 179) <= 0; playAgain_W(8, 180) <= 0; playAgain_W(8, 181) <= 0; playAgain_W(8, 182) <= 0; playAgain_W(8, 183) <= 0; playAgain_W(8, 184) <= 0; playAgain_W(8, 185) <= 0; playAgain_W(8, 186) <= 0; playAgain_W(8, 187) <= 0; playAgain_W(8, 188) <= 0; playAgain_W(8, 189) <= 0; playAgain_W(8, 190) <= 0; playAgain_W(8, 191) <= 0; playAgain_W(8, 192) <= 0; playAgain_W(8, 193) <= 0; playAgain_W(8, 194) <= 0; playAgain_W(8, 195) <= 0; playAgain_W(8, 196) <= 0; playAgain_W(8, 197) <= 0; playAgain_W(8, 198) <= 0; playAgain_W(8, 199) <= 0; playAgain_W(8, 200) <= 0; playAgain_W(8, 201) <= 0; playAgain_W(8, 202) <= 0; playAgain_W(8, 203) <= 0; playAgain_W(8, 204) <= 0; playAgain_W(8, 205) <= 0; playAgain_W(8, 206) <= 0; playAgain_W(8, 207) <= 0; playAgain_W(8, 208) <= 0; playAgain_W(8, 209) <= 0; playAgain_W(8, 210) <= 0; playAgain_W(8, 211) <= 0; playAgain_W(8, 212) <= 0; playAgain_W(8, 213) <= 0; playAgain_W(8, 214) <= 0; playAgain_W(8, 215) <= 0; playAgain_W(8, 216) <= 0; playAgain_W(8, 217) <= 0; playAgain_W(8, 218) <= 1; playAgain_W(8, 219) <= 1; playAgain_W(8, 220) <= 1; playAgain_W(8, 221) <= 1; playAgain_W(8, 222) <= 1; playAgain_W(8, 223) <= 1; playAgain_W(8, 224) <= 1; playAgain_W(8, 225) <= 1; playAgain_W(8, 226) <= 1; playAgain_W(8, 227) <= 1; playAgain_W(8, 228) <= 0; playAgain_W(8, 229) <= 0; playAgain_W(8, 230) <= 0; playAgain_W(8, 231) <= 0; playAgain_W(8, 232) <= 0; playAgain_W(8, 233) <= 0; playAgain_W(8, 234) <= 0; playAgain_W(8, 235) <= 0; playAgain_W(8, 236) <= 0; playAgain_W(8, 237) <= 0; playAgain_W(8, 238) <= 0; playAgain_W(8, 239) <= 0; playAgain_W(8, 240) <= 1; playAgain_W(8, 241) <= 1; playAgain_W(8, 242) <= 1; playAgain_W(8, 243) <= 1; playAgain_W(8, 244) <= 0; playAgain_W(8, 245) <= 0; playAgain_W(8, 246) <= 0; playAgain_W(8, 247) <= 0; playAgain_W(8, 248) <= 0; playAgain_W(8, 249) <= 0; playAgain_W(8, 250) <= 0; playAgain_W(8, 251) <= 0; playAgain_W(8, 252) <= 1; playAgain_W(8, 253) <= 1; playAgain_W(8, 254) <= 1; playAgain_W(8, 255) <= 1; playAgain_W(8, 256) <= 0; playAgain_W(8, 257) <= 0; playAgain_W(8, 258) <= 1; playAgain_W(8, 259) <= 1; playAgain_W(8, 260) <= 1; playAgain_W(8, 261) <= 1; playAgain_W(8, 262) <= 1; playAgain_W(8, 263) <= 1; playAgain_W(8, 264) <= 1; playAgain_W(8, 265) <= 1; playAgain_W(8, 266) <= 0; playAgain_W(8, 267) <= 0; playAgain_W(8, 268) <= 0; playAgain_W(8, 269) <= 0; playAgain_W(8, 270) <= 0; playAgain_W(8, 271) <= 0; playAgain_W(8, 272) <= 1; playAgain_W(8, 273) <= 1; playAgain_W(8, 274) <= 1; playAgain_W(8, 275) <= 1; playAgain_W(8, 276) <= 0; playAgain_W(8, 277) <= 0; playAgain_W(8, 278) <= 0; playAgain_W(8, 279) <= 0; playAgain_W(8, 280) <= 1; playAgain_W(8, 281) <= 1; playAgain_W(8, 282) <= 1; playAgain_W(8, 283) <= 1; playAgain_W(8, 284) <= 0; playAgain_W(8, 285) <= 0; playAgain_W(8, 286) <= 0; playAgain_W(8, 287) <= 0; 
playAgain_W(9, 0) <= 0; playAgain_W(9, 1) <= 0; playAgain_W(9, 2) <= 1; playAgain_W(9, 3) <= 1; playAgain_W(9, 4) <= 1; playAgain_W(9, 5) <= 1; playAgain_W(9, 6) <= 1; playAgain_W(9, 7) <= 1; playAgain_W(9, 8) <= 1; playAgain_W(9, 9) <= 1; playAgain_W(9, 10) <= 1; playAgain_W(9, 11) <= 1; playAgain_W(9, 12) <= 0; playAgain_W(9, 13) <= 0; playAgain_W(9, 14) <= 0; playAgain_W(9, 15) <= 0; playAgain_W(9, 16) <= 0; playAgain_W(9, 17) <= 0; playAgain_W(9, 18) <= 0; playAgain_W(9, 19) <= 0; playAgain_W(9, 20) <= 1; playAgain_W(9, 21) <= 1; playAgain_W(9, 22) <= 1; playAgain_W(9, 23) <= 1; playAgain_W(9, 24) <= 0; playAgain_W(9, 25) <= 0; playAgain_W(9, 26) <= 0; playAgain_W(9, 27) <= 0; playAgain_W(9, 28) <= 0; playAgain_W(9, 29) <= 0; playAgain_W(9, 30) <= 0; playAgain_W(9, 31) <= 0; playAgain_W(9, 32) <= 0; playAgain_W(9, 33) <= 0; playAgain_W(9, 34) <= 0; playAgain_W(9, 35) <= 0; playAgain_W(9, 36) <= 1; playAgain_W(9, 37) <= 1; playAgain_W(9, 38) <= 1; playAgain_W(9, 39) <= 1; playAgain_W(9, 40) <= 0; playAgain_W(9, 41) <= 0; playAgain_W(9, 42) <= 0; playAgain_W(9, 43) <= 0; playAgain_W(9, 44) <= 0; playAgain_W(9, 45) <= 0; playAgain_W(9, 46) <= 1; playAgain_W(9, 47) <= 1; playAgain_W(9, 48) <= 1; playAgain_W(9, 49) <= 1; playAgain_W(9, 50) <= 0; playAgain_W(9, 51) <= 0; playAgain_W(9, 52) <= 0; playAgain_W(9, 53) <= 0; playAgain_W(9, 54) <= 0; playAgain_W(9, 55) <= 0; playAgain_W(9, 56) <= 0; playAgain_W(9, 57) <= 0; playAgain_W(9, 58) <= 1; playAgain_W(9, 59) <= 1; playAgain_W(9, 60) <= 1; playAgain_W(9, 61) <= 1; playAgain_W(9, 62) <= 1; playAgain_W(9, 63) <= 1; playAgain_W(9, 64) <= 1; playAgain_W(9, 65) <= 1; playAgain_W(9, 66) <= 0; playAgain_W(9, 67) <= 0; playAgain_W(9, 68) <= 0; playAgain_W(9, 69) <= 0; playAgain_W(9, 70) <= 0; playAgain_W(9, 71) <= 0; playAgain_W(9, 72) <= 0; playAgain_W(9, 73) <= 0; playAgain_W(9, 74) <= 0; playAgain_W(9, 75) <= 0; playAgain_W(9, 76) <= 0; playAgain_W(9, 77) <= 0; playAgain_W(9, 78) <= 0; playAgain_W(9, 79) <= 0; playAgain_W(9, 80) <= 0; playAgain_W(9, 81) <= 0; playAgain_W(9, 82) <= 0; playAgain_W(9, 83) <= 0; playAgain_W(9, 84) <= 0; playAgain_W(9, 85) <= 0; playAgain_W(9, 86) <= 0; playAgain_W(9, 87) <= 0; playAgain_W(9, 88) <= 0; playAgain_W(9, 89) <= 0; playAgain_W(9, 90) <= 1; playAgain_W(9, 91) <= 1; playAgain_W(9, 92) <= 1; playAgain_W(9, 93) <= 1; playAgain_W(9, 94) <= 0; playAgain_W(9, 95) <= 0; playAgain_W(9, 96) <= 0; playAgain_W(9, 97) <= 0; playAgain_W(9, 98) <= 0; playAgain_W(9, 99) <= 0; playAgain_W(9, 100) <= 1; playAgain_W(9, 101) <= 1; playAgain_W(9, 102) <= 1; playAgain_W(9, 103) <= 1; playAgain_W(9, 104) <= 0; playAgain_W(9, 105) <= 0; playAgain_W(9, 106) <= 0; playAgain_W(9, 107) <= 0; playAgain_W(9, 108) <= 1; playAgain_W(9, 109) <= 1; playAgain_W(9, 110) <= 1; playAgain_W(9, 111) <= 1; playAgain_W(9, 112) <= 0; playAgain_W(9, 113) <= 0; playAgain_W(9, 114) <= 0; playAgain_W(9, 115) <= 0; playAgain_W(9, 116) <= 0; playAgain_W(9, 117) <= 0; playAgain_W(9, 118) <= 0; playAgain_W(9, 119) <= 0; playAgain_W(9, 120) <= 0; playAgain_W(9, 121) <= 0; playAgain_W(9, 122) <= 0; playAgain_W(9, 123) <= 0; playAgain_W(9, 124) <= 0; playAgain_W(9, 125) <= 0; playAgain_W(9, 126) <= 1; playAgain_W(9, 127) <= 1; playAgain_W(9, 128) <= 1; playAgain_W(9, 129) <= 1; playAgain_W(9, 130) <= 0; playAgain_W(9, 131) <= 0; playAgain_W(9, 132) <= 0; playAgain_W(9, 133) <= 0; playAgain_W(9, 134) <= 0; playAgain_W(9, 135) <= 0; playAgain_W(9, 136) <= 1; playAgain_W(9, 137) <= 1; playAgain_W(9, 138) <= 1; playAgain_W(9, 139) <= 1; playAgain_W(9, 140) <= 0; playAgain_W(9, 141) <= 0; playAgain_W(9, 142) <= 0; playAgain_W(9, 143) <= 0; playAgain_W(9, 144) <= 0; playAgain_W(9, 145) <= 0; playAgain_W(9, 146) <= 0; playAgain_W(9, 147) <= 0; playAgain_W(9, 148) <= 0; playAgain_W(9, 149) <= 0; playAgain_W(9, 150) <= 1; playAgain_W(9, 151) <= 1; playAgain_W(9, 152) <= 1; playAgain_W(9, 153) <= 1; playAgain_W(9, 154) <= 0; playAgain_W(9, 155) <= 0; playAgain_W(9, 156) <= 0; playAgain_W(9, 157) <= 0; playAgain_W(9, 158) <= 0; playAgain_W(9, 159) <= 0; playAgain_W(9, 160) <= 0; playAgain_W(9, 161) <= 0; playAgain_W(9, 162) <= 1; playAgain_W(9, 163) <= 1; playAgain_W(9, 164) <= 1; playAgain_W(9, 165) <= 1; playAgain_W(9, 166) <= 0; playAgain_W(9, 167) <= 0; playAgain_W(9, 168) <= 1; playAgain_W(9, 169) <= 1; playAgain_W(9, 170) <= 1; playAgain_W(9, 171) <= 1; playAgain_W(9, 172) <= 1; playAgain_W(9, 173) <= 1; playAgain_W(9, 174) <= 1; playAgain_W(9, 175) <= 1; playAgain_W(9, 176) <= 0; playAgain_W(9, 177) <= 0; playAgain_W(9, 178) <= 0; playAgain_W(9, 179) <= 0; playAgain_W(9, 180) <= 0; playAgain_W(9, 181) <= 0; playAgain_W(9, 182) <= 0; playAgain_W(9, 183) <= 0; playAgain_W(9, 184) <= 0; playAgain_W(9, 185) <= 0; playAgain_W(9, 186) <= 0; playAgain_W(9, 187) <= 0; playAgain_W(9, 188) <= 0; playAgain_W(9, 189) <= 0; playAgain_W(9, 190) <= 0; playAgain_W(9, 191) <= 0; playAgain_W(9, 192) <= 0; playAgain_W(9, 193) <= 0; playAgain_W(9, 194) <= 0; playAgain_W(9, 195) <= 0; playAgain_W(9, 196) <= 0; playAgain_W(9, 197) <= 0; playAgain_W(9, 198) <= 0; playAgain_W(9, 199) <= 0; playAgain_W(9, 200) <= 0; playAgain_W(9, 201) <= 0; playAgain_W(9, 202) <= 0; playAgain_W(9, 203) <= 0; playAgain_W(9, 204) <= 0; playAgain_W(9, 205) <= 0; playAgain_W(9, 206) <= 0; playAgain_W(9, 207) <= 0; playAgain_W(9, 208) <= 0; playAgain_W(9, 209) <= 0; playAgain_W(9, 210) <= 0; playAgain_W(9, 211) <= 0; playAgain_W(9, 212) <= 0; playAgain_W(9, 213) <= 0; playAgain_W(9, 214) <= 0; playAgain_W(9, 215) <= 0; playAgain_W(9, 216) <= 0; playAgain_W(9, 217) <= 0; playAgain_W(9, 218) <= 1; playAgain_W(9, 219) <= 1; playAgain_W(9, 220) <= 1; playAgain_W(9, 221) <= 1; playAgain_W(9, 222) <= 1; playAgain_W(9, 223) <= 1; playAgain_W(9, 224) <= 1; playAgain_W(9, 225) <= 1; playAgain_W(9, 226) <= 1; playAgain_W(9, 227) <= 1; playAgain_W(9, 228) <= 0; playAgain_W(9, 229) <= 0; playAgain_W(9, 230) <= 0; playAgain_W(9, 231) <= 0; playAgain_W(9, 232) <= 0; playAgain_W(9, 233) <= 0; playAgain_W(9, 234) <= 0; playAgain_W(9, 235) <= 0; playAgain_W(9, 236) <= 0; playAgain_W(9, 237) <= 0; playAgain_W(9, 238) <= 0; playAgain_W(9, 239) <= 0; playAgain_W(9, 240) <= 1; playAgain_W(9, 241) <= 1; playAgain_W(9, 242) <= 1; playAgain_W(9, 243) <= 1; playAgain_W(9, 244) <= 0; playAgain_W(9, 245) <= 0; playAgain_W(9, 246) <= 0; playAgain_W(9, 247) <= 0; playAgain_W(9, 248) <= 0; playAgain_W(9, 249) <= 0; playAgain_W(9, 250) <= 0; playAgain_W(9, 251) <= 0; playAgain_W(9, 252) <= 1; playAgain_W(9, 253) <= 1; playAgain_W(9, 254) <= 1; playAgain_W(9, 255) <= 1; playAgain_W(9, 256) <= 0; playAgain_W(9, 257) <= 0; playAgain_W(9, 258) <= 1; playAgain_W(9, 259) <= 1; playAgain_W(9, 260) <= 1; playAgain_W(9, 261) <= 1; playAgain_W(9, 262) <= 1; playAgain_W(9, 263) <= 1; playAgain_W(9, 264) <= 1; playAgain_W(9, 265) <= 1; playAgain_W(9, 266) <= 0; playAgain_W(9, 267) <= 0; playAgain_W(9, 268) <= 0; playAgain_W(9, 269) <= 0; playAgain_W(9, 270) <= 0; playAgain_W(9, 271) <= 0; playAgain_W(9, 272) <= 1; playAgain_W(9, 273) <= 1; playAgain_W(9, 274) <= 1; playAgain_W(9, 275) <= 1; playAgain_W(9, 276) <= 0; playAgain_W(9, 277) <= 0; playAgain_W(9, 278) <= 0; playAgain_W(9, 279) <= 0; playAgain_W(9, 280) <= 1; playAgain_W(9, 281) <= 1; playAgain_W(9, 282) <= 1; playAgain_W(9, 283) <= 1; playAgain_W(9, 284) <= 0; playAgain_W(9, 285) <= 0; playAgain_W(9, 286) <= 0; playAgain_W(9, 287) <= 0; 
playAgain_W(10, 0) <= 0; playAgain_W(10, 1) <= 0; playAgain_W(10, 2) <= 1; playAgain_W(10, 3) <= 1; playAgain_W(10, 4) <= 1; playAgain_W(10, 5) <= 1; playAgain_W(10, 6) <= 0; playAgain_W(10, 7) <= 0; playAgain_W(10, 8) <= 0; playAgain_W(10, 9) <= 0; playAgain_W(10, 10) <= 0; playAgain_W(10, 11) <= 0; playAgain_W(10, 12) <= 0; playAgain_W(10, 13) <= 0; playAgain_W(10, 14) <= 0; playAgain_W(10, 15) <= 0; playAgain_W(10, 16) <= 0; playAgain_W(10, 17) <= 0; playAgain_W(10, 18) <= 0; playAgain_W(10, 19) <= 0; playAgain_W(10, 20) <= 1; playAgain_W(10, 21) <= 1; playAgain_W(10, 22) <= 1; playAgain_W(10, 23) <= 1; playAgain_W(10, 24) <= 0; playAgain_W(10, 25) <= 0; playAgain_W(10, 26) <= 0; playAgain_W(10, 27) <= 0; playAgain_W(10, 28) <= 0; playAgain_W(10, 29) <= 0; playAgain_W(10, 30) <= 0; playAgain_W(10, 31) <= 0; playAgain_W(10, 32) <= 0; playAgain_W(10, 33) <= 0; playAgain_W(10, 34) <= 0; playAgain_W(10, 35) <= 0; playAgain_W(10, 36) <= 1; playAgain_W(10, 37) <= 1; playAgain_W(10, 38) <= 1; playAgain_W(10, 39) <= 1; playAgain_W(10, 40) <= 1; playAgain_W(10, 41) <= 1; playAgain_W(10, 42) <= 1; playAgain_W(10, 43) <= 1; playAgain_W(10, 44) <= 1; playAgain_W(10, 45) <= 1; playAgain_W(10, 46) <= 1; playAgain_W(10, 47) <= 1; playAgain_W(10, 48) <= 1; playAgain_W(10, 49) <= 1; playAgain_W(10, 50) <= 0; playAgain_W(10, 51) <= 0; playAgain_W(10, 52) <= 0; playAgain_W(10, 53) <= 0; playAgain_W(10, 54) <= 0; playAgain_W(10, 55) <= 0; playAgain_W(10, 56) <= 0; playAgain_W(10, 57) <= 0; playAgain_W(10, 58) <= 0; playAgain_W(10, 59) <= 0; playAgain_W(10, 60) <= 1; playAgain_W(10, 61) <= 1; playAgain_W(10, 62) <= 1; playAgain_W(10, 63) <= 1; playAgain_W(10, 64) <= 0; playAgain_W(10, 65) <= 0; playAgain_W(10, 66) <= 0; playAgain_W(10, 67) <= 0; playAgain_W(10, 68) <= 0; playAgain_W(10, 69) <= 0; playAgain_W(10, 70) <= 0; playAgain_W(10, 71) <= 0; playAgain_W(10, 72) <= 0; playAgain_W(10, 73) <= 0; playAgain_W(10, 74) <= 0; playAgain_W(10, 75) <= 0; playAgain_W(10, 76) <= 0; playAgain_W(10, 77) <= 0; playAgain_W(10, 78) <= 0; playAgain_W(10, 79) <= 0; playAgain_W(10, 80) <= 0; playAgain_W(10, 81) <= 0; playAgain_W(10, 82) <= 0; playAgain_W(10, 83) <= 0; playAgain_W(10, 84) <= 0; playAgain_W(10, 85) <= 0; playAgain_W(10, 86) <= 0; playAgain_W(10, 87) <= 0; playAgain_W(10, 88) <= 0; playAgain_W(10, 89) <= 0; playAgain_W(10, 90) <= 1; playAgain_W(10, 91) <= 1; playAgain_W(10, 92) <= 1; playAgain_W(10, 93) <= 1; playAgain_W(10, 94) <= 1; playAgain_W(10, 95) <= 1; playAgain_W(10, 96) <= 1; playAgain_W(10, 97) <= 1; playAgain_W(10, 98) <= 1; playAgain_W(10, 99) <= 1; playAgain_W(10, 100) <= 1; playAgain_W(10, 101) <= 1; playAgain_W(10, 102) <= 1; playAgain_W(10, 103) <= 1; playAgain_W(10, 104) <= 0; playAgain_W(10, 105) <= 0; playAgain_W(10, 106) <= 0; playAgain_W(10, 107) <= 0; playAgain_W(10, 108) <= 1; playAgain_W(10, 109) <= 1; playAgain_W(10, 110) <= 1; playAgain_W(10, 111) <= 1; playAgain_W(10, 112) <= 0; playAgain_W(10, 113) <= 0; playAgain_W(10, 114) <= 1; playAgain_W(10, 115) <= 1; playAgain_W(10, 116) <= 1; playAgain_W(10, 117) <= 1; playAgain_W(10, 118) <= 1; playAgain_W(10, 119) <= 1; playAgain_W(10, 120) <= 1; playAgain_W(10, 121) <= 1; playAgain_W(10, 122) <= 0; playAgain_W(10, 123) <= 0; playAgain_W(10, 124) <= 0; playAgain_W(10, 125) <= 0; playAgain_W(10, 126) <= 1; playAgain_W(10, 127) <= 1; playAgain_W(10, 128) <= 1; playAgain_W(10, 129) <= 1; playAgain_W(10, 130) <= 1; playAgain_W(10, 131) <= 1; playAgain_W(10, 132) <= 1; playAgain_W(10, 133) <= 1; playAgain_W(10, 134) <= 1; playAgain_W(10, 135) <= 1; playAgain_W(10, 136) <= 1; playAgain_W(10, 137) <= 1; playAgain_W(10, 138) <= 1; playAgain_W(10, 139) <= 1; playAgain_W(10, 140) <= 0; playAgain_W(10, 141) <= 0; playAgain_W(10, 142) <= 0; playAgain_W(10, 143) <= 0; playAgain_W(10, 144) <= 0; playAgain_W(10, 145) <= 0; playAgain_W(10, 146) <= 0; playAgain_W(10, 147) <= 0; playAgain_W(10, 148) <= 0; playAgain_W(10, 149) <= 0; playAgain_W(10, 150) <= 1; playAgain_W(10, 151) <= 1; playAgain_W(10, 152) <= 1; playAgain_W(10, 153) <= 1; playAgain_W(10, 154) <= 0; playAgain_W(10, 155) <= 0; playAgain_W(10, 156) <= 0; playAgain_W(10, 157) <= 0; playAgain_W(10, 158) <= 0; playAgain_W(10, 159) <= 0; playAgain_W(10, 160) <= 0; playAgain_W(10, 161) <= 0; playAgain_W(10, 162) <= 1; playAgain_W(10, 163) <= 1; playAgain_W(10, 164) <= 1; playAgain_W(10, 165) <= 1; playAgain_W(10, 166) <= 0; playAgain_W(10, 167) <= 0; playAgain_W(10, 168) <= 0; playAgain_W(10, 169) <= 0; playAgain_W(10, 170) <= 1; playAgain_W(10, 171) <= 1; playAgain_W(10, 172) <= 1; playAgain_W(10, 173) <= 1; playAgain_W(10, 174) <= 1; playAgain_W(10, 175) <= 1; playAgain_W(10, 176) <= 0; playAgain_W(10, 177) <= 0; playAgain_W(10, 178) <= 0; playAgain_W(10, 179) <= 0; playAgain_W(10, 180) <= 0; playAgain_W(10, 181) <= 0; playAgain_W(10, 182) <= 0; playAgain_W(10, 183) <= 0; playAgain_W(10, 184) <= 0; playAgain_W(10, 185) <= 0; playAgain_W(10, 186) <= 0; playAgain_W(10, 187) <= 0; playAgain_W(10, 188) <= 0; playAgain_W(10, 189) <= 0; playAgain_W(10, 190) <= 0; playAgain_W(10, 191) <= 0; playAgain_W(10, 192) <= 0; playAgain_W(10, 193) <= 0; playAgain_W(10, 194) <= 0; playAgain_W(10, 195) <= 0; playAgain_W(10, 196) <= 0; playAgain_W(10, 197) <= 0; playAgain_W(10, 198) <= 0; playAgain_W(10, 199) <= 0; playAgain_W(10, 200) <= 0; playAgain_W(10, 201) <= 0; playAgain_W(10, 202) <= 0; playAgain_W(10, 203) <= 0; playAgain_W(10, 204) <= 0; playAgain_W(10, 205) <= 0; playAgain_W(10, 206) <= 0; playAgain_W(10, 207) <= 0; playAgain_W(10, 208) <= 0; playAgain_W(10, 209) <= 0; playAgain_W(10, 210) <= 0; playAgain_W(10, 211) <= 0; playAgain_W(10, 212) <= 0; playAgain_W(10, 213) <= 0; playAgain_W(10, 214) <= 0; playAgain_W(10, 215) <= 0; playAgain_W(10, 216) <= 0; playAgain_W(10, 217) <= 0; playAgain_W(10, 218) <= 1; playAgain_W(10, 219) <= 1; playAgain_W(10, 220) <= 1; playAgain_W(10, 221) <= 1; playAgain_W(10, 222) <= 0; playAgain_W(10, 223) <= 0; playAgain_W(10, 224) <= 0; playAgain_W(10, 225) <= 0; playAgain_W(10, 226) <= 1; playAgain_W(10, 227) <= 1; playAgain_W(10, 228) <= 1; playAgain_W(10, 229) <= 1; playAgain_W(10, 230) <= 0; playAgain_W(10, 231) <= 0; playAgain_W(10, 232) <= 0; playAgain_W(10, 233) <= 0; playAgain_W(10, 234) <= 0; playAgain_W(10, 235) <= 0; playAgain_W(10, 236) <= 0; playAgain_W(10, 237) <= 0; playAgain_W(10, 238) <= 0; playAgain_W(10, 239) <= 0; playAgain_W(10, 240) <= 1; playAgain_W(10, 241) <= 1; playAgain_W(10, 242) <= 1; playAgain_W(10, 243) <= 1; playAgain_W(10, 244) <= 0; playAgain_W(10, 245) <= 0; playAgain_W(10, 246) <= 0; playAgain_W(10, 247) <= 0; playAgain_W(10, 248) <= 0; playAgain_W(10, 249) <= 0; playAgain_W(10, 250) <= 0; playAgain_W(10, 251) <= 0; playAgain_W(10, 252) <= 1; playAgain_W(10, 253) <= 1; playAgain_W(10, 254) <= 1; playAgain_W(10, 255) <= 1; playAgain_W(10, 256) <= 0; playAgain_W(10, 257) <= 0; playAgain_W(10, 258) <= 0; playAgain_W(10, 259) <= 0; playAgain_W(10, 260) <= 1; playAgain_W(10, 261) <= 1; playAgain_W(10, 262) <= 1; playAgain_W(10, 263) <= 1; playAgain_W(10, 264) <= 1; playAgain_W(10, 265) <= 1; playAgain_W(10, 266) <= 0; playAgain_W(10, 267) <= 0; playAgain_W(10, 268) <= 0; playAgain_W(10, 269) <= 0; playAgain_W(10, 270) <= 0; playAgain_W(10, 271) <= 0; playAgain_W(10, 272) <= 1; playAgain_W(10, 273) <= 1; playAgain_W(10, 274) <= 1; playAgain_W(10, 275) <= 1; playAgain_W(10, 276) <= 0; playAgain_W(10, 277) <= 0; playAgain_W(10, 278) <= 0; playAgain_W(10, 279) <= 0; playAgain_W(10, 280) <= 1; playAgain_W(10, 281) <= 1; playAgain_W(10, 282) <= 1; playAgain_W(10, 283) <= 1; playAgain_W(10, 284) <= 0; playAgain_W(10, 285) <= 0; playAgain_W(10, 286) <= 0; playAgain_W(10, 287) <= 0; 
playAgain_W(11, 0) <= 0; playAgain_W(11, 1) <= 0; playAgain_W(11, 2) <= 1; playAgain_W(11, 3) <= 1; playAgain_W(11, 4) <= 1; playAgain_W(11, 5) <= 1; playAgain_W(11, 6) <= 0; playAgain_W(11, 7) <= 0; playAgain_W(11, 8) <= 0; playAgain_W(11, 9) <= 0; playAgain_W(11, 10) <= 0; playAgain_W(11, 11) <= 0; playAgain_W(11, 12) <= 0; playAgain_W(11, 13) <= 0; playAgain_W(11, 14) <= 0; playAgain_W(11, 15) <= 0; playAgain_W(11, 16) <= 0; playAgain_W(11, 17) <= 0; playAgain_W(11, 18) <= 0; playAgain_W(11, 19) <= 0; playAgain_W(11, 20) <= 1; playAgain_W(11, 21) <= 1; playAgain_W(11, 22) <= 1; playAgain_W(11, 23) <= 1; playAgain_W(11, 24) <= 0; playAgain_W(11, 25) <= 0; playAgain_W(11, 26) <= 0; playAgain_W(11, 27) <= 0; playAgain_W(11, 28) <= 0; playAgain_W(11, 29) <= 0; playAgain_W(11, 30) <= 0; playAgain_W(11, 31) <= 0; playAgain_W(11, 32) <= 0; playAgain_W(11, 33) <= 0; playAgain_W(11, 34) <= 0; playAgain_W(11, 35) <= 0; playAgain_W(11, 36) <= 1; playAgain_W(11, 37) <= 1; playAgain_W(11, 38) <= 1; playAgain_W(11, 39) <= 1; playAgain_W(11, 40) <= 1; playAgain_W(11, 41) <= 1; playAgain_W(11, 42) <= 1; playAgain_W(11, 43) <= 1; playAgain_W(11, 44) <= 1; playAgain_W(11, 45) <= 1; playAgain_W(11, 46) <= 1; playAgain_W(11, 47) <= 1; playAgain_W(11, 48) <= 1; playAgain_W(11, 49) <= 1; playAgain_W(11, 50) <= 0; playAgain_W(11, 51) <= 0; playAgain_W(11, 52) <= 0; playAgain_W(11, 53) <= 0; playAgain_W(11, 54) <= 0; playAgain_W(11, 55) <= 0; playAgain_W(11, 56) <= 0; playAgain_W(11, 57) <= 0; playAgain_W(11, 58) <= 0; playAgain_W(11, 59) <= 0; playAgain_W(11, 60) <= 1; playAgain_W(11, 61) <= 1; playAgain_W(11, 62) <= 1; playAgain_W(11, 63) <= 1; playAgain_W(11, 64) <= 0; playAgain_W(11, 65) <= 0; playAgain_W(11, 66) <= 0; playAgain_W(11, 67) <= 0; playAgain_W(11, 68) <= 0; playAgain_W(11, 69) <= 0; playAgain_W(11, 70) <= 0; playAgain_W(11, 71) <= 0; playAgain_W(11, 72) <= 0; playAgain_W(11, 73) <= 0; playAgain_W(11, 74) <= 0; playAgain_W(11, 75) <= 0; playAgain_W(11, 76) <= 0; playAgain_W(11, 77) <= 0; playAgain_W(11, 78) <= 0; playAgain_W(11, 79) <= 0; playAgain_W(11, 80) <= 0; playAgain_W(11, 81) <= 0; playAgain_W(11, 82) <= 0; playAgain_W(11, 83) <= 0; playAgain_W(11, 84) <= 0; playAgain_W(11, 85) <= 0; playAgain_W(11, 86) <= 0; playAgain_W(11, 87) <= 0; playAgain_W(11, 88) <= 0; playAgain_W(11, 89) <= 0; playAgain_W(11, 90) <= 1; playAgain_W(11, 91) <= 1; playAgain_W(11, 92) <= 1; playAgain_W(11, 93) <= 1; playAgain_W(11, 94) <= 1; playAgain_W(11, 95) <= 1; playAgain_W(11, 96) <= 1; playAgain_W(11, 97) <= 1; playAgain_W(11, 98) <= 1; playAgain_W(11, 99) <= 1; playAgain_W(11, 100) <= 1; playAgain_W(11, 101) <= 1; playAgain_W(11, 102) <= 1; playAgain_W(11, 103) <= 1; playAgain_W(11, 104) <= 0; playAgain_W(11, 105) <= 0; playAgain_W(11, 106) <= 0; playAgain_W(11, 107) <= 0; playAgain_W(11, 108) <= 1; playAgain_W(11, 109) <= 1; playAgain_W(11, 110) <= 1; playAgain_W(11, 111) <= 1; playAgain_W(11, 112) <= 0; playAgain_W(11, 113) <= 0; playAgain_W(11, 114) <= 1; playAgain_W(11, 115) <= 1; playAgain_W(11, 116) <= 1; playAgain_W(11, 117) <= 1; playAgain_W(11, 118) <= 1; playAgain_W(11, 119) <= 1; playAgain_W(11, 120) <= 1; playAgain_W(11, 121) <= 1; playAgain_W(11, 122) <= 0; playAgain_W(11, 123) <= 0; playAgain_W(11, 124) <= 0; playAgain_W(11, 125) <= 0; playAgain_W(11, 126) <= 1; playAgain_W(11, 127) <= 1; playAgain_W(11, 128) <= 1; playAgain_W(11, 129) <= 1; playAgain_W(11, 130) <= 1; playAgain_W(11, 131) <= 1; playAgain_W(11, 132) <= 1; playAgain_W(11, 133) <= 1; playAgain_W(11, 134) <= 1; playAgain_W(11, 135) <= 1; playAgain_W(11, 136) <= 1; playAgain_W(11, 137) <= 1; playAgain_W(11, 138) <= 1; playAgain_W(11, 139) <= 1; playAgain_W(11, 140) <= 0; playAgain_W(11, 141) <= 0; playAgain_W(11, 142) <= 0; playAgain_W(11, 143) <= 0; playAgain_W(11, 144) <= 0; playAgain_W(11, 145) <= 0; playAgain_W(11, 146) <= 0; playAgain_W(11, 147) <= 0; playAgain_W(11, 148) <= 0; playAgain_W(11, 149) <= 0; playAgain_W(11, 150) <= 1; playAgain_W(11, 151) <= 1; playAgain_W(11, 152) <= 1; playAgain_W(11, 153) <= 1; playAgain_W(11, 154) <= 0; playAgain_W(11, 155) <= 0; playAgain_W(11, 156) <= 0; playAgain_W(11, 157) <= 0; playAgain_W(11, 158) <= 0; playAgain_W(11, 159) <= 0; playAgain_W(11, 160) <= 0; playAgain_W(11, 161) <= 0; playAgain_W(11, 162) <= 1; playAgain_W(11, 163) <= 1; playAgain_W(11, 164) <= 1; playAgain_W(11, 165) <= 1; playAgain_W(11, 166) <= 0; playAgain_W(11, 167) <= 0; playAgain_W(11, 168) <= 0; playAgain_W(11, 169) <= 0; playAgain_W(11, 170) <= 1; playAgain_W(11, 171) <= 1; playAgain_W(11, 172) <= 1; playAgain_W(11, 173) <= 1; playAgain_W(11, 174) <= 1; playAgain_W(11, 175) <= 1; playAgain_W(11, 176) <= 0; playAgain_W(11, 177) <= 0; playAgain_W(11, 178) <= 0; playAgain_W(11, 179) <= 0; playAgain_W(11, 180) <= 0; playAgain_W(11, 181) <= 0; playAgain_W(11, 182) <= 0; playAgain_W(11, 183) <= 0; playAgain_W(11, 184) <= 0; playAgain_W(11, 185) <= 0; playAgain_W(11, 186) <= 0; playAgain_W(11, 187) <= 0; playAgain_W(11, 188) <= 0; playAgain_W(11, 189) <= 0; playAgain_W(11, 190) <= 0; playAgain_W(11, 191) <= 0; playAgain_W(11, 192) <= 0; playAgain_W(11, 193) <= 0; playAgain_W(11, 194) <= 0; playAgain_W(11, 195) <= 0; playAgain_W(11, 196) <= 0; playAgain_W(11, 197) <= 0; playAgain_W(11, 198) <= 0; playAgain_W(11, 199) <= 0; playAgain_W(11, 200) <= 0; playAgain_W(11, 201) <= 0; playAgain_W(11, 202) <= 0; playAgain_W(11, 203) <= 0; playAgain_W(11, 204) <= 0; playAgain_W(11, 205) <= 0; playAgain_W(11, 206) <= 0; playAgain_W(11, 207) <= 0; playAgain_W(11, 208) <= 0; playAgain_W(11, 209) <= 0; playAgain_W(11, 210) <= 0; playAgain_W(11, 211) <= 0; playAgain_W(11, 212) <= 0; playAgain_W(11, 213) <= 0; playAgain_W(11, 214) <= 0; playAgain_W(11, 215) <= 0; playAgain_W(11, 216) <= 0; playAgain_W(11, 217) <= 0; playAgain_W(11, 218) <= 1; playAgain_W(11, 219) <= 1; playAgain_W(11, 220) <= 1; playAgain_W(11, 221) <= 1; playAgain_W(11, 222) <= 0; playAgain_W(11, 223) <= 0; playAgain_W(11, 224) <= 0; playAgain_W(11, 225) <= 0; playAgain_W(11, 226) <= 1; playAgain_W(11, 227) <= 1; playAgain_W(11, 228) <= 1; playAgain_W(11, 229) <= 1; playAgain_W(11, 230) <= 0; playAgain_W(11, 231) <= 0; playAgain_W(11, 232) <= 0; playAgain_W(11, 233) <= 0; playAgain_W(11, 234) <= 0; playAgain_W(11, 235) <= 0; playAgain_W(11, 236) <= 0; playAgain_W(11, 237) <= 0; playAgain_W(11, 238) <= 0; playAgain_W(11, 239) <= 0; playAgain_W(11, 240) <= 1; playAgain_W(11, 241) <= 1; playAgain_W(11, 242) <= 1; playAgain_W(11, 243) <= 1; playAgain_W(11, 244) <= 0; playAgain_W(11, 245) <= 0; playAgain_W(11, 246) <= 0; playAgain_W(11, 247) <= 0; playAgain_W(11, 248) <= 0; playAgain_W(11, 249) <= 0; playAgain_W(11, 250) <= 0; playAgain_W(11, 251) <= 0; playAgain_W(11, 252) <= 1; playAgain_W(11, 253) <= 1; playAgain_W(11, 254) <= 1; playAgain_W(11, 255) <= 1; playAgain_W(11, 256) <= 0; playAgain_W(11, 257) <= 0; playAgain_W(11, 258) <= 0; playAgain_W(11, 259) <= 0; playAgain_W(11, 260) <= 1; playAgain_W(11, 261) <= 1; playAgain_W(11, 262) <= 1; playAgain_W(11, 263) <= 1; playAgain_W(11, 264) <= 1; playAgain_W(11, 265) <= 1; playAgain_W(11, 266) <= 0; playAgain_W(11, 267) <= 0; playAgain_W(11, 268) <= 0; playAgain_W(11, 269) <= 0; playAgain_W(11, 270) <= 0; playAgain_W(11, 271) <= 0; playAgain_W(11, 272) <= 1; playAgain_W(11, 273) <= 1; playAgain_W(11, 274) <= 1; playAgain_W(11, 275) <= 1; playAgain_W(11, 276) <= 0; playAgain_W(11, 277) <= 0; playAgain_W(11, 278) <= 0; playAgain_W(11, 279) <= 0; playAgain_W(11, 280) <= 1; playAgain_W(11, 281) <= 1; playAgain_W(11, 282) <= 1; playAgain_W(11, 283) <= 1; playAgain_W(11, 284) <= 0; playAgain_W(11, 285) <= 0; playAgain_W(11, 286) <= 0; playAgain_W(11, 287) <= 0; 
playAgain_W(12, 0) <= 0; playAgain_W(12, 1) <= 0; playAgain_W(12, 2) <= 1; playAgain_W(12, 3) <= 1; playAgain_W(12, 4) <= 1; playAgain_W(12, 5) <= 1; playAgain_W(12, 6) <= 0; playAgain_W(12, 7) <= 0; playAgain_W(12, 8) <= 0; playAgain_W(12, 9) <= 0; playAgain_W(12, 10) <= 0; playAgain_W(12, 11) <= 0; playAgain_W(12, 12) <= 0; playAgain_W(12, 13) <= 0; playAgain_W(12, 14) <= 0; playAgain_W(12, 15) <= 0; playAgain_W(12, 16) <= 0; playAgain_W(12, 17) <= 0; playAgain_W(12, 18) <= 0; playAgain_W(12, 19) <= 0; playAgain_W(12, 20) <= 1; playAgain_W(12, 21) <= 1; playAgain_W(12, 22) <= 1; playAgain_W(12, 23) <= 1; playAgain_W(12, 24) <= 0; playAgain_W(12, 25) <= 0; playAgain_W(12, 26) <= 0; playAgain_W(12, 27) <= 0; playAgain_W(12, 28) <= 0; playAgain_W(12, 29) <= 0; playAgain_W(12, 30) <= 0; playAgain_W(12, 31) <= 0; playAgain_W(12, 32) <= 0; playAgain_W(12, 33) <= 0; playAgain_W(12, 34) <= 0; playAgain_W(12, 35) <= 0; playAgain_W(12, 36) <= 1; playAgain_W(12, 37) <= 1; playAgain_W(12, 38) <= 1; playAgain_W(12, 39) <= 1; playAgain_W(12, 40) <= 0; playAgain_W(12, 41) <= 0; playAgain_W(12, 42) <= 0; playAgain_W(12, 43) <= 0; playAgain_W(12, 44) <= 0; playAgain_W(12, 45) <= 0; playAgain_W(12, 46) <= 1; playAgain_W(12, 47) <= 1; playAgain_W(12, 48) <= 1; playAgain_W(12, 49) <= 1; playAgain_W(12, 50) <= 0; playAgain_W(12, 51) <= 0; playAgain_W(12, 52) <= 0; playAgain_W(12, 53) <= 0; playAgain_W(12, 54) <= 0; playAgain_W(12, 55) <= 0; playAgain_W(12, 56) <= 0; playAgain_W(12, 57) <= 0; playAgain_W(12, 58) <= 0; playAgain_W(12, 59) <= 0; playAgain_W(12, 60) <= 1; playAgain_W(12, 61) <= 1; playAgain_W(12, 62) <= 1; playAgain_W(12, 63) <= 1; playAgain_W(12, 64) <= 0; playAgain_W(12, 65) <= 0; playAgain_W(12, 66) <= 0; playAgain_W(12, 67) <= 0; playAgain_W(12, 68) <= 0; playAgain_W(12, 69) <= 0; playAgain_W(12, 70) <= 0; playAgain_W(12, 71) <= 0; playAgain_W(12, 72) <= 0; playAgain_W(12, 73) <= 0; playAgain_W(12, 74) <= 0; playAgain_W(12, 75) <= 0; playAgain_W(12, 76) <= 0; playAgain_W(12, 77) <= 0; playAgain_W(12, 78) <= 0; playAgain_W(12, 79) <= 0; playAgain_W(12, 80) <= 0; playAgain_W(12, 81) <= 0; playAgain_W(12, 82) <= 0; playAgain_W(12, 83) <= 0; playAgain_W(12, 84) <= 0; playAgain_W(12, 85) <= 0; playAgain_W(12, 86) <= 0; playAgain_W(12, 87) <= 0; playAgain_W(12, 88) <= 0; playAgain_W(12, 89) <= 0; playAgain_W(12, 90) <= 1; playAgain_W(12, 91) <= 1; playAgain_W(12, 92) <= 1; playAgain_W(12, 93) <= 1; playAgain_W(12, 94) <= 0; playAgain_W(12, 95) <= 0; playAgain_W(12, 96) <= 0; playAgain_W(12, 97) <= 0; playAgain_W(12, 98) <= 0; playAgain_W(12, 99) <= 0; playAgain_W(12, 100) <= 1; playAgain_W(12, 101) <= 1; playAgain_W(12, 102) <= 1; playAgain_W(12, 103) <= 1; playAgain_W(12, 104) <= 0; playAgain_W(12, 105) <= 0; playAgain_W(12, 106) <= 0; playAgain_W(12, 107) <= 0; playAgain_W(12, 108) <= 1; playAgain_W(12, 109) <= 1; playAgain_W(12, 110) <= 1; playAgain_W(12, 111) <= 1; playAgain_W(12, 112) <= 0; playAgain_W(12, 113) <= 0; playAgain_W(12, 114) <= 0; playAgain_W(12, 115) <= 0; playAgain_W(12, 116) <= 0; playAgain_W(12, 117) <= 0; playAgain_W(12, 118) <= 1; playAgain_W(12, 119) <= 1; playAgain_W(12, 120) <= 1; playAgain_W(12, 121) <= 1; playAgain_W(12, 122) <= 0; playAgain_W(12, 123) <= 0; playAgain_W(12, 124) <= 0; playAgain_W(12, 125) <= 0; playAgain_W(12, 126) <= 1; playAgain_W(12, 127) <= 1; playAgain_W(12, 128) <= 1; playAgain_W(12, 129) <= 1; playAgain_W(12, 130) <= 0; playAgain_W(12, 131) <= 0; playAgain_W(12, 132) <= 0; playAgain_W(12, 133) <= 0; playAgain_W(12, 134) <= 0; playAgain_W(12, 135) <= 0; playAgain_W(12, 136) <= 1; playAgain_W(12, 137) <= 1; playAgain_W(12, 138) <= 1; playAgain_W(12, 139) <= 1; playAgain_W(12, 140) <= 0; playAgain_W(12, 141) <= 0; playAgain_W(12, 142) <= 0; playAgain_W(12, 143) <= 0; playAgain_W(12, 144) <= 0; playAgain_W(12, 145) <= 0; playAgain_W(12, 146) <= 0; playAgain_W(12, 147) <= 0; playAgain_W(12, 148) <= 0; playAgain_W(12, 149) <= 0; playAgain_W(12, 150) <= 1; playAgain_W(12, 151) <= 1; playAgain_W(12, 152) <= 1; playAgain_W(12, 153) <= 1; playAgain_W(12, 154) <= 0; playAgain_W(12, 155) <= 0; playAgain_W(12, 156) <= 0; playAgain_W(12, 157) <= 0; playAgain_W(12, 158) <= 0; playAgain_W(12, 159) <= 0; playAgain_W(12, 160) <= 0; playAgain_W(12, 161) <= 0; playAgain_W(12, 162) <= 1; playAgain_W(12, 163) <= 1; playAgain_W(12, 164) <= 1; playAgain_W(12, 165) <= 1; playAgain_W(12, 166) <= 0; playAgain_W(12, 167) <= 0; playAgain_W(12, 168) <= 0; playAgain_W(12, 169) <= 0; playAgain_W(12, 170) <= 0; playAgain_W(12, 171) <= 0; playAgain_W(12, 172) <= 1; playAgain_W(12, 173) <= 1; playAgain_W(12, 174) <= 1; playAgain_W(12, 175) <= 1; playAgain_W(12, 176) <= 0; playAgain_W(12, 177) <= 0; playAgain_W(12, 178) <= 0; playAgain_W(12, 179) <= 0; playAgain_W(12, 180) <= 0; playAgain_W(12, 181) <= 0; playAgain_W(12, 182) <= 0; playAgain_W(12, 183) <= 0; playAgain_W(12, 184) <= 0; playAgain_W(12, 185) <= 0; playAgain_W(12, 186) <= 1; playAgain_W(12, 187) <= 1; playAgain_W(12, 188) <= 1; playAgain_W(12, 189) <= 1; playAgain_W(12, 190) <= 0; playAgain_W(12, 191) <= 0; playAgain_W(12, 192) <= 0; playAgain_W(12, 193) <= 0; playAgain_W(12, 194) <= 0; playAgain_W(12, 195) <= 0; playAgain_W(12, 196) <= 0; playAgain_W(12, 197) <= 0; playAgain_W(12, 198) <= 0; playAgain_W(12, 199) <= 0; playAgain_W(12, 200) <= 0; playAgain_W(12, 201) <= 0; playAgain_W(12, 202) <= 0; playAgain_W(12, 203) <= 0; playAgain_W(12, 204) <= 0; playAgain_W(12, 205) <= 0; playAgain_W(12, 206) <= 0; playAgain_W(12, 207) <= 0; playAgain_W(12, 208) <= 0; playAgain_W(12, 209) <= 0; playAgain_W(12, 210) <= 0; playAgain_W(12, 211) <= 0; playAgain_W(12, 212) <= 0; playAgain_W(12, 213) <= 0; playAgain_W(12, 214) <= 0; playAgain_W(12, 215) <= 0; playAgain_W(12, 216) <= 0; playAgain_W(12, 217) <= 0; playAgain_W(12, 218) <= 1; playAgain_W(12, 219) <= 1; playAgain_W(12, 220) <= 1; playAgain_W(12, 221) <= 1; playAgain_W(12, 222) <= 0; playAgain_W(12, 223) <= 0; playAgain_W(12, 224) <= 0; playAgain_W(12, 225) <= 0; playAgain_W(12, 226) <= 1; playAgain_W(12, 227) <= 1; playAgain_W(12, 228) <= 1; playAgain_W(12, 229) <= 1; playAgain_W(12, 230) <= 0; playAgain_W(12, 231) <= 0; playAgain_W(12, 232) <= 0; playAgain_W(12, 233) <= 0; playAgain_W(12, 234) <= 0; playAgain_W(12, 235) <= 0; playAgain_W(12, 236) <= 0; playAgain_W(12, 237) <= 0; playAgain_W(12, 238) <= 0; playAgain_W(12, 239) <= 0; playAgain_W(12, 240) <= 1; playAgain_W(12, 241) <= 1; playAgain_W(12, 242) <= 1; playAgain_W(12, 243) <= 1; playAgain_W(12, 244) <= 0; playAgain_W(12, 245) <= 0; playAgain_W(12, 246) <= 0; playAgain_W(12, 247) <= 0; playAgain_W(12, 248) <= 0; playAgain_W(12, 249) <= 0; playAgain_W(12, 250) <= 0; playAgain_W(12, 251) <= 0; playAgain_W(12, 252) <= 1; playAgain_W(12, 253) <= 1; playAgain_W(12, 254) <= 1; playAgain_W(12, 255) <= 1; playAgain_W(12, 256) <= 0; playAgain_W(12, 257) <= 0; playAgain_W(12, 258) <= 0; playAgain_W(12, 259) <= 0; playAgain_W(12, 260) <= 0; playAgain_W(12, 261) <= 0; playAgain_W(12, 262) <= 1; playAgain_W(12, 263) <= 1; playAgain_W(12, 264) <= 1; playAgain_W(12, 265) <= 1; playAgain_W(12, 266) <= 0; playAgain_W(12, 267) <= 0; playAgain_W(12, 268) <= 0; playAgain_W(12, 269) <= 0; playAgain_W(12, 270) <= 0; playAgain_W(12, 271) <= 0; playAgain_W(12, 272) <= 1; playAgain_W(12, 273) <= 1; playAgain_W(12, 274) <= 1; playAgain_W(12, 275) <= 1; playAgain_W(12, 276) <= 0; playAgain_W(12, 277) <= 0; playAgain_W(12, 278) <= 0; playAgain_W(12, 279) <= 0; playAgain_W(12, 280) <= 1; playAgain_W(12, 281) <= 1; playAgain_W(12, 282) <= 1; playAgain_W(12, 283) <= 1; playAgain_W(12, 284) <= 0; playAgain_W(12, 285) <= 0; playAgain_W(12, 286) <= 0; playAgain_W(12, 287) <= 0; 
playAgain_W(13, 0) <= 0; playAgain_W(13, 1) <= 0; playAgain_W(13, 2) <= 1; playAgain_W(13, 3) <= 1; playAgain_W(13, 4) <= 1; playAgain_W(13, 5) <= 1; playAgain_W(13, 6) <= 0; playAgain_W(13, 7) <= 0; playAgain_W(13, 8) <= 0; playAgain_W(13, 9) <= 0; playAgain_W(13, 10) <= 0; playAgain_W(13, 11) <= 0; playAgain_W(13, 12) <= 0; playAgain_W(13, 13) <= 0; playAgain_W(13, 14) <= 0; playAgain_W(13, 15) <= 0; playAgain_W(13, 16) <= 0; playAgain_W(13, 17) <= 0; playAgain_W(13, 18) <= 0; playAgain_W(13, 19) <= 0; playAgain_W(13, 20) <= 1; playAgain_W(13, 21) <= 1; playAgain_W(13, 22) <= 1; playAgain_W(13, 23) <= 1; playAgain_W(13, 24) <= 0; playAgain_W(13, 25) <= 0; playAgain_W(13, 26) <= 0; playAgain_W(13, 27) <= 0; playAgain_W(13, 28) <= 0; playAgain_W(13, 29) <= 0; playAgain_W(13, 30) <= 0; playAgain_W(13, 31) <= 0; playAgain_W(13, 32) <= 0; playAgain_W(13, 33) <= 0; playAgain_W(13, 34) <= 0; playAgain_W(13, 35) <= 0; playAgain_W(13, 36) <= 1; playAgain_W(13, 37) <= 1; playAgain_W(13, 38) <= 1; playAgain_W(13, 39) <= 1; playAgain_W(13, 40) <= 0; playAgain_W(13, 41) <= 0; playAgain_W(13, 42) <= 0; playAgain_W(13, 43) <= 0; playAgain_W(13, 44) <= 0; playAgain_W(13, 45) <= 0; playAgain_W(13, 46) <= 1; playAgain_W(13, 47) <= 1; playAgain_W(13, 48) <= 1; playAgain_W(13, 49) <= 1; playAgain_W(13, 50) <= 0; playAgain_W(13, 51) <= 0; playAgain_W(13, 52) <= 0; playAgain_W(13, 53) <= 0; playAgain_W(13, 54) <= 0; playAgain_W(13, 55) <= 0; playAgain_W(13, 56) <= 0; playAgain_W(13, 57) <= 0; playAgain_W(13, 58) <= 0; playAgain_W(13, 59) <= 0; playAgain_W(13, 60) <= 1; playAgain_W(13, 61) <= 1; playAgain_W(13, 62) <= 1; playAgain_W(13, 63) <= 1; playAgain_W(13, 64) <= 0; playAgain_W(13, 65) <= 0; playAgain_W(13, 66) <= 0; playAgain_W(13, 67) <= 0; playAgain_W(13, 68) <= 0; playAgain_W(13, 69) <= 0; playAgain_W(13, 70) <= 0; playAgain_W(13, 71) <= 0; playAgain_W(13, 72) <= 0; playAgain_W(13, 73) <= 0; playAgain_W(13, 74) <= 0; playAgain_W(13, 75) <= 0; playAgain_W(13, 76) <= 0; playAgain_W(13, 77) <= 0; playAgain_W(13, 78) <= 0; playAgain_W(13, 79) <= 0; playAgain_W(13, 80) <= 0; playAgain_W(13, 81) <= 0; playAgain_W(13, 82) <= 0; playAgain_W(13, 83) <= 0; playAgain_W(13, 84) <= 0; playAgain_W(13, 85) <= 0; playAgain_W(13, 86) <= 0; playAgain_W(13, 87) <= 0; playAgain_W(13, 88) <= 0; playAgain_W(13, 89) <= 0; playAgain_W(13, 90) <= 1; playAgain_W(13, 91) <= 1; playAgain_W(13, 92) <= 1; playAgain_W(13, 93) <= 1; playAgain_W(13, 94) <= 0; playAgain_W(13, 95) <= 0; playAgain_W(13, 96) <= 0; playAgain_W(13, 97) <= 0; playAgain_W(13, 98) <= 0; playAgain_W(13, 99) <= 0; playAgain_W(13, 100) <= 1; playAgain_W(13, 101) <= 1; playAgain_W(13, 102) <= 1; playAgain_W(13, 103) <= 1; playAgain_W(13, 104) <= 0; playAgain_W(13, 105) <= 0; playAgain_W(13, 106) <= 0; playAgain_W(13, 107) <= 0; playAgain_W(13, 108) <= 1; playAgain_W(13, 109) <= 1; playAgain_W(13, 110) <= 1; playAgain_W(13, 111) <= 1; playAgain_W(13, 112) <= 0; playAgain_W(13, 113) <= 0; playAgain_W(13, 114) <= 0; playAgain_W(13, 115) <= 0; playAgain_W(13, 116) <= 0; playAgain_W(13, 117) <= 0; playAgain_W(13, 118) <= 1; playAgain_W(13, 119) <= 1; playAgain_W(13, 120) <= 1; playAgain_W(13, 121) <= 1; playAgain_W(13, 122) <= 0; playAgain_W(13, 123) <= 0; playAgain_W(13, 124) <= 0; playAgain_W(13, 125) <= 0; playAgain_W(13, 126) <= 1; playAgain_W(13, 127) <= 1; playAgain_W(13, 128) <= 1; playAgain_W(13, 129) <= 1; playAgain_W(13, 130) <= 0; playAgain_W(13, 131) <= 0; playAgain_W(13, 132) <= 0; playAgain_W(13, 133) <= 0; playAgain_W(13, 134) <= 0; playAgain_W(13, 135) <= 0; playAgain_W(13, 136) <= 1; playAgain_W(13, 137) <= 1; playAgain_W(13, 138) <= 1; playAgain_W(13, 139) <= 1; playAgain_W(13, 140) <= 0; playAgain_W(13, 141) <= 0; playAgain_W(13, 142) <= 0; playAgain_W(13, 143) <= 0; playAgain_W(13, 144) <= 0; playAgain_W(13, 145) <= 0; playAgain_W(13, 146) <= 0; playAgain_W(13, 147) <= 0; playAgain_W(13, 148) <= 0; playAgain_W(13, 149) <= 0; playAgain_W(13, 150) <= 1; playAgain_W(13, 151) <= 1; playAgain_W(13, 152) <= 1; playAgain_W(13, 153) <= 1; playAgain_W(13, 154) <= 0; playAgain_W(13, 155) <= 0; playAgain_W(13, 156) <= 0; playAgain_W(13, 157) <= 0; playAgain_W(13, 158) <= 0; playAgain_W(13, 159) <= 0; playAgain_W(13, 160) <= 0; playAgain_W(13, 161) <= 0; playAgain_W(13, 162) <= 1; playAgain_W(13, 163) <= 1; playAgain_W(13, 164) <= 1; playAgain_W(13, 165) <= 1; playAgain_W(13, 166) <= 0; playAgain_W(13, 167) <= 0; playAgain_W(13, 168) <= 0; playAgain_W(13, 169) <= 0; playAgain_W(13, 170) <= 0; playAgain_W(13, 171) <= 0; playAgain_W(13, 172) <= 1; playAgain_W(13, 173) <= 1; playAgain_W(13, 174) <= 1; playAgain_W(13, 175) <= 1; playAgain_W(13, 176) <= 0; playAgain_W(13, 177) <= 0; playAgain_W(13, 178) <= 0; playAgain_W(13, 179) <= 0; playAgain_W(13, 180) <= 0; playAgain_W(13, 181) <= 0; playAgain_W(13, 182) <= 0; playAgain_W(13, 183) <= 0; playAgain_W(13, 184) <= 0; playAgain_W(13, 185) <= 0; playAgain_W(13, 186) <= 1; playAgain_W(13, 187) <= 1; playAgain_W(13, 188) <= 1; playAgain_W(13, 189) <= 1; playAgain_W(13, 190) <= 0; playAgain_W(13, 191) <= 0; playAgain_W(13, 192) <= 0; playAgain_W(13, 193) <= 0; playAgain_W(13, 194) <= 0; playAgain_W(13, 195) <= 0; playAgain_W(13, 196) <= 0; playAgain_W(13, 197) <= 0; playAgain_W(13, 198) <= 0; playAgain_W(13, 199) <= 0; playAgain_W(13, 200) <= 0; playAgain_W(13, 201) <= 0; playAgain_W(13, 202) <= 0; playAgain_W(13, 203) <= 0; playAgain_W(13, 204) <= 0; playAgain_W(13, 205) <= 0; playAgain_W(13, 206) <= 0; playAgain_W(13, 207) <= 0; playAgain_W(13, 208) <= 0; playAgain_W(13, 209) <= 0; playAgain_W(13, 210) <= 0; playAgain_W(13, 211) <= 0; playAgain_W(13, 212) <= 0; playAgain_W(13, 213) <= 0; playAgain_W(13, 214) <= 0; playAgain_W(13, 215) <= 0; playAgain_W(13, 216) <= 0; playAgain_W(13, 217) <= 0; playAgain_W(13, 218) <= 1; playAgain_W(13, 219) <= 1; playAgain_W(13, 220) <= 1; playAgain_W(13, 221) <= 1; playAgain_W(13, 222) <= 0; playAgain_W(13, 223) <= 0; playAgain_W(13, 224) <= 0; playAgain_W(13, 225) <= 0; playAgain_W(13, 226) <= 1; playAgain_W(13, 227) <= 1; playAgain_W(13, 228) <= 1; playAgain_W(13, 229) <= 1; playAgain_W(13, 230) <= 0; playAgain_W(13, 231) <= 0; playAgain_W(13, 232) <= 0; playAgain_W(13, 233) <= 0; playAgain_W(13, 234) <= 0; playAgain_W(13, 235) <= 0; playAgain_W(13, 236) <= 0; playAgain_W(13, 237) <= 0; playAgain_W(13, 238) <= 0; playAgain_W(13, 239) <= 0; playAgain_W(13, 240) <= 1; playAgain_W(13, 241) <= 1; playAgain_W(13, 242) <= 1; playAgain_W(13, 243) <= 1; playAgain_W(13, 244) <= 0; playAgain_W(13, 245) <= 0; playAgain_W(13, 246) <= 0; playAgain_W(13, 247) <= 0; playAgain_W(13, 248) <= 0; playAgain_W(13, 249) <= 0; playAgain_W(13, 250) <= 0; playAgain_W(13, 251) <= 0; playAgain_W(13, 252) <= 1; playAgain_W(13, 253) <= 1; playAgain_W(13, 254) <= 1; playAgain_W(13, 255) <= 1; playAgain_W(13, 256) <= 0; playAgain_W(13, 257) <= 0; playAgain_W(13, 258) <= 0; playAgain_W(13, 259) <= 0; playAgain_W(13, 260) <= 0; playAgain_W(13, 261) <= 0; playAgain_W(13, 262) <= 1; playAgain_W(13, 263) <= 1; playAgain_W(13, 264) <= 1; playAgain_W(13, 265) <= 1; playAgain_W(13, 266) <= 0; playAgain_W(13, 267) <= 0; playAgain_W(13, 268) <= 0; playAgain_W(13, 269) <= 0; playAgain_W(13, 270) <= 0; playAgain_W(13, 271) <= 0; playAgain_W(13, 272) <= 1; playAgain_W(13, 273) <= 1; playAgain_W(13, 274) <= 1; playAgain_W(13, 275) <= 1; playAgain_W(13, 276) <= 0; playAgain_W(13, 277) <= 0; playAgain_W(13, 278) <= 0; playAgain_W(13, 279) <= 0; playAgain_W(13, 280) <= 1; playAgain_W(13, 281) <= 1; playAgain_W(13, 282) <= 1; playAgain_W(13, 283) <= 1; playAgain_W(13, 284) <= 0; playAgain_W(13, 285) <= 0; playAgain_W(13, 286) <= 0; playAgain_W(13, 287) <= 0; 
playAgain_W(14, 0) <= 0; playAgain_W(14, 1) <= 0; playAgain_W(14, 2) <= 1; playAgain_W(14, 3) <= 1; playAgain_W(14, 4) <= 1; playAgain_W(14, 5) <= 1; playAgain_W(14, 6) <= 0; playAgain_W(14, 7) <= 0; playAgain_W(14, 8) <= 0; playAgain_W(14, 9) <= 0; playAgain_W(14, 10) <= 0; playAgain_W(14, 11) <= 0; playAgain_W(14, 12) <= 0; playAgain_W(14, 13) <= 0; playAgain_W(14, 14) <= 0; playAgain_W(14, 15) <= 0; playAgain_W(14, 16) <= 0; playAgain_W(14, 17) <= 0; playAgain_W(14, 18) <= 0; playAgain_W(14, 19) <= 0; playAgain_W(14, 20) <= 1; playAgain_W(14, 21) <= 1; playAgain_W(14, 22) <= 1; playAgain_W(14, 23) <= 1; playAgain_W(14, 24) <= 0; playAgain_W(14, 25) <= 0; playAgain_W(14, 26) <= 0; playAgain_W(14, 27) <= 0; playAgain_W(14, 28) <= 0; playAgain_W(14, 29) <= 0; playAgain_W(14, 30) <= 1; playAgain_W(14, 31) <= 1; playAgain_W(14, 32) <= 0; playAgain_W(14, 33) <= 0; playAgain_W(14, 34) <= 0; playAgain_W(14, 35) <= 0; playAgain_W(14, 36) <= 1; playAgain_W(14, 37) <= 1; playAgain_W(14, 38) <= 1; playAgain_W(14, 39) <= 1; playAgain_W(14, 40) <= 0; playAgain_W(14, 41) <= 0; playAgain_W(14, 42) <= 0; playAgain_W(14, 43) <= 0; playAgain_W(14, 44) <= 0; playAgain_W(14, 45) <= 0; playAgain_W(14, 46) <= 1; playAgain_W(14, 47) <= 1; playAgain_W(14, 48) <= 1; playAgain_W(14, 49) <= 1; playAgain_W(14, 50) <= 0; playAgain_W(14, 51) <= 0; playAgain_W(14, 52) <= 0; playAgain_W(14, 53) <= 0; playAgain_W(14, 54) <= 0; playAgain_W(14, 55) <= 0; playAgain_W(14, 56) <= 0; playAgain_W(14, 57) <= 0; playAgain_W(14, 58) <= 0; playAgain_W(14, 59) <= 0; playAgain_W(14, 60) <= 1; playAgain_W(14, 61) <= 1; playAgain_W(14, 62) <= 1; playAgain_W(14, 63) <= 1; playAgain_W(14, 64) <= 0; playAgain_W(14, 65) <= 0; playAgain_W(14, 66) <= 0; playAgain_W(14, 67) <= 0; playAgain_W(14, 68) <= 0; playAgain_W(14, 69) <= 0; playAgain_W(14, 70) <= 0; playAgain_W(14, 71) <= 0; playAgain_W(14, 72) <= 0; playAgain_W(14, 73) <= 0; playAgain_W(14, 74) <= 0; playAgain_W(14, 75) <= 0; playAgain_W(14, 76) <= 0; playAgain_W(14, 77) <= 0; playAgain_W(14, 78) <= 0; playAgain_W(14, 79) <= 0; playAgain_W(14, 80) <= 0; playAgain_W(14, 81) <= 0; playAgain_W(14, 82) <= 0; playAgain_W(14, 83) <= 0; playAgain_W(14, 84) <= 0; playAgain_W(14, 85) <= 0; playAgain_W(14, 86) <= 0; playAgain_W(14, 87) <= 0; playAgain_W(14, 88) <= 0; playAgain_W(14, 89) <= 0; playAgain_W(14, 90) <= 1; playAgain_W(14, 91) <= 1; playAgain_W(14, 92) <= 1; playAgain_W(14, 93) <= 1; playAgain_W(14, 94) <= 0; playAgain_W(14, 95) <= 0; playAgain_W(14, 96) <= 0; playAgain_W(14, 97) <= 0; playAgain_W(14, 98) <= 0; playAgain_W(14, 99) <= 0; playAgain_W(14, 100) <= 1; playAgain_W(14, 101) <= 1; playAgain_W(14, 102) <= 1; playAgain_W(14, 103) <= 1; playAgain_W(14, 104) <= 0; playAgain_W(14, 105) <= 0; playAgain_W(14, 106) <= 0; playAgain_W(14, 107) <= 0; playAgain_W(14, 108) <= 1; playAgain_W(14, 109) <= 1; playAgain_W(14, 110) <= 1; playAgain_W(14, 111) <= 1; playAgain_W(14, 112) <= 0; playAgain_W(14, 113) <= 0; playAgain_W(14, 114) <= 0; playAgain_W(14, 115) <= 0; playAgain_W(14, 116) <= 0; playAgain_W(14, 117) <= 0; playAgain_W(14, 118) <= 1; playAgain_W(14, 119) <= 1; playAgain_W(14, 120) <= 1; playAgain_W(14, 121) <= 1; playAgain_W(14, 122) <= 0; playAgain_W(14, 123) <= 0; playAgain_W(14, 124) <= 0; playAgain_W(14, 125) <= 0; playAgain_W(14, 126) <= 1; playAgain_W(14, 127) <= 1; playAgain_W(14, 128) <= 1; playAgain_W(14, 129) <= 1; playAgain_W(14, 130) <= 0; playAgain_W(14, 131) <= 0; playAgain_W(14, 132) <= 0; playAgain_W(14, 133) <= 0; playAgain_W(14, 134) <= 0; playAgain_W(14, 135) <= 0; playAgain_W(14, 136) <= 1; playAgain_W(14, 137) <= 1; playAgain_W(14, 138) <= 1; playAgain_W(14, 139) <= 1; playAgain_W(14, 140) <= 0; playAgain_W(14, 141) <= 0; playAgain_W(14, 142) <= 0; playAgain_W(14, 143) <= 0; playAgain_W(14, 144) <= 0; playAgain_W(14, 145) <= 0; playAgain_W(14, 146) <= 0; playAgain_W(14, 147) <= 0; playAgain_W(14, 148) <= 0; playAgain_W(14, 149) <= 0; playAgain_W(14, 150) <= 1; playAgain_W(14, 151) <= 1; playAgain_W(14, 152) <= 1; playAgain_W(14, 153) <= 1; playAgain_W(14, 154) <= 0; playAgain_W(14, 155) <= 0; playAgain_W(14, 156) <= 0; playAgain_W(14, 157) <= 0; playAgain_W(14, 158) <= 0; playAgain_W(14, 159) <= 0; playAgain_W(14, 160) <= 0; playAgain_W(14, 161) <= 0; playAgain_W(14, 162) <= 1; playAgain_W(14, 163) <= 1; playAgain_W(14, 164) <= 1; playAgain_W(14, 165) <= 1; playAgain_W(14, 166) <= 0; playAgain_W(14, 167) <= 0; playAgain_W(14, 168) <= 0; playAgain_W(14, 169) <= 0; playAgain_W(14, 170) <= 0; playAgain_W(14, 171) <= 0; playAgain_W(14, 172) <= 1; playAgain_W(14, 173) <= 1; playAgain_W(14, 174) <= 1; playAgain_W(14, 175) <= 1; playAgain_W(14, 176) <= 0; playAgain_W(14, 177) <= 0; playAgain_W(14, 178) <= 0; playAgain_W(14, 179) <= 0; playAgain_W(14, 180) <= 0; playAgain_W(14, 181) <= 0; playAgain_W(14, 182) <= 0; playAgain_W(14, 183) <= 0; playAgain_W(14, 184) <= 0; playAgain_W(14, 185) <= 0; playAgain_W(14, 186) <= 1; playAgain_W(14, 187) <= 1; playAgain_W(14, 188) <= 1; playAgain_W(14, 189) <= 1; playAgain_W(14, 190) <= 0; playAgain_W(14, 191) <= 0; playAgain_W(14, 192) <= 0; playAgain_W(14, 193) <= 0; playAgain_W(14, 194) <= 0; playAgain_W(14, 195) <= 0; playAgain_W(14, 196) <= 0; playAgain_W(14, 197) <= 0; playAgain_W(14, 198) <= 0; playAgain_W(14, 199) <= 0; playAgain_W(14, 200) <= 0; playAgain_W(14, 201) <= 0; playAgain_W(14, 202) <= 0; playAgain_W(14, 203) <= 0; playAgain_W(14, 204) <= 0; playAgain_W(14, 205) <= 0; playAgain_W(14, 206) <= 0; playAgain_W(14, 207) <= 0; playAgain_W(14, 208) <= 0; playAgain_W(14, 209) <= 0; playAgain_W(14, 210) <= 0; playAgain_W(14, 211) <= 0; playAgain_W(14, 212) <= 0; playAgain_W(14, 213) <= 0; playAgain_W(14, 214) <= 0; playAgain_W(14, 215) <= 0; playAgain_W(14, 216) <= 0; playAgain_W(14, 217) <= 0; playAgain_W(14, 218) <= 1; playAgain_W(14, 219) <= 1; playAgain_W(14, 220) <= 1; playAgain_W(14, 221) <= 1; playAgain_W(14, 222) <= 0; playAgain_W(14, 223) <= 0; playAgain_W(14, 224) <= 0; playAgain_W(14, 225) <= 0; playAgain_W(14, 226) <= 1; playAgain_W(14, 227) <= 1; playAgain_W(14, 228) <= 1; playAgain_W(14, 229) <= 1; playAgain_W(14, 230) <= 0; playAgain_W(14, 231) <= 0; playAgain_W(14, 232) <= 0; playAgain_W(14, 233) <= 0; playAgain_W(14, 234) <= 0; playAgain_W(14, 235) <= 0; playAgain_W(14, 236) <= 0; playAgain_W(14, 237) <= 0; playAgain_W(14, 238) <= 0; playAgain_W(14, 239) <= 0; playAgain_W(14, 240) <= 1; playAgain_W(14, 241) <= 1; playAgain_W(14, 242) <= 1; playAgain_W(14, 243) <= 1; playAgain_W(14, 244) <= 0; playAgain_W(14, 245) <= 0; playAgain_W(14, 246) <= 0; playAgain_W(14, 247) <= 0; playAgain_W(14, 248) <= 0; playAgain_W(14, 249) <= 0; playAgain_W(14, 250) <= 0; playAgain_W(14, 251) <= 0; playAgain_W(14, 252) <= 1; playAgain_W(14, 253) <= 1; playAgain_W(14, 254) <= 1; playAgain_W(14, 255) <= 1; playAgain_W(14, 256) <= 0; playAgain_W(14, 257) <= 0; playAgain_W(14, 258) <= 0; playAgain_W(14, 259) <= 0; playAgain_W(14, 260) <= 0; playAgain_W(14, 261) <= 0; playAgain_W(14, 262) <= 1; playAgain_W(14, 263) <= 1; playAgain_W(14, 264) <= 1; playAgain_W(14, 265) <= 1; playAgain_W(14, 266) <= 0; playAgain_W(14, 267) <= 0; playAgain_W(14, 268) <= 0; playAgain_W(14, 269) <= 0; playAgain_W(14, 270) <= 0; playAgain_W(14, 271) <= 0; playAgain_W(14, 272) <= 1; playAgain_W(14, 273) <= 1; playAgain_W(14, 274) <= 1; playAgain_W(14, 275) <= 1; playAgain_W(14, 276) <= 0; playAgain_W(14, 277) <= 0; playAgain_W(14, 278) <= 0; playAgain_W(14, 279) <= 0; playAgain_W(14, 280) <= 1; playAgain_W(14, 281) <= 1; playAgain_W(14, 282) <= 1; playAgain_W(14, 283) <= 1; playAgain_W(14, 284) <= 0; playAgain_W(14, 285) <= 0; playAgain_W(14, 286) <= 0; playAgain_W(14, 287) <= 0; 
playAgain_W(15, 0) <= 0; playAgain_W(15, 1) <= 0; playAgain_W(15, 2) <= 1; playAgain_W(15, 3) <= 1; playAgain_W(15, 4) <= 1; playAgain_W(15, 5) <= 1; playAgain_W(15, 6) <= 0; playAgain_W(15, 7) <= 0; playAgain_W(15, 8) <= 0; playAgain_W(15, 9) <= 0; playAgain_W(15, 10) <= 0; playAgain_W(15, 11) <= 0; playAgain_W(15, 12) <= 0; playAgain_W(15, 13) <= 0; playAgain_W(15, 14) <= 0; playAgain_W(15, 15) <= 0; playAgain_W(15, 16) <= 0; playAgain_W(15, 17) <= 0; playAgain_W(15, 18) <= 0; playAgain_W(15, 19) <= 0; playAgain_W(15, 20) <= 1; playAgain_W(15, 21) <= 1; playAgain_W(15, 22) <= 1; playAgain_W(15, 23) <= 1; playAgain_W(15, 24) <= 0; playAgain_W(15, 25) <= 0; playAgain_W(15, 26) <= 0; playAgain_W(15, 27) <= 0; playAgain_W(15, 28) <= 0; playAgain_W(15, 29) <= 0; playAgain_W(15, 30) <= 1; playAgain_W(15, 31) <= 1; playAgain_W(15, 32) <= 0; playAgain_W(15, 33) <= 0; playAgain_W(15, 34) <= 0; playAgain_W(15, 35) <= 0; playAgain_W(15, 36) <= 1; playAgain_W(15, 37) <= 1; playAgain_W(15, 38) <= 1; playAgain_W(15, 39) <= 1; playAgain_W(15, 40) <= 0; playAgain_W(15, 41) <= 0; playAgain_W(15, 42) <= 0; playAgain_W(15, 43) <= 0; playAgain_W(15, 44) <= 0; playAgain_W(15, 45) <= 0; playAgain_W(15, 46) <= 1; playAgain_W(15, 47) <= 1; playAgain_W(15, 48) <= 1; playAgain_W(15, 49) <= 1; playAgain_W(15, 50) <= 0; playAgain_W(15, 51) <= 0; playAgain_W(15, 52) <= 0; playAgain_W(15, 53) <= 0; playAgain_W(15, 54) <= 0; playAgain_W(15, 55) <= 0; playAgain_W(15, 56) <= 0; playAgain_W(15, 57) <= 0; playAgain_W(15, 58) <= 0; playAgain_W(15, 59) <= 0; playAgain_W(15, 60) <= 1; playAgain_W(15, 61) <= 1; playAgain_W(15, 62) <= 1; playAgain_W(15, 63) <= 1; playAgain_W(15, 64) <= 0; playAgain_W(15, 65) <= 0; playAgain_W(15, 66) <= 0; playAgain_W(15, 67) <= 0; playAgain_W(15, 68) <= 0; playAgain_W(15, 69) <= 0; playAgain_W(15, 70) <= 0; playAgain_W(15, 71) <= 0; playAgain_W(15, 72) <= 0; playAgain_W(15, 73) <= 0; playAgain_W(15, 74) <= 0; playAgain_W(15, 75) <= 0; playAgain_W(15, 76) <= 0; playAgain_W(15, 77) <= 0; playAgain_W(15, 78) <= 0; playAgain_W(15, 79) <= 0; playAgain_W(15, 80) <= 0; playAgain_W(15, 81) <= 0; playAgain_W(15, 82) <= 0; playAgain_W(15, 83) <= 0; playAgain_W(15, 84) <= 0; playAgain_W(15, 85) <= 0; playAgain_W(15, 86) <= 0; playAgain_W(15, 87) <= 0; playAgain_W(15, 88) <= 0; playAgain_W(15, 89) <= 0; playAgain_W(15, 90) <= 1; playAgain_W(15, 91) <= 1; playAgain_W(15, 92) <= 1; playAgain_W(15, 93) <= 1; playAgain_W(15, 94) <= 0; playAgain_W(15, 95) <= 0; playAgain_W(15, 96) <= 0; playAgain_W(15, 97) <= 0; playAgain_W(15, 98) <= 0; playAgain_W(15, 99) <= 0; playAgain_W(15, 100) <= 1; playAgain_W(15, 101) <= 1; playAgain_W(15, 102) <= 1; playAgain_W(15, 103) <= 1; playAgain_W(15, 104) <= 0; playAgain_W(15, 105) <= 0; playAgain_W(15, 106) <= 0; playAgain_W(15, 107) <= 0; playAgain_W(15, 108) <= 1; playAgain_W(15, 109) <= 1; playAgain_W(15, 110) <= 1; playAgain_W(15, 111) <= 1; playAgain_W(15, 112) <= 0; playAgain_W(15, 113) <= 0; playAgain_W(15, 114) <= 0; playAgain_W(15, 115) <= 0; playAgain_W(15, 116) <= 0; playAgain_W(15, 117) <= 0; playAgain_W(15, 118) <= 1; playAgain_W(15, 119) <= 1; playAgain_W(15, 120) <= 1; playAgain_W(15, 121) <= 1; playAgain_W(15, 122) <= 0; playAgain_W(15, 123) <= 0; playAgain_W(15, 124) <= 0; playAgain_W(15, 125) <= 0; playAgain_W(15, 126) <= 1; playAgain_W(15, 127) <= 1; playAgain_W(15, 128) <= 1; playAgain_W(15, 129) <= 1; playAgain_W(15, 130) <= 0; playAgain_W(15, 131) <= 0; playAgain_W(15, 132) <= 0; playAgain_W(15, 133) <= 0; playAgain_W(15, 134) <= 0; playAgain_W(15, 135) <= 0; playAgain_W(15, 136) <= 1; playAgain_W(15, 137) <= 1; playAgain_W(15, 138) <= 1; playAgain_W(15, 139) <= 1; playAgain_W(15, 140) <= 0; playAgain_W(15, 141) <= 0; playAgain_W(15, 142) <= 0; playAgain_W(15, 143) <= 0; playAgain_W(15, 144) <= 0; playAgain_W(15, 145) <= 0; playAgain_W(15, 146) <= 0; playAgain_W(15, 147) <= 0; playAgain_W(15, 148) <= 0; playAgain_W(15, 149) <= 0; playAgain_W(15, 150) <= 1; playAgain_W(15, 151) <= 1; playAgain_W(15, 152) <= 1; playAgain_W(15, 153) <= 1; playAgain_W(15, 154) <= 0; playAgain_W(15, 155) <= 0; playAgain_W(15, 156) <= 0; playAgain_W(15, 157) <= 0; playAgain_W(15, 158) <= 0; playAgain_W(15, 159) <= 0; playAgain_W(15, 160) <= 0; playAgain_W(15, 161) <= 0; playAgain_W(15, 162) <= 1; playAgain_W(15, 163) <= 1; playAgain_W(15, 164) <= 1; playAgain_W(15, 165) <= 1; playAgain_W(15, 166) <= 0; playAgain_W(15, 167) <= 0; playAgain_W(15, 168) <= 0; playAgain_W(15, 169) <= 0; playAgain_W(15, 170) <= 0; playAgain_W(15, 171) <= 0; playAgain_W(15, 172) <= 1; playAgain_W(15, 173) <= 1; playAgain_W(15, 174) <= 1; playAgain_W(15, 175) <= 1; playAgain_W(15, 176) <= 0; playAgain_W(15, 177) <= 0; playAgain_W(15, 178) <= 0; playAgain_W(15, 179) <= 0; playAgain_W(15, 180) <= 0; playAgain_W(15, 181) <= 0; playAgain_W(15, 182) <= 0; playAgain_W(15, 183) <= 0; playAgain_W(15, 184) <= 0; playAgain_W(15, 185) <= 0; playAgain_W(15, 186) <= 1; playAgain_W(15, 187) <= 1; playAgain_W(15, 188) <= 1; playAgain_W(15, 189) <= 1; playAgain_W(15, 190) <= 0; playAgain_W(15, 191) <= 0; playAgain_W(15, 192) <= 0; playAgain_W(15, 193) <= 0; playAgain_W(15, 194) <= 0; playAgain_W(15, 195) <= 0; playAgain_W(15, 196) <= 0; playAgain_W(15, 197) <= 0; playAgain_W(15, 198) <= 0; playAgain_W(15, 199) <= 0; playAgain_W(15, 200) <= 0; playAgain_W(15, 201) <= 0; playAgain_W(15, 202) <= 0; playAgain_W(15, 203) <= 0; playAgain_W(15, 204) <= 0; playAgain_W(15, 205) <= 0; playAgain_W(15, 206) <= 0; playAgain_W(15, 207) <= 0; playAgain_W(15, 208) <= 0; playAgain_W(15, 209) <= 0; playAgain_W(15, 210) <= 0; playAgain_W(15, 211) <= 0; playAgain_W(15, 212) <= 0; playAgain_W(15, 213) <= 0; playAgain_W(15, 214) <= 0; playAgain_W(15, 215) <= 0; playAgain_W(15, 216) <= 0; playAgain_W(15, 217) <= 0; playAgain_W(15, 218) <= 1; playAgain_W(15, 219) <= 1; playAgain_W(15, 220) <= 1; playAgain_W(15, 221) <= 1; playAgain_W(15, 222) <= 0; playAgain_W(15, 223) <= 0; playAgain_W(15, 224) <= 0; playAgain_W(15, 225) <= 0; playAgain_W(15, 226) <= 1; playAgain_W(15, 227) <= 1; playAgain_W(15, 228) <= 1; playAgain_W(15, 229) <= 1; playAgain_W(15, 230) <= 0; playAgain_W(15, 231) <= 0; playAgain_W(15, 232) <= 0; playAgain_W(15, 233) <= 0; playAgain_W(15, 234) <= 0; playAgain_W(15, 235) <= 0; playAgain_W(15, 236) <= 0; playAgain_W(15, 237) <= 0; playAgain_W(15, 238) <= 0; playAgain_W(15, 239) <= 0; playAgain_W(15, 240) <= 1; playAgain_W(15, 241) <= 1; playAgain_W(15, 242) <= 1; playAgain_W(15, 243) <= 1; playAgain_W(15, 244) <= 0; playAgain_W(15, 245) <= 0; playAgain_W(15, 246) <= 0; playAgain_W(15, 247) <= 0; playAgain_W(15, 248) <= 0; playAgain_W(15, 249) <= 0; playAgain_W(15, 250) <= 0; playAgain_W(15, 251) <= 0; playAgain_W(15, 252) <= 1; playAgain_W(15, 253) <= 1; playAgain_W(15, 254) <= 1; playAgain_W(15, 255) <= 1; playAgain_W(15, 256) <= 0; playAgain_W(15, 257) <= 0; playAgain_W(15, 258) <= 0; playAgain_W(15, 259) <= 0; playAgain_W(15, 260) <= 0; playAgain_W(15, 261) <= 0; playAgain_W(15, 262) <= 1; playAgain_W(15, 263) <= 1; playAgain_W(15, 264) <= 1; playAgain_W(15, 265) <= 1; playAgain_W(15, 266) <= 0; playAgain_W(15, 267) <= 0; playAgain_W(15, 268) <= 0; playAgain_W(15, 269) <= 0; playAgain_W(15, 270) <= 0; playAgain_W(15, 271) <= 0; playAgain_W(15, 272) <= 1; playAgain_W(15, 273) <= 1; playAgain_W(15, 274) <= 1; playAgain_W(15, 275) <= 1; playAgain_W(15, 276) <= 0; playAgain_W(15, 277) <= 0; playAgain_W(15, 278) <= 0; playAgain_W(15, 279) <= 0; playAgain_W(15, 280) <= 1; playAgain_W(15, 281) <= 1; playAgain_W(15, 282) <= 1; playAgain_W(15, 283) <= 1; playAgain_W(15, 284) <= 0; playAgain_W(15, 285) <= 0; playAgain_W(15, 286) <= 0; playAgain_W(15, 287) <= 0; 
playAgain_W(16, 0) <= 0; playAgain_W(16, 1) <= 0; playAgain_W(16, 2) <= 1; playAgain_W(16, 3) <= 1; playAgain_W(16, 4) <= 1; playAgain_W(16, 5) <= 1; playAgain_W(16, 6) <= 0; playAgain_W(16, 7) <= 0; playAgain_W(16, 8) <= 0; playAgain_W(16, 9) <= 0; playAgain_W(16, 10) <= 0; playAgain_W(16, 11) <= 0; playAgain_W(16, 12) <= 0; playAgain_W(16, 13) <= 0; playAgain_W(16, 14) <= 0; playAgain_W(16, 15) <= 0; playAgain_W(16, 16) <= 0; playAgain_W(16, 17) <= 0; playAgain_W(16, 18) <= 0; playAgain_W(16, 19) <= 0; playAgain_W(16, 20) <= 1; playAgain_W(16, 21) <= 1; playAgain_W(16, 22) <= 1; playAgain_W(16, 23) <= 1; playAgain_W(16, 24) <= 0; playAgain_W(16, 25) <= 0; playAgain_W(16, 26) <= 0; playAgain_W(16, 27) <= 0; playAgain_W(16, 28) <= 1; playAgain_W(16, 29) <= 1; playAgain_W(16, 30) <= 1; playAgain_W(16, 31) <= 1; playAgain_W(16, 32) <= 0; playAgain_W(16, 33) <= 0; playAgain_W(16, 34) <= 0; playAgain_W(16, 35) <= 0; playAgain_W(16, 36) <= 1; playAgain_W(16, 37) <= 1; playAgain_W(16, 38) <= 1; playAgain_W(16, 39) <= 1; playAgain_W(16, 40) <= 0; playAgain_W(16, 41) <= 0; playAgain_W(16, 42) <= 0; playAgain_W(16, 43) <= 0; playAgain_W(16, 44) <= 0; playAgain_W(16, 45) <= 0; playAgain_W(16, 46) <= 1; playAgain_W(16, 47) <= 1; playAgain_W(16, 48) <= 1; playAgain_W(16, 49) <= 1; playAgain_W(16, 50) <= 0; playAgain_W(16, 51) <= 0; playAgain_W(16, 52) <= 0; playAgain_W(16, 53) <= 0; playAgain_W(16, 54) <= 0; playAgain_W(16, 55) <= 0; playAgain_W(16, 56) <= 0; playAgain_W(16, 57) <= 0; playAgain_W(16, 58) <= 0; playAgain_W(16, 59) <= 0; playAgain_W(16, 60) <= 1; playAgain_W(16, 61) <= 1; playAgain_W(16, 62) <= 1; playAgain_W(16, 63) <= 1; playAgain_W(16, 64) <= 0; playAgain_W(16, 65) <= 0; playAgain_W(16, 66) <= 0; playAgain_W(16, 67) <= 0; playAgain_W(16, 68) <= 0; playAgain_W(16, 69) <= 0; playAgain_W(16, 70) <= 0; playAgain_W(16, 71) <= 0; playAgain_W(16, 72) <= 0; playAgain_W(16, 73) <= 0; playAgain_W(16, 74) <= 0; playAgain_W(16, 75) <= 0; playAgain_W(16, 76) <= 0; playAgain_W(16, 77) <= 0; playAgain_W(16, 78) <= 0; playAgain_W(16, 79) <= 0; playAgain_W(16, 80) <= 0; playAgain_W(16, 81) <= 0; playAgain_W(16, 82) <= 0; playAgain_W(16, 83) <= 0; playAgain_W(16, 84) <= 0; playAgain_W(16, 85) <= 0; playAgain_W(16, 86) <= 0; playAgain_W(16, 87) <= 0; playAgain_W(16, 88) <= 0; playAgain_W(16, 89) <= 0; playAgain_W(16, 90) <= 1; playAgain_W(16, 91) <= 1; playAgain_W(16, 92) <= 1; playAgain_W(16, 93) <= 1; playAgain_W(16, 94) <= 0; playAgain_W(16, 95) <= 0; playAgain_W(16, 96) <= 0; playAgain_W(16, 97) <= 0; playAgain_W(16, 98) <= 0; playAgain_W(16, 99) <= 0; playAgain_W(16, 100) <= 1; playAgain_W(16, 101) <= 1; playAgain_W(16, 102) <= 1; playAgain_W(16, 103) <= 1; playAgain_W(16, 104) <= 0; playAgain_W(16, 105) <= 0; playAgain_W(16, 106) <= 0; playAgain_W(16, 107) <= 0; playAgain_W(16, 108) <= 0; playAgain_W(16, 109) <= 0; playAgain_W(16, 110) <= 1; playAgain_W(16, 111) <= 1; playAgain_W(16, 112) <= 1; playAgain_W(16, 113) <= 1; playAgain_W(16, 114) <= 0; playAgain_W(16, 115) <= 0; playAgain_W(16, 116) <= 0; playAgain_W(16, 117) <= 0; playAgain_W(16, 118) <= 1; playAgain_W(16, 119) <= 1; playAgain_W(16, 120) <= 1; playAgain_W(16, 121) <= 1; playAgain_W(16, 122) <= 0; playAgain_W(16, 123) <= 0; playAgain_W(16, 124) <= 0; playAgain_W(16, 125) <= 0; playAgain_W(16, 126) <= 1; playAgain_W(16, 127) <= 1; playAgain_W(16, 128) <= 1; playAgain_W(16, 129) <= 1; playAgain_W(16, 130) <= 0; playAgain_W(16, 131) <= 0; playAgain_W(16, 132) <= 0; playAgain_W(16, 133) <= 0; playAgain_W(16, 134) <= 0; playAgain_W(16, 135) <= 0; playAgain_W(16, 136) <= 1; playAgain_W(16, 137) <= 1; playAgain_W(16, 138) <= 1; playAgain_W(16, 139) <= 1; playAgain_W(16, 140) <= 0; playAgain_W(16, 141) <= 0; playAgain_W(16, 142) <= 0; playAgain_W(16, 143) <= 0; playAgain_W(16, 144) <= 0; playAgain_W(16, 145) <= 0; playAgain_W(16, 146) <= 0; playAgain_W(16, 147) <= 0; playAgain_W(16, 148) <= 0; playAgain_W(16, 149) <= 0; playAgain_W(16, 150) <= 1; playAgain_W(16, 151) <= 1; playAgain_W(16, 152) <= 1; playAgain_W(16, 153) <= 1; playAgain_W(16, 154) <= 0; playAgain_W(16, 155) <= 0; playAgain_W(16, 156) <= 0; playAgain_W(16, 157) <= 0; playAgain_W(16, 158) <= 0; playAgain_W(16, 159) <= 0; playAgain_W(16, 160) <= 0; playAgain_W(16, 161) <= 0; playAgain_W(16, 162) <= 1; playAgain_W(16, 163) <= 1; playAgain_W(16, 164) <= 1; playAgain_W(16, 165) <= 1; playAgain_W(16, 166) <= 0; playAgain_W(16, 167) <= 0; playAgain_W(16, 168) <= 0; playAgain_W(16, 169) <= 0; playAgain_W(16, 170) <= 0; playAgain_W(16, 171) <= 0; playAgain_W(16, 172) <= 1; playAgain_W(16, 173) <= 1; playAgain_W(16, 174) <= 1; playAgain_W(16, 175) <= 1; playAgain_W(16, 176) <= 0; playAgain_W(16, 177) <= 0; playAgain_W(16, 178) <= 0; playAgain_W(16, 179) <= 0; playAgain_W(16, 180) <= 0; playAgain_W(16, 181) <= 0; playAgain_W(16, 182) <= 0; playAgain_W(16, 183) <= 0; playAgain_W(16, 184) <= 0; playAgain_W(16, 185) <= 0; playAgain_W(16, 186) <= 0; playAgain_W(16, 187) <= 0; playAgain_W(16, 188) <= 0; playAgain_W(16, 189) <= 0; playAgain_W(16, 190) <= 0; playAgain_W(16, 191) <= 0; playAgain_W(16, 192) <= 0; playAgain_W(16, 193) <= 0; playAgain_W(16, 194) <= 0; playAgain_W(16, 195) <= 0; playAgain_W(16, 196) <= 0; playAgain_W(16, 197) <= 0; playAgain_W(16, 198) <= 0; playAgain_W(16, 199) <= 0; playAgain_W(16, 200) <= 0; playAgain_W(16, 201) <= 0; playAgain_W(16, 202) <= 0; playAgain_W(16, 203) <= 0; playAgain_W(16, 204) <= 0; playAgain_W(16, 205) <= 0; playAgain_W(16, 206) <= 0; playAgain_W(16, 207) <= 0; playAgain_W(16, 208) <= 0; playAgain_W(16, 209) <= 0; playAgain_W(16, 210) <= 0; playAgain_W(16, 211) <= 0; playAgain_W(16, 212) <= 0; playAgain_W(16, 213) <= 0; playAgain_W(16, 214) <= 0; playAgain_W(16, 215) <= 0; playAgain_W(16, 216) <= 0; playAgain_W(16, 217) <= 0; playAgain_W(16, 218) <= 1; playAgain_W(16, 219) <= 1; playAgain_W(16, 220) <= 1; playAgain_W(16, 221) <= 1; playAgain_W(16, 222) <= 0; playAgain_W(16, 223) <= 0; playAgain_W(16, 224) <= 0; playAgain_W(16, 225) <= 0; playAgain_W(16, 226) <= 1; playAgain_W(16, 227) <= 1; playAgain_W(16, 228) <= 1; playAgain_W(16, 229) <= 1; playAgain_W(16, 230) <= 0; playAgain_W(16, 231) <= 0; playAgain_W(16, 232) <= 0; playAgain_W(16, 233) <= 0; playAgain_W(16, 234) <= 0; playAgain_W(16, 235) <= 0; playAgain_W(16, 236) <= 0; playAgain_W(16, 237) <= 0; playAgain_W(16, 238) <= 0; playAgain_W(16, 239) <= 0; playAgain_W(16, 240) <= 1; playAgain_W(16, 241) <= 1; playAgain_W(16, 242) <= 1; playAgain_W(16, 243) <= 1; playAgain_W(16, 244) <= 0; playAgain_W(16, 245) <= 0; playAgain_W(16, 246) <= 0; playAgain_W(16, 247) <= 0; playAgain_W(16, 248) <= 0; playAgain_W(16, 249) <= 0; playAgain_W(16, 250) <= 0; playAgain_W(16, 251) <= 0; playAgain_W(16, 252) <= 1; playAgain_W(16, 253) <= 1; playAgain_W(16, 254) <= 1; playAgain_W(16, 255) <= 1; playAgain_W(16, 256) <= 0; playAgain_W(16, 257) <= 0; playAgain_W(16, 258) <= 0; playAgain_W(16, 259) <= 0; playAgain_W(16, 260) <= 0; playAgain_W(16, 261) <= 0; playAgain_W(16, 262) <= 1; playAgain_W(16, 263) <= 1; playAgain_W(16, 264) <= 1; playAgain_W(16, 265) <= 1; playAgain_W(16, 266) <= 0; playAgain_W(16, 267) <= 0; playAgain_W(16, 268) <= 0; playAgain_W(16, 269) <= 0; playAgain_W(16, 270) <= 0; playAgain_W(16, 271) <= 0; playAgain_W(16, 272) <= 1; playAgain_W(16, 273) <= 1; playAgain_W(16, 274) <= 1; playAgain_W(16, 275) <= 1; playAgain_W(16, 276) <= 0; playAgain_W(16, 277) <= 0; playAgain_W(16, 278) <= 1; playAgain_W(16, 279) <= 1; playAgain_W(16, 280) <= 1; playAgain_W(16, 281) <= 1; playAgain_W(16, 282) <= 0; playAgain_W(16, 283) <= 0; playAgain_W(16, 284) <= 0; playAgain_W(16, 285) <= 0; playAgain_W(16, 286) <= 0; playAgain_W(16, 287) <= 0; 
playAgain_W(17, 0) <= 0; playAgain_W(17, 1) <= 0; playAgain_W(17, 2) <= 1; playAgain_W(17, 3) <= 1; playAgain_W(17, 4) <= 1; playAgain_W(17, 5) <= 1; playAgain_W(17, 6) <= 0; playAgain_W(17, 7) <= 0; playAgain_W(17, 8) <= 0; playAgain_W(17, 9) <= 0; playAgain_W(17, 10) <= 0; playAgain_W(17, 11) <= 0; playAgain_W(17, 12) <= 0; playAgain_W(17, 13) <= 0; playAgain_W(17, 14) <= 0; playAgain_W(17, 15) <= 0; playAgain_W(17, 16) <= 0; playAgain_W(17, 17) <= 0; playAgain_W(17, 18) <= 0; playAgain_W(17, 19) <= 0; playAgain_W(17, 20) <= 1; playAgain_W(17, 21) <= 1; playAgain_W(17, 22) <= 1; playAgain_W(17, 23) <= 1; playAgain_W(17, 24) <= 0; playAgain_W(17, 25) <= 0; playAgain_W(17, 26) <= 0; playAgain_W(17, 27) <= 0; playAgain_W(17, 28) <= 1; playAgain_W(17, 29) <= 1; playAgain_W(17, 30) <= 1; playAgain_W(17, 31) <= 1; playAgain_W(17, 32) <= 0; playAgain_W(17, 33) <= 0; playAgain_W(17, 34) <= 0; playAgain_W(17, 35) <= 0; playAgain_W(17, 36) <= 1; playAgain_W(17, 37) <= 1; playAgain_W(17, 38) <= 1; playAgain_W(17, 39) <= 1; playAgain_W(17, 40) <= 0; playAgain_W(17, 41) <= 0; playAgain_W(17, 42) <= 0; playAgain_W(17, 43) <= 0; playAgain_W(17, 44) <= 0; playAgain_W(17, 45) <= 0; playAgain_W(17, 46) <= 1; playAgain_W(17, 47) <= 1; playAgain_W(17, 48) <= 1; playAgain_W(17, 49) <= 1; playAgain_W(17, 50) <= 0; playAgain_W(17, 51) <= 0; playAgain_W(17, 52) <= 0; playAgain_W(17, 53) <= 0; playAgain_W(17, 54) <= 0; playAgain_W(17, 55) <= 0; playAgain_W(17, 56) <= 0; playAgain_W(17, 57) <= 0; playAgain_W(17, 58) <= 0; playAgain_W(17, 59) <= 0; playAgain_W(17, 60) <= 1; playAgain_W(17, 61) <= 1; playAgain_W(17, 62) <= 1; playAgain_W(17, 63) <= 1; playAgain_W(17, 64) <= 0; playAgain_W(17, 65) <= 0; playAgain_W(17, 66) <= 0; playAgain_W(17, 67) <= 0; playAgain_W(17, 68) <= 0; playAgain_W(17, 69) <= 0; playAgain_W(17, 70) <= 0; playAgain_W(17, 71) <= 0; playAgain_W(17, 72) <= 0; playAgain_W(17, 73) <= 0; playAgain_W(17, 74) <= 0; playAgain_W(17, 75) <= 0; playAgain_W(17, 76) <= 0; playAgain_W(17, 77) <= 0; playAgain_W(17, 78) <= 0; playAgain_W(17, 79) <= 0; playAgain_W(17, 80) <= 0; playAgain_W(17, 81) <= 0; playAgain_W(17, 82) <= 0; playAgain_W(17, 83) <= 0; playAgain_W(17, 84) <= 0; playAgain_W(17, 85) <= 0; playAgain_W(17, 86) <= 0; playAgain_W(17, 87) <= 0; playAgain_W(17, 88) <= 0; playAgain_W(17, 89) <= 0; playAgain_W(17, 90) <= 1; playAgain_W(17, 91) <= 1; playAgain_W(17, 92) <= 1; playAgain_W(17, 93) <= 1; playAgain_W(17, 94) <= 0; playAgain_W(17, 95) <= 0; playAgain_W(17, 96) <= 0; playAgain_W(17, 97) <= 0; playAgain_W(17, 98) <= 0; playAgain_W(17, 99) <= 0; playAgain_W(17, 100) <= 1; playAgain_W(17, 101) <= 1; playAgain_W(17, 102) <= 1; playAgain_W(17, 103) <= 1; playAgain_W(17, 104) <= 0; playAgain_W(17, 105) <= 0; playAgain_W(17, 106) <= 0; playAgain_W(17, 107) <= 0; playAgain_W(17, 108) <= 0; playAgain_W(17, 109) <= 0; playAgain_W(17, 110) <= 1; playAgain_W(17, 111) <= 1; playAgain_W(17, 112) <= 1; playAgain_W(17, 113) <= 1; playAgain_W(17, 114) <= 0; playAgain_W(17, 115) <= 0; playAgain_W(17, 116) <= 0; playAgain_W(17, 117) <= 0; playAgain_W(17, 118) <= 1; playAgain_W(17, 119) <= 1; playAgain_W(17, 120) <= 1; playAgain_W(17, 121) <= 1; playAgain_W(17, 122) <= 0; playAgain_W(17, 123) <= 0; playAgain_W(17, 124) <= 0; playAgain_W(17, 125) <= 0; playAgain_W(17, 126) <= 1; playAgain_W(17, 127) <= 1; playAgain_W(17, 128) <= 1; playAgain_W(17, 129) <= 1; playAgain_W(17, 130) <= 0; playAgain_W(17, 131) <= 0; playAgain_W(17, 132) <= 0; playAgain_W(17, 133) <= 0; playAgain_W(17, 134) <= 0; playAgain_W(17, 135) <= 0; playAgain_W(17, 136) <= 1; playAgain_W(17, 137) <= 1; playAgain_W(17, 138) <= 1; playAgain_W(17, 139) <= 1; playAgain_W(17, 140) <= 0; playAgain_W(17, 141) <= 0; playAgain_W(17, 142) <= 0; playAgain_W(17, 143) <= 0; playAgain_W(17, 144) <= 0; playAgain_W(17, 145) <= 0; playAgain_W(17, 146) <= 0; playAgain_W(17, 147) <= 0; playAgain_W(17, 148) <= 0; playAgain_W(17, 149) <= 0; playAgain_W(17, 150) <= 1; playAgain_W(17, 151) <= 1; playAgain_W(17, 152) <= 1; playAgain_W(17, 153) <= 1; playAgain_W(17, 154) <= 0; playAgain_W(17, 155) <= 0; playAgain_W(17, 156) <= 0; playAgain_W(17, 157) <= 0; playAgain_W(17, 158) <= 0; playAgain_W(17, 159) <= 0; playAgain_W(17, 160) <= 0; playAgain_W(17, 161) <= 0; playAgain_W(17, 162) <= 1; playAgain_W(17, 163) <= 1; playAgain_W(17, 164) <= 1; playAgain_W(17, 165) <= 1; playAgain_W(17, 166) <= 0; playAgain_W(17, 167) <= 0; playAgain_W(17, 168) <= 0; playAgain_W(17, 169) <= 0; playAgain_W(17, 170) <= 0; playAgain_W(17, 171) <= 0; playAgain_W(17, 172) <= 1; playAgain_W(17, 173) <= 1; playAgain_W(17, 174) <= 1; playAgain_W(17, 175) <= 1; playAgain_W(17, 176) <= 0; playAgain_W(17, 177) <= 0; playAgain_W(17, 178) <= 0; playAgain_W(17, 179) <= 0; playAgain_W(17, 180) <= 0; playAgain_W(17, 181) <= 0; playAgain_W(17, 182) <= 0; playAgain_W(17, 183) <= 0; playAgain_W(17, 184) <= 0; playAgain_W(17, 185) <= 0; playAgain_W(17, 186) <= 0; playAgain_W(17, 187) <= 0; playAgain_W(17, 188) <= 0; playAgain_W(17, 189) <= 0; playAgain_W(17, 190) <= 0; playAgain_W(17, 191) <= 0; playAgain_W(17, 192) <= 0; playAgain_W(17, 193) <= 0; playAgain_W(17, 194) <= 0; playAgain_W(17, 195) <= 0; playAgain_W(17, 196) <= 0; playAgain_W(17, 197) <= 0; playAgain_W(17, 198) <= 0; playAgain_W(17, 199) <= 0; playAgain_W(17, 200) <= 0; playAgain_W(17, 201) <= 0; playAgain_W(17, 202) <= 0; playAgain_W(17, 203) <= 0; playAgain_W(17, 204) <= 0; playAgain_W(17, 205) <= 0; playAgain_W(17, 206) <= 0; playAgain_W(17, 207) <= 0; playAgain_W(17, 208) <= 0; playAgain_W(17, 209) <= 0; playAgain_W(17, 210) <= 0; playAgain_W(17, 211) <= 0; playAgain_W(17, 212) <= 0; playAgain_W(17, 213) <= 0; playAgain_W(17, 214) <= 0; playAgain_W(17, 215) <= 0; playAgain_W(17, 216) <= 0; playAgain_W(17, 217) <= 0; playAgain_W(17, 218) <= 1; playAgain_W(17, 219) <= 1; playAgain_W(17, 220) <= 1; playAgain_W(17, 221) <= 1; playAgain_W(17, 222) <= 0; playAgain_W(17, 223) <= 0; playAgain_W(17, 224) <= 0; playAgain_W(17, 225) <= 0; playAgain_W(17, 226) <= 1; playAgain_W(17, 227) <= 1; playAgain_W(17, 228) <= 1; playAgain_W(17, 229) <= 1; playAgain_W(17, 230) <= 0; playAgain_W(17, 231) <= 0; playAgain_W(17, 232) <= 0; playAgain_W(17, 233) <= 0; playAgain_W(17, 234) <= 0; playAgain_W(17, 235) <= 0; playAgain_W(17, 236) <= 0; playAgain_W(17, 237) <= 0; playAgain_W(17, 238) <= 0; playAgain_W(17, 239) <= 0; playAgain_W(17, 240) <= 1; playAgain_W(17, 241) <= 1; playAgain_W(17, 242) <= 1; playAgain_W(17, 243) <= 1; playAgain_W(17, 244) <= 0; playAgain_W(17, 245) <= 0; playAgain_W(17, 246) <= 0; playAgain_W(17, 247) <= 0; playAgain_W(17, 248) <= 0; playAgain_W(17, 249) <= 0; playAgain_W(17, 250) <= 0; playAgain_W(17, 251) <= 0; playAgain_W(17, 252) <= 1; playAgain_W(17, 253) <= 1; playAgain_W(17, 254) <= 1; playAgain_W(17, 255) <= 1; playAgain_W(17, 256) <= 0; playAgain_W(17, 257) <= 0; playAgain_W(17, 258) <= 0; playAgain_W(17, 259) <= 0; playAgain_W(17, 260) <= 0; playAgain_W(17, 261) <= 0; playAgain_W(17, 262) <= 1; playAgain_W(17, 263) <= 1; playAgain_W(17, 264) <= 1; playAgain_W(17, 265) <= 1; playAgain_W(17, 266) <= 0; playAgain_W(17, 267) <= 0; playAgain_W(17, 268) <= 0; playAgain_W(17, 269) <= 0; playAgain_W(17, 270) <= 0; playAgain_W(17, 271) <= 0; playAgain_W(17, 272) <= 1; playAgain_W(17, 273) <= 1; playAgain_W(17, 274) <= 1; playAgain_W(17, 275) <= 1; playAgain_W(17, 276) <= 0; playAgain_W(17, 277) <= 0; playAgain_W(17, 278) <= 1; playAgain_W(17, 279) <= 1; playAgain_W(17, 280) <= 1; playAgain_W(17, 281) <= 1; playAgain_W(17, 282) <= 0; playAgain_W(17, 283) <= 0; playAgain_W(17, 284) <= 0; playAgain_W(17, 285) <= 0; playAgain_W(17, 286) <= 0; playAgain_W(17, 287) <= 0; 
playAgain_W(18, 0) <= 1; playAgain_W(18, 1) <= 1; playAgain_W(18, 2) <= 1; playAgain_W(18, 3) <= 1; playAgain_W(18, 4) <= 1; playAgain_W(18, 5) <= 1; playAgain_W(18, 6) <= 1; playAgain_W(18, 7) <= 1; playAgain_W(18, 8) <= 0; playAgain_W(18, 9) <= 0; playAgain_W(18, 10) <= 0; playAgain_W(18, 11) <= 0; playAgain_W(18, 12) <= 0; playAgain_W(18, 13) <= 0; playAgain_W(18, 14) <= 0; playAgain_W(18, 15) <= 0; playAgain_W(18, 16) <= 0; playAgain_W(18, 17) <= 0; playAgain_W(18, 18) <= 1; playAgain_W(18, 19) <= 1; playAgain_W(18, 20) <= 1; playAgain_W(18, 21) <= 1; playAgain_W(18, 22) <= 1; playAgain_W(18, 23) <= 1; playAgain_W(18, 24) <= 1; playAgain_W(18, 25) <= 1; playAgain_W(18, 26) <= 1; playAgain_W(18, 27) <= 1; playAgain_W(18, 28) <= 1; playAgain_W(18, 29) <= 1; playAgain_W(18, 30) <= 1; playAgain_W(18, 31) <= 1; playAgain_W(18, 32) <= 0; playAgain_W(18, 33) <= 0; playAgain_W(18, 34) <= 0; playAgain_W(18, 35) <= 0; playAgain_W(18, 36) <= 1; playAgain_W(18, 37) <= 1; playAgain_W(18, 38) <= 1; playAgain_W(18, 39) <= 1; playAgain_W(18, 40) <= 0; playAgain_W(18, 41) <= 0; playAgain_W(18, 42) <= 0; playAgain_W(18, 43) <= 0; playAgain_W(18, 44) <= 0; playAgain_W(18, 45) <= 0; playAgain_W(18, 46) <= 1; playAgain_W(18, 47) <= 1; playAgain_W(18, 48) <= 1; playAgain_W(18, 49) <= 1; playAgain_W(18, 50) <= 0; playAgain_W(18, 51) <= 0; playAgain_W(18, 52) <= 0; playAgain_W(18, 53) <= 0; playAgain_W(18, 54) <= 0; playAgain_W(18, 55) <= 0; playAgain_W(18, 56) <= 0; playAgain_W(18, 57) <= 0; playAgain_W(18, 58) <= 1; playAgain_W(18, 59) <= 1; playAgain_W(18, 60) <= 1; playAgain_W(18, 61) <= 1; playAgain_W(18, 62) <= 1; playAgain_W(18, 63) <= 1; playAgain_W(18, 64) <= 1; playAgain_W(18, 65) <= 1; playAgain_W(18, 66) <= 0; playAgain_W(18, 67) <= 0; playAgain_W(18, 68) <= 0; playAgain_W(18, 69) <= 0; playAgain_W(18, 70) <= 0; playAgain_W(18, 71) <= 0; playAgain_W(18, 72) <= 0; playAgain_W(18, 73) <= 0; playAgain_W(18, 74) <= 0; playAgain_W(18, 75) <= 0; playAgain_W(18, 76) <= 0; playAgain_W(18, 77) <= 0; playAgain_W(18, 78) <= 0; playAgain_W(18, 79) <= 0; playAgain_W(18, 80) <= 0; playAgain_W(18, 81) <= 0; playAgain_W(18, 82) <= 0; playAgain_W(18, 83) <= 0; playAgain_W(18, 84) <= 0; playAgain_W(18, 85) <= 0; playAgain_W(18, 86) <= 0; playAgain_W(18, 87) <= 0; playAgain_W(18, 88) <= 0; playAgain_W(18, 89) <= 0; playAgain_W(18, 90) <= 1; playAgain_W(18, 91) <= 1; playAgain_W(18, 92) <= 1; playAgain_W(18, 93) <= 1; playAgain_W(18, 94) <= 0; playAgain_W(18, 95) <= 0; playAgain_W(18, 96) <= 0; playAgain_W(18, 97) <= 0; playAgain_W(18, 98) <= 0; playAgain_W(18, 99) <= 0; playAgain_W(18, 100) <= 1; playAgain_W(18, 101) <= 1; playAgain_W(18, 102) <= 1; playAgain_W(18, 103) <= 1; playAgain_W(18, 104) <= 0; playAgain_W(18, 105) <= 0; playAgain_W(18, 106) <= 0; playAgain_W(18, 107) <= 0; playAgain_W(18, 108) <= 0; playAgain_W(18, 109) <= 0; playAgain_W(18, 110) <= 0; playAgain_W(18, 111) <= 0; playAgain_W(18, 112) <= 1; playAgain_W(18, 113) <= 1; playAgain_W(18, 114) <= 1; playAgain_W(18, 115) <= 1; playAgain_W(18, 116) <= 1; playAgain_W(18, 117) <= 1; playAgain_W(18, 118) <= 0; playAgain_W(18, 119) <= 0; playAgain_W(18, 120) <= 1; playAgain_W(18, 121) <= 1; playAgain_W(18, 122) <= 0; playAgain_W(18, 123) <= 0; playAgain_W(18, 124) <= 0; playAgain_W(18, 125) <= 0; playAgain_W(18, 126) <= 1; playAgain_W(18, 127) <= 1; playAgain_W(18, 128) <= 1; playAgain_W(18, 129) <= 1; playAgain_W(18, 130) <= 0; playAgain_W(18, 131) <= 0; playAgain_W(18, 132) <= 0; playAgain_W(18, 133) <= 0; playAgain_W(18, 134) <= 0; playAgain_W(18, 135) <= 0; playAgain_W(18, 136) <= 1; playAgain_W(18, 137) <= 1; playAgain_W(18, 138) <= 1; playAgain_W(18, 139) <= 1; playAgain_W(18, 140) <= 0; playAgain_W(18, 141) <= 0; playAgain_W(18, 142) <= 0; playAgain_W(18, 143) <= 0; playAgain_W(18, 144) <= 0; playAgain_W(18, 145) <= 0; playAgain_W(18, 146) <= 0; playAgain_W(18, 147) <= 0; playAgain_W(18, 148) <= 1; playAgain_W(18, 149) <= 1; playAgain_W(18, 150) <= 1; playAgain_W(18, 151) <= 1; playAgain_W(18, 152) <= 1; playAgain_W(18, 153) <= 1; playAgain_W(18, 154) <= 1; playAgain_W(18, 155) <= 1; playAgain_W(18, 156) <= 0; playAgain_W(18, 157) <= 0; playAgain_W(18, 158) <= 0; playAgain_W(18, 159) <= 0; playAgain_W(18, 160) <= 0; playAgain_W(18, 161) <= 0; playAgain_W(18, 162) <= 1; playAgain_W(18, 163) <= 1; playAgain_W(18, 164) <= 1; playAgain_W(18, 165) <= 1; playAgain_W(18, 166) <= 0; playAgain_W(18, 167) <= 0; playAgain_W(18, 168) <= 0; playAgain_W(18, 169) <= 0; playAgain_W(18, 170) <= 0; playAgain_W(18, 171) <= 0; playAgain_W(18, 172) <= 1; playAgain_W(18, 173) <= 1; playAgain_W(18, 174) <= 1; playAgain_W(18, 175) <= 1; playAgain_W(18, 176) <= 0; playAgain_W(18, 177) <= 0; playAgain_W(18, 178) <= 0; playAgain_W(18, 179) <= 0; playAgain_W(18, 180) <= 0; playAgain_W(18, 181) <= 0; playAgain_W(18, 182) <= 0; playAgain_W(18, 183) <= 0; playAgain_W(18, 184) <= 0; playAgain_W(18, 185) <= 0; playAgain_W(18, 186) <= 0; playAgain_W(18, 187) <= 0; playAgain_W(18, 188) <= 0; playAgain_W(18, 189) <= 0; playAgain_W(18, 190) <= 0; playAgain_W(18, 191) <= 0; playAgain_W(18, 192) <= 0; playAgain_W(18, 193) <= 0; playAgain_W(18, 194) <= 0; playAgain_W(18, 195) <= 0; playAgain_W(18, 196) <= 0; playAgain_W(18, 197) <= 0; playAgain_W(18, 198) <= 0; playAgain_W(18, 199) <= 0; playAgain_W(18, 200) <= 0; playAgain_W(18, 201) <= 0; playAgain_W(18, 202) <= 0; playAgain_W(18, 203) <= 0; playAgain_W(18, 204) <= 0; playAgain_W(18, 205) <= 0; playAgain_W(18, 206) <= 0; playAgain_W(18, 207) <= 0; playAgain_W(18, 208) <= 0; playAgain_W(18, 209) <= 0; playAgain_W(18, 210) <= 0; playAgain_W(18, 211) <= 0; playAgain_W(18, 212) <= 0; playAgain_W(18, 213) <= 0; playAgain_W(18, 214) <= 0; playAgain_W(18, 215) <= 0; playAgain_W(18, 216) <= 1; playAgain_W(18, 217) <= 1; playAgain_W(18, 218) <= 1; playAgain_W(18, 219) <= 1; playAgain_W(18, 220) <= 1; playAgain_W(18, 221) <= 1; playAgain_W(18, 222) <= 1; playAgain_W(18, 223) <= 1; playAgain_W(18, 224) <= 1; playAgain_W(18, 225) <= 1; playAgain_W(18, 226) <= 1; playAgain_W(18, 227) <= 1; playAgain_W(18, 228) <= 0; playAgain_W(18, 229) <= 0; playAgain_W(18, 230) <= 0; playAgain_W(18, 231) <= 0; playAgain_W(18, 232) <= 0; playAgain_W(18, 233) <= 0; playAgain_W(18, 234) <= 0; playAgain_W(18, 235) <= 0; playAgain_W(18, 236) <= 0; playAgain_W(18, 237) <= 0; playAgain_W(18, 238) <= 1; playAgain_W(18, 239) <= 1; playAgain_W(18, 240) <= 1; playAgain_W(18, 241) <= 1; playAgain_W(18, 242) <= 1; playAgain_W(18, 243) <= 1; playAgain_W(18, 244) <= 1; playAgain_W(18, 245) <= 1; playAgain_W(18, 246) <= 0; playAgain_W(18, 247) <= 0; playAgain_W(18, 248) <= 0; playAgain_W(18, 249) <= 0; playAgain_W(18, 250) <= 0; playAgain_W(18, 251) <= 0; playAgain_W(18, 252) <= 1; playAgain_W(18, 253) <= 1; playAgain_W(18, 254) <= 1; playAgain_W(18, 255) <= 1; playAgain_W(18, 256) <= 0; playAgain_W(18, 257) <= 0; playAgain_W(18, 258) <= 0; playAgain_W(18, 259) <= 0; playAgain_W(18, 260) <= 0; playAgain_W(18, 261) <= 0; playAgain_W(18, 262) <= 1; playAgain_W(18, 263) <= 1; playAgain_W(18, 264) <= 1; playAgain_W(18, 265) <= 1; playAgain_W(18, 266) <= 0; playAgain_W(18, 267) <= 0; playAgain_W(18, 268) <= 0; playAgain_W(18, 269) <= 0; playAgain_W(18, 270) <= 1; playAgain_W(18, 271) <= 1; playAgain_W(18, 272) <= 1; playAgain_W(18, 273) <= 1; playAgain_W(18, 274) <= 1; playAgain_W(18, 275) <= 1; playAgain_W(18, 276) <= 1; playAgain_W(18, 277) <= 1; playAgain_W(18, 278) <= 1; playAgain_W(18, 279) <= 1; playAgain_W(18, 280) <= 0; playAgain_W(18, 281) <= 0; playAgain_W(18, 282) <= 0; playAgain_W(18, 283) <= 0; playAgain_W(18, 284) <= 0; playAgain_W(18, 285) <= 0; playAgain_W(18, 286) <= 0; playAgain_W(18, 287) <= 0; 
playAgain_W(19, 0) <= 1; playAgain_W(19, 1) <= 1; playAgain_W(19, 2) <= 1; playAgain_W(19, 3) <= 1; playAgain_W(19, 4) <= 1; playAgain_W(19, 5) <= 1; playAgain_W(19, 6) <= 1; playAgain_W(19, 7) <= 1; playAgain_W(19, 8) <= 0; playAgain_W(19, 9) <= 0; playAgain_W(19, 10) <= 0; playAgain_W(19, 11) <= 0; playAgain_W(19, 12) <= 0; playAgain_W(19, 13) <= 0; playAgain_W(19, 14) <= 0; playAgain_W(19, 15) <= 0; playAgain_W(19, 16) <= 0; playAgain_W(19, 17) <= 0; playAgain_W(19, 18) <= 1; playAgain_W(19, 19) <= 1; playAgain_W(19, 20) <= 1; playAgain_W(19, 21) <= 1; playAgain_W(19, 22) <= 1; playAgain_W(19, 23) <= 1; playAgain_W(19, 24) <= 1; playAgain_W(19, 25) <= 1; playAgain_W(19, 26) <= 1; playAgain_W(19, 27) <= 1; playAgain_W(19, 28) <= 1; playAgain_W(19, 29) <= 1; playAgain_W(19, 30) <= 1; playAgain_W(19, 31) <= 1; playAgain_W(19, 32) <= 0; playAgain_W(19, 33) <= 0; playAgain_W(19, 34) <= 0; playAgain_W(19, 35) <= 0; playAgain_W(19, 36) <= 1; playAgain_W(19, 37) <= 1; playAgain_W(19, 38) <= 1; playAgain_W(19, 39) <= 1; playAgain_W(19, 40) <= 0; playAgain_W(19, 41) <= 0; playAgain_W(19, 42) <= 0; playAgain_W(19, 43) <= 0; playAgain_W(19, 44) <= 0; playAgain_W(19, 45) <= 0; playAgain_W(19, 46) <= 1; playAgain_W(19, 47) <= 1; playAgain_W(19, 48) <= 1; playAgain_W(19, 49) <= 1; playAgain_W(19, 50) <= 0; playAgain_W(19, 51) <= 0; playAgain_W(19, 52) <= 0; playAgain_W(19, 53) <= 0; playAgain_W(19, 54) <= 0; playAgain_W(19, 55) <= 0; playAgain_W(19, 56) <= 0; playAgain_W(19, 57) <= 0; playAgain_W(19, 58) <= 1; playAgain_W(19, 59) <= 1; playAgain_W(19, 60) <= 1; playAgain_W(19, 61) <= 1; playAgain_W(19, 62) <= 1; playAgain_W(19, 63) <= 1; playAgain_W(19, 64) <= 1; playAgain_W(19, 65) <= 1; playAgain_W(19, 66) <= 0; playAgain_W(19, 67) <= 0; playAgain_W(19, 68) <= 0; playAgain_W(19, 69) <= 0; playAgain_W(19, 70) <= 0; playAgain_W(19, 71) <= 0; playAgain_W(19, 72) <= 0; playAgain_W(19, 73) <= 0; playAgain_W(19, 74) <= 0; playAgain_W(19, 75) <= 0; playAgain_W(19, 76) <= 0; playAgain_W(19, 77) <= 0; playAgain_W(19, 78) <= 0; playAgain_W(19, 79) <= 0; playAgain_W(19, 80) <= 0; playAgain_W(19, 81) <= 0; playAgain_W(19, 82) <= 0; playAgain_W(19, 83) <= 0; playAgain_W(19, 84) <= 0; playAgain_W(19, 85) <= 0; playAgain_W(19, 86) <= 0; playAgain_W(19, 87) <= 0; playAgain_W(19, 88) <= 0; playAgain_W(19, 89) <= 0; playAgain_W(19, 90) <= 1; playAgain_W(19, 91) <= 1; playAgain_W(19, 92) <= 1; playAgain_W(19, 93) <= 1; playAgain_W(19, 94) <= 0; playAgain_W(19, 95) <= 0; playAgain_W(19, 96) <= 0; playAgain_W(19, 97) <= 0; playAgain_W(19, 98) <= 0; playAgain_W(19, 99) <= 0; playAgain_W(19, 100) <= 1; playAgain_W(19, 101) <= 1; playAgain_W(19, 102) <= 1; playAgain_W(19, 103) <= 1; playAgain_W(19, 104) <= 0; playAgain_W(19, 105) <= 0; playAgain_W(19, 106) <= 0; playAgain_W(19, 107) <= 0; playAgain_W(19, 108) <= 0; playAgain_W(19, 109) <= 0; playAgain_W(19, 110) <= 0; playAgain_W(19, 111) <= 0; playAgain_W(19, 112) <= 1; playAgain_W(19, 113) <= 1; playAgain_W(19, 114) <= 1; playAgain_W(19, 115) <= 1; playAgain_W(19, 116) <= 1; playAgain_W(19, 117) <= 1; playAgain_W(19, 118) <= 0; playAgain_W(19, 119) <= 0; playAgain_W(19, 120) <= 1; playAgain_W(19, 121) <= 1; playAgain_W(19, 122) <= 0; playAgain_W(19, 123) <= 0; playAgain_W(19, 124) <= 0; playAgain_W(19, 125) <= 0; playAgain_W(19, 126) <= 1; playAgain_W(19, 127) <= 1; playAgain_W(19, 128) <= 1; playAgain_W(19, 129) <= 1; playAgain_W(19, 130) <= 0; playAgain_W(19, 131) <= 0; playAgain_W(19, 132) <= 0; playAgain_W(19, 133) <= 0; playAgain_W(19, 134) <= 0; playAgain_W(19, 135) <= 0; playAgain_W(19, 136) <= 1; playAgain_W(19, 137) <= 1; playAgain_W(19, 138) <= 1; playAgain_W(19, 139) <= 1; playAgain_W(19, 140) <= 0; playAgain_W(19, 141) <= 0; playAgain_W(19, 142) <= 0; playAgain_W(19, 143) <= 0; playAgain_W(19, 144) <= 0; playAgain_W(19, 145) <= 0; playAgain_W(19, 146) <= 0; playAgain_W(19, 147) <= 0; playAgain_W(19, 148) <= 1; playAgain_W(19, 149) <= 1; playAgain_W(19, 150) <= 1; playAgain_W(19, 151) <= 1; playAgain_W(19, 152) <= 1; playAgain_W(19, 153) <= 1; playAgain_W(19, 154) <= 1; playAgain_W(19, 155) <= 1; playAgain_W(19, 156) <= 0; playAgain_W(19, 157) <= 0; playAgain_W(19, 158) <= 0; playAgain_W(19, 159) <= 0; playAgain_W(19, 160) <= 0; playAgain_W(19, 161) <= 0; playAgain_W(19, 162) <= 1; playAgain_W(19, 163) <= 1; playAgain_W(19, 164) <= 1; playAgain_W(19, 165) <= 1; playAgain_W(19, 166) <= 0; playAgain_W(19, 167) <= 0; playAgain_W(19, 168) <= 0; playAgain_W(19, 169) <= 0; playAgain_W(19, 170) <= 0; playAgain_W(19, 171) <= 0; playAgain_W(19, 172) <= 1; playAgain_W(19, 173) <= 1; playAgain_W(19, 174) <= 1; playAgain_W(19, 175) <= 1; playAgain_W(19, 176) <= 0; playAgain_W(19, 177) <= 0; playAgain_W(19, 178) <= 0; playAgain_W(19, 179) <= 0; playAgain_W(19, 180) <= 0; playAgain_W(19, 181) <= 0; playAgain_W(19, 182) <= 0; playAgain_W(19, 183) <= 0; playAgain_W(19, 184) <= 0; playAgain_W(19, 185) <= 0; playAgain_W(19, 186) <= 0; playAgain_W(19, 187) <= 0; playAgain_W(19, 188) <= 0; playAgain_W(19, 189) <= 0; playAgain_W(19, 190) <= 0; playAgain_W(19, 191) <= 0; playAgain_W(19, 192) <= 0; playAgain_W(19, 193) <= 0; playAgain_W(19, 194) <= 0; playAgain_W(19, 195) <= 0; playAgain_W(19, 196) <= 0; playAgain_W(19, 197) <= 0; playAgain_W(19, 198) <= 0; playAgain_W(19, 199) <= 0; playAgain_W(19, 200) <= 0; playAgain_W(19, 201) <= 0; playAgain_W(19, 202) <= 0; playAgain_W(19, 203) <= 0; playAgain_W(19, 204) <= 0; playAgain_W(19, 205) <= 0; playAgain_W(19, 206) <= 0; playAgain_W(19, 207) <= 0; playAgain_W(19, 208) <= 0; playAgain_W(19, 209) <= 0; playAgain_W(19, 210) <= 0; playAgain_W(19, 211) <= 0; playAgain_W(19, 212) <= 0; playAgain_W(19, 213) <= 0; playAgain_W(19, 214) <= 0; playAgain_W(19, 215) <= 0; playAgain_W(19, 216) <= 1; playAgain_W(19, 217) <= 1; playAgain_W(19, 218) <= 1; playAgain_W(19, 219) <= 1; playAgain_W(19, 220) <= 1; playAgain_W(19, 221) <= 1; playAgain_W(19, 222) <= 1; playAgain_W(19, 223) <= 1; playAgain_W(19, 224) <= 1; playAgain_W(19, 225) <= 1; playAgain_W(19, 226) <= 1; playAgain_W(19, 227) <= 1; playAgain_W(19, 228) <= 0; playAgain_W(19, 229) <= 0; playAgain_W(19, 230) <= 0; playAgain_W(19, 231) <= 0; playAgain_W(19, 232) <= 0; playAgain_W(19, 233) <= 0; playAgain_W(19, 234) <= 0; playAgain_W(19, 235) <= 0; playAgain_W(19, 236) <= 0; playAgain_W(19, 237) <= 0; playAgain_W(19, 238) <= 1; playAgain_W(19, 239) <= 1; playAgain_W(19, 240) <= 1; playAgain_W(19, 241) <= 1; playAgain_W(19, 242) <= 1; playAgain_W(19, 243) <= 1; playAgain_W(19, 244) <= 1; playAgain_W(19, 245) <= 1; playAgain_W(19, 246) <= 0; playAgain_W(19, 247) <= 0; playAgain_W(19, 248) <= 0; playAgain_W(19, 249) <= 0; playAgain_W(19, 250) <= 0; playAgain_W(19, 251) <= 0; playAgain_W(19, 252) <= 1; playAgain_W(19, 253) <= 1; playAgain_W(19, 254) <= 1; playAgain_W(19, 255) <= 1; playAgain_W(19, 256) <= 0; playAgain_W(19, 257) <= 0; playAgain_W(19, 258) <= 0; playAgain_W(19, 259) <= 0; playAgain_W(19, 260) <= 0; playAgain_W(19, 261) <= 0; playAgain_W(19, 262) <= 1; playAgain_W(19, 263) <= 1; playAgain_W(19, 264) <= 1; playAgain_W(19, 265) <= 1; playAgain_W(19, 266) <= 0; playAgain_W(19, 267) <= 0; playAgain_W(19, 268) <= 0; playAgain_W(19, 269) <= 0; playAgain_W(19, 270) <= 1; playAgain_W(19, 271) <= 1; playAgain_W(19, 272) <= 1; playAgain_W(19, 273) <= 1; playAgain_W(19, 274) <= 1; playAgain_W(19, 275) <= 1; playAgain_W(19, 276) <= 1; playAgain_W(19, 277) <= 1; playAgain_W(19, 278) <= 1; playAgain_W(19, 279) <= 1; playAgain_W(19, 280) <= 0; playAgain_W(19, 281) <= 0; playAgain_W(19, 282) <= 0; playAgain_W(19, 283) <= 0; playAgain_W(19, 284) <= 0; playAgain_W(19, 285) <= 0; playAgain_W(19, 286) <= 0; playAgain_W(19, 287) <= 0; 



end Behavioral;
