
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package endpkg is
    type end2D is array(0 to 39, 0 to 323) of integer;
end package;

use work.endpkg.all;

entity gameover is
    Port (end_W: out end2D);
end gameover;

architecture Behavioral of gameover is

begin

end_W(0, 0) <= 0; end_W(0, 1) <= 0; end_W(0, 2) <= 0; end_W(0, 3) <= 0; end_W(0, 4) <= 0; end_W(0, 5) <= 0; end_W(0, 6) <= 0; end_W(0, 7) <= 0; 
end_W(0, 8) <= 1; end_W(0, 9) <= 1; end_W(0, 10) <= 1; end_W(0, 11) <= 1; end_W(0, 12) <= 1; end_W(0, 13) <= 1; end_W(0, 14) <= 1; end_W(0, 15) <= 1; 
end_W(0, 16) <= 1; end_W(0, 17) <= 1; end_W(0, 18) <= 1; end_W(0, 19) <= 1; end_W(0, 20) <= 1; end_W(0, 21) <= 1; end_W(0, 22) <= 1; end_W(0, 23) <= 1; 
end_W(0, 24) <= 0; end_W(0, 25) <= 0; end_W(0, 26) <= 0; end_W(0, 27) <= 0; end_W(0, 28) <= 0; end_W(0, 29) <= 0; end_W(0, 30) <= 0; end_W(0, 31) <= 0; 
end_W(0, 32) <= 0; end_W(0, 33) <= 0; end_W(0, 34) <= 0; end_W(0, 35) <= 0; end_W(0, 36) <= 0; end_W(0, 37) <= 0; end_W(0, 38) <= 0; end_W(0, 39) <= 0; 
end_W(0, 40) <= 0; end_W(0, 41) <= 0; end_W(0, 42) <= 0; end_W(0, 43) <= 0; end_W(0, 44) <= 0; end_W(0, 45) <= 0; end_W(0, 46) <= 0; end_W(0, 47) <= 0; 
end_W(0, 48) <= 1; end_W(0, 49) <= 1; end_W(0, 50) <= 1; end_W(0, 51) <= 1; end_W(0, 52) <= 0; end_W(0, 53) <= 0; end_W(0, 54) <= 0; end_W(0, 55) <= 0; 
end_W(0, 56) <= 0; end_W(0, 57) <= 0; end_W(0, 58) <= 0; end_W(0, 59) <= 0; end_W(0, 60) <= 0; end_W(0, 61) <= 0; end_W(0, 62) <= 0; end_W(0, 63) <= 0; 
end_W(0, 64) <= 0; end_W(0, 65) <= 0; end_W(0, 66) <= 0; end_W(0, 67) <= 0; end_W(0, 68) <= 0; end_W(0, 69) <= 0; end_W(0, 70) <= 0; end_W(0, 71) <= 0; 
end_W(0, 72) <= 1; end_W(0, 73) <= 1; end_W(0, 74) <= 1; end_W(0, 75) <= 1; end_W(0, 76) <= 1; end_W(0, 77) <= 1; end_W(0, 78) <= 1; end_W(0, 79) <= 1; 
end_W(0, 80) <= 0; end_W(0, 81) <= 0; end_W(0, 82) <= 0; end_W(0, 83) <= 0; end_W(0, 84) <= 0; end_W(0, 85) <= 0; end_W(0, 86) <= 0; end_W(0, 87) <= 0; 
end_W(0, 88) <= 0; end_W(0, 89) <= 0; end_W(0, 90) <= 0; end_W(0, 91) <= 0; end_W(0, 92) <= 0; end_W(0, 93) <= 0; end_W(0, 94) <= 0; end_W(0, 95) <= 0; 
end_W(0, 96) <= 1; end_W(0, 97) <= 1; end_W(0, 98) <= 1; end_W(0, 99) <= 1; end_W(0, 100) <= 1; end_W(0, 101) <= 1; end_W(0, 102) <= 1; end_W(0, 103) <= 1; 
end_W(0, 104) <= 0; end_W(0, 105) <= 0; end_W(0, 106) <= 0; end_W(0, 107) <= 0; end_W(0, 108) <= 1; end_W(0, 109) <= 1; end_W(0, 110) <= 1; end_W(0, 111) <= 1; 
end_W(0, 112) <= 1; end_W(0, 113) <= 1; end_W(0, 114) <= 1; end_W(0, 115) <= 1; end_W(0, 116) <= 1; end_W(0, 117) <= 1; end_W(0, 118) <= 1; end_W(0, 119) <= 1; 
end_W(0, 120) <= 1; end_W(0, 121) <= 1; end_W(0, 122) <= 1; end_W(0, 123) <= 1; end_W(0, 124) <= 1; end_W(0, 125) <= 1; end_W(0, 126) <= 1; end_W(0, 127) <= 1; 
end_W(0, 128) <= 1; end_W(0, 129) <= 1; end_W(0, 130) <= 1; end_W(0, 131) <= 1; end_W(0, 132) <= 1; end_W(0, 133) <= 1; end_W(0, 134) <= 1; end_W(0, 135) <= 1; 
end_W(0, 136) <= 0; end_W(0, 137) <= 0; end_W(0, 138) <= 0; end_W(0, 139) <= 0; end_W(0, 140) <= 0; end_W(0, 141) <= 0; end_W(0, 142) <= 0; end_W(0, 143) <= 0; 
end_W(0, 144) <= 0; end_W(0, 145) <= 0; end_W(0, 146) <= 0; end_W(0, 147) <= 0; end_W(0, 148) <= 0; end_W(0, 149) <= 0; end_W(0, 150) <= 0; end_W(0, 151) <= 0; 
end_W(0, 152) <= 0; end_W(0, 153) <= 0; end_W(0, 154) <= 0; end_W(0, 155) <= 0; end_W(0, 156) <= 0; end_W(0, 157) <= 0; end_W(0, 158) <= 0; end_W(0, 159) <= 0; 
end_W(0, 160) <= 0; end_W(0, 161) <= 0; end_W(0, 162) <= 0; end_W(0, 163) <= 0; end_W(0, 164) <= 0; end_W(0, 165) <= 0; end_W(0, 166) <= 0; end_W(0, 167) <= 0; 
end_W(0, 168) <= 0; end_W(0, 169) <= 0; end_W(0, 170) <= 0; end_W(0, 171) <= 0; end_W(0, 172) <= 0; end_W(0, 173) <= 0; end_W(0, 174) <= 0; end_W(0, 175) <= 0; 
end_W(0, 176) <= 0; end_W(0, 177) <= 0; end_W(0, 178) <= 0; end_W(0, 179) <= 0; end_W(0, 180) <= 0; end_W(0, 181) <= 0; end_W(0, 182) <= 0; end_W(0, 183) <= 0; 
end_W(0, 184) <= 1; end_W(0, 185) <= 1; end_W(0, 186) <= 1; end_W(0, 187) <= 1; end_W(0, 188) <= 1; end_W(0, 189) <= 1; end_W(0, 190) <= 1; end_W(0, 191) <= 1; 
end_W(0, 192) <= 1; end_W(0, 193) <= 1; end_W(0, 194) <= 1; end_W(0, 195) <= 1; end_W(0, 196) <= 1; end_W(0, 197) <= 1; end_W(0, 198) <= 1; end_W(0, 199) <= 1; 
end_W(0, 200) <= 1; end_W(0, 201) <= 1; end_W(0, 202) <= 1; end_W(0, 203) <= 1; end_W(0, 204) <= 0; end_W(0, 205) <= 0; end_W(0, 206) <= 0; end_W(0, 207) <= 0; 
end_W(0, 208) <= 0; end_W(0, 209) <= 0; end_W(0, 210) <= 0; end_W(0, 211) <= 0; end_W(0, 212) <= 0; end_W(0, 213) <= 0; end_W(0, 214) <= 0; end_W(0, 215) <= 0; 
end_W(0, 216) <= 1; end_W(0, 217) <= 1; end_W(0, 218) <= 1; end_W(0, 219) <= 1; end_W(0, 220) <= 1; end_W(0, 221) <= 1; end_W(0, 222) <= 1; end_W(0, 223) <= 1; 
end_W(0, 224) <= 0; end_W(0, 225) <= 0; end_W(0, 226) <= 0; end_W(0, 227) <= 0; end_W(0, 228) <= 0; end_W(0, 229) <= 0; end_W(0, 230) <= 0; end_W(0, 231) <= 0; 
end_W(0, 232) <= 0; end_W(0, 233) <= 0; end_W(0, 234) <= 0; end_W(0, 235) <= 0; end_W(0, 236) <= 0; end_W(0, 237) <= 0; end_W(0, 238) <= 0; end_W(0, 239) <= 0; 
end_W(0, 240) <= 1; end_W(0, 241) <= 1; end_W(0, 242) <= 1; end_W(0, 243) <= 1; end_W(0, 244) <= 1; end_W(0, 245) <= 1; end_W(0, 246) <= 1; end_W(0, 247) <= 1; 
end_W(0, 248) <= 0; end_W(0, 249) <= 0; end_W(0, 250) <= 0; end_W(0, 251) <= 0; end_W(0, 252) <= 1; end_W(0, 253) <= 1; end_W(0, 254) <= 1; end_W(0, 255) <= 1; 
end_W(0, 256) <= 1; end_W(0, 257) <= 1; end_W(0, 258) <= 1; end_W(0, 259) <= 1; end_W(0, 260) <= 1; end_W(0, 261) <= 1; end_W(0, 262) <= 1; end_W(0, 263) <= 1; 
end_W(0, 264) <= 1; end_W(0, 265) <= 1; end_W(0, 266) <= 1; end_W(0, 267) <= 1; end_W(0, 268) <= 1; end_W(0, 269) <= 1; end_W(0, 270) <= 1; end_W(0, 271) <= 1; 
end_W(0, 272) <= 1; end_W(0, 273) <= 1; end_W(0, 274) <= 1; end_W(0, 275) <= 1; end_W(0, 276) <= 1; end_W(0, 277) <= 1; end_W(0, 278) <= 1; end_W(0, 279) <= 1; 
end_W(0, 280) <= 0; end_W(0, 281) <= 0; end_W(0, 282) <= 0; end_W(0, 283) <= 0; end_W(0, 284) <= 0; end_W(0, 285) <= 0; end_W(0, 286) <= 0; end_W(0, 287) <= 0; 
end_W(0, 288) <= 1; end_W(0, 289) <= 1; end_W(0, 290) <= 1; end_W(0, 291) <= 1; end_W(0, 292) <= 1; end_W(0, 293) <= 1; end_W(0, 294) <= 1; end_W(0, 295) <= 1; 
end_W(0, 296) <= 1; end_W(0, 297) <= 1; end_W(0, 298) <= 1; end_W(0, 299) <= 1; end_W(0, 300) <= 1; end_W(0, 301) <= 1; end_W(0, 302) <= 1; end_W(0, 303) <= 1; 
end_W(0, 304) <= 1; end_W(0, 305) <= 1; end_W(0, 306) <= 1; end_W(0, 307) <= 1; end_W(0, 308) <= 1; end_W(0, 309) <= 1; end_W(0, 310) <= 1; end_W(0, 311) <= 1; 
end_W(0, 312) <= 0; end_W(0, 313) <= 0; end_W(0, 314) <= 0; end_W(0, 315) <= 0; end_W(0, 316) <= 0; end_W(0, 317) <= 0; end_W(0, 318) <= 0; end_W(0, 319) <= 0; 
end_W(0, 320) <= 0; end_W(0, 321) <= 0; end_W(0, 322) <= 0; end_W(0, 323) <= 0; end_W(1, 0) <= 0; end_W(1, 1) <= 0; end_W(1, 2) <= 0; end_W(1, 3) <= 0; end_W(1, 4) <= 0; end_W(1, 5) <= 0; end_W(1, 6) <= 0; end_W(1, 7) <= 0; 
end_W(1, 8) <= 1; end_W(1, 9) <= 1; end_W(1, 10) <= 1; end_W(1, 11) <= 1; end_W(1, 12) <= 1; end_W(1, 13) <= 1; end_W(1, 14) <= 1; end_W(1, 15) <= 1; 
end_W(1, 16) <= 1; end_W(1, 17) <= 1; end_W(1, 18) <= 1; end_W(1, 19) <= 1; end_W(1, 20) <= 1; end_W(1, 21) <= 1; end_W(1, 22) <= 1; end_W(1, 23) <= 1; 
end_W(1, 24) <= 0; end_W(1, 25) <= 0; end_W(1, 26) <= 0; end_W(1, 27) <= 0; end_W(1, 28) <= 0; end_W(1, 29) <= 0; end_W(1, 30) <= 0; end_W(1, 31) <= 0; 
end_W(1, 32) <= 0; end_W(1, 33) <= 0; end_W(1, 34) <= 0; end_W(1, 35) <= 0; end_W(1, 36) <= 0; end_W(1, 37) <= 0; end_W(1, 38) <= 0; end_W(1, 39) <= 0; 
end_W(1, 40) <= 0; end_W(1, 41) <= 0; end_W(1, 42) <= 0; end_W(1, 43) <= 0; end_W(1, 44) <= 0; end_W(1, 45) <= 0; end_W(1, 46) <= 0; end_W(1, 47) <= 0; 
end_W(1, 48) <= 1; end_W(1, 49) <= 1; end_W(1, 50) <= 1; end_W(1, 51) <= 1; end_W(1, 52) <= 0; end_W(1, 53) <= 0; end_W(1, 54) <= 0; end_W(1, 55) <= 0; 
end_W(1, 56) <= 0; end_W(1, 57) <= 0; end_W(1, 58) <= 0; end_W(1, 59) <= 0; end_W(1, 60) <= 0; end_W(1, 61) <= 0; end_W(1, 62) <= 0; end_W(1, 63) <= 0; 
end_W(1, 64) <= 0; end_W(1, 65) <= 0; end_W(1, 66) <= 0; end_W(1, 67) <= 0; end_W(1, 68) <= 0; end_W(1, 69) <= 0; end_W(1, 70) <= 0; end_W(1, 71) <= 0; 
end_W(1, 72) <= 1; end_W(1, 73) <= 1; end_W(1, 74) <= 1; end_W(1, 75) <= 1; end_W(1, 76) <= 1; end_W(1, 77) <= 1; end_W(1, 78) <= 1; end_W(1, 79) <= 1; 
end_W(1, 80) <= 0; end_W(1, 81) <= 0; end_W(1, 82) <= 0; end_W(1, 83) <= 0; end_W(1, 84) <= 0; end_W(1, 85) <= 0; end_W(1, 86) <= 0; end_W(1, 87) <= 0; 
end_W(1, 88) <= 0; end_W(1, 89) <= 0; end_W(1, 90) <= 0; end_W(1, 91) <= 0; end_W(1, 92) <= 0; end_W(1, 93) <= 0; end_W(1, 94) <= 0; end_W(1, 95) <= 0; 
end_W(1, 96) <= 1; end_W(1, 97) <= 1; end_W(1, 98) <= 1; end_W(1, 99) <= 1; end_W(1, 100) <= 1; end_W(1, 101) <= 1; end_W(1, 102) <= 1; end_W(1, 103) <= 1; 
end_W(1, 104) <= 0; end_W(1, 105) <= 0; end_W(1, 106) <= 0; end_W(1, 107) <= 0; end_W(1, 108) <= 1; end_W(1, 109) <= 1; end_W(1, 110) <= 1; end_W(1, 111) <= 1; 
end_W(1, 112) <= 1; end_W(1, 113) <= 1; end_W(1, 114) <= 1; end_W(1, 115) <= 1; end_W(1, 116) <= 1; end_W(1, 117) <= 1; end_W(1, 118) <= 1; end_W(1, 119) <= 1; 
end_W(1, 120) <= 1; end_W(1, 121) <= 1; end_W(1, 122) <= 1; end_W(1, 123) <= 1; end_W(1, 124) <= 1; end_W(1, 125) <= 1; end_W(1, 126) <= 1; end_W(1, 127) <= 1; 
end_W(1, 128) <= 1; end_W(1, 129) <= 1; end_W(1, 130) <= 1; end_W(1, 131) <= 1; end_W(1, 132) <= 1; end_W(1, 133) <= 1; end_W(1, 134) <= 1; end_W(1, 135) <= 1; 
end_W(1, 136) <= 0; end_W(1, 137) <= 0; end_W(1, 138) <= 0; end_W(1, 139) <= 0; end_W(1, 140) <= 0; end_W(1, 141) <= 0; end_W(1, 142) <= 0; end_W(1, 143) <= 0; 
end_W(1, 144) <= 0; end_W(1, 145) <= 0; end_W(1, 146) <= 0; end_W(1, 147) <= 0; end_W(1, 148) <= 0; end_W(1, 149) <= 0; end_W(1, 150) <= 0; end_W(1, 151) <= 0; 
end_W(1, 152) <= 0; end_W(1, 153) <= 0; end_W(1, 154) <= 0; end_W(1, 155) <= 0; end_W(1, 156) <= 0; end_W(1, 157) <= 0; end_W(1, 158) <= 0; end_W(1, 159) <= 0; 
end_W(1, 160) <= 0; end_W(1, 161) <= 0; end_W(1, 162) <= 0; end_W(1, 163) <= 0; end_W(1, 164) <= 0; end_W(1, 165) <= 0; end_W(1, 166) <= 0; end_W(1, 167) <= 0; 
end_W(1, 168) <= 0; end_W(1, 169) <= 0; end_W(1, 170) <= 0; end_W(1, 171) <= 0; end_W(1, 172) <= 0; end_W(1, 173) <= 0; end_W(1, 174) <= 0; end_W(1, 175) <= 0; 
end_W(1, 176) <= 0; end_W(1, 177) <= 0; end_W(1, 178) <= 0; end_W(1, 179) <= 0; end_W(1, 180) <= 0; end_W(1, 181) <= 0; end_W(1, 182) <= 0; end_W(1, 183) <= 0; 
end_W(1, 184) <= 1; end_W(1, 185) <= 1; end_W(1, 186) <= 1; end_W(1, 187) <= 1; end_W(1, 188) <= 1; end_W(1, 189) <= 1; end_W(1, 190) <= 1; end_W(1, 191) <= 1; 
end_W(1, 192) <= 1; end_W(1, 193) <= 1; end_W(1, 194) <= 1; end_W(1, 195) <= 1; end_W(1, 196) <= 1; end_W(1, 197) <= 1; end_W(1, 198) <= 1; end_W(1, 199) <= 1; 
end_W(1, 200) <= 1; end_W(1, 201) <= 1; end_W(1, 202) <= 1; end_W(1, 203) <= 1; end_W(1, 204) <= 0; end_W(1, 205) <= 0; end_W(1, 206) <= 0; end_W(1, 207) <= 0; 
end_W(1, 208) <= 0; end_W(1, 209) <= 0; end_W(1, 210) <= 0; end_W(1, 211) <= 0; end_W(1, 212) <= 0; end_W(1, 213) <= 0; end_W(1, 214) <= 0; end_W(1, 215) <= 0; 
end_W(1, 216) <= 1; end_W(1, 217) <= 1; end_W(1, 218) <= 1; end_W(1, 219) <= 1; end_W(1, 220) <= 1; end_W(1, 221) <= 1; end_W(1, 222) <= 1; end_W(1, 223) <= 1; 
end_W(1, 224) <= 0; end_W(1, 225) <= 0; end_W(1, 226) <= 0; end_W(1, 227) <= 0; end_W(1, 228) <= 0; end_W(1, 229) <= 0; end_W(1, 230) <= 0; end_W(1, 231) <= 0; 
end_W(1, 232) <= 0; end_W(1, 233) <= 0; end_W(1, 234) <= 0; end_W(1, 235) <= 0; end_W(1, 236) <= 0; end_W(1, 237) <= 0; end_W(1, 238) <= 0; end_W(1, 239) <= 0; 
end_W(1, 240) <= 1; end_W(1, 241) <= 1; end_W(1, 242) <= 1; end_W(1, 243) <= 1; end_W(1, 244) <= 1; end_W(1, 245) <= 1; end_W(1, 246) <= 1; end_W(1, 247) <= 1; 
end_W(1, 248) <= 0; end_W(1, 249) <= 0; end_W(1, 250) <= 0; end_W(1, 251) <= 0; end_W(1, 252) <= 1; end_W(1, 253) <= 1; end_W(1, 254) <= 1; end_W(1, 255) <= 1; 
end_W(1, 256) <= 1; end_W(1, 257) <= 1; end_W(1, 258) <= 1; end_W(1, 259) <= 1; end_W(1, 260) <= 1; end_W(1, 261) <= 1; end_W(1, 262) <= 1; end_W(1, 263) <= 1; 
end_W(1, 264) <= 1; end_W(1, 265) <= 1; end_W(1, 266) <= 1; end_W(1, 267) <= 1; end_W(1, 268) <= 1; end_W(1, 269) <= 1; end_W(1, 270) <= 1; end_W(1, 271) <= 1; 
end_W(1, 272) <= 1; end_W(1, 273) <= 1; end_W(1, 274) <= 1; end_W(1, 275) <= 1; end_W(1, 276) <= 1; end_W(1, 277) <= 1; end_W(1, 278) <= 1; end_W(1, 279) <= 1; 
end_W(1, 280) <= 0; end_W(1, 281) <= 0; end_W(1, 282) <= 0; end_W(1, 283) <= 0; end_W(1, 284) <= 0; end_W(1, 285) <= 0; end_W(1, 286) <= 0; end_W(1, 287) <= 0; 
end_W(1, 288) <= 1; end_W(1, 289) <= 1; end_W(1, 290) <= 1; end_W(1, 291) <= 1; end_W(1, 292) <= 1; end_W(1, 293) <= 1; end_W(1, 294) <= 1; end_W(1, 295) <= 1; 
end_W(1, 296) <= 1; end_W(1, 297) <= 1; end_W(1, 298) <= 1; end_W(1, 299) <= 1; end_W(1, 300) <= 1; end_W(1, 301) <= 1; end_W(1, 302) <= 1; end_W(1, 303) <= 1; 
end_W(1, 304) <= 1; end_W(1, 305) <= 1; end_W(1, 306) <= 1; end_W(1, 307) <= 1; end_W(1, 308) <= 1; end_W(1, 309) <= 1; end_W(1, 310) <= 1; end_W(1, 311) <= 1; 
end_W(1, 312) <= 0; end_W(1, 313) <= 0; end_W(1, 314) <= 0; end_W(1, 315) <= 0; end_W(1, 316) <= 0; end_W(1, 317) <= 0; end_W(1, 318) <= 0; end_W(1, 319) <= 0; 
end_W(1, 320) <= 0; end_W(1, 321) <= 0; end_W(1, 322) <= 0; end_W(1, 323) <= 0; end_W(2, 0) <= 0; end_W(2, 1) <= 0; end_W(2, 2) <= 0; end_W(2, 3) <= 0; end_W(2, 4) <= 0; end_W(2, 5) <= 0; end_W(2, 6) <= 0; end_W(2, 7) <= 0; 
end_W(2, 8) <= 1; end_W(2, 9) <= 1; end_W(2, 10) <= 1; end_W(2, 11) <= 1; end_W(2, 12) <= 1; end_W(2, 13) <= 1; end_W(2, 14) <= 1; end_W(2, 15) <= 1; 
end_W(2, 16) <= 1; end_W(2, 17) <= 1; end_W(2, 18) <= 1; end_W(2, 19) <= 1; end_W(2, 20) <= 1; end_W(2, 21) <= 1; end_W(2, 22) <= 1; end_W(2, 23) <= 1; 
end_W(2, 24) <= 0; end_W(2, 25) <= 0; end_W(2, 26) <= 0; end_W(2, 27) <= 0; end_W(2, 28) <= 0; end_W(2, 29) <= 0; end_W(2, 30) <= 0; end_W(2, 31) <= 0; 
end_W(2, 32) <= 0; end_W(2, 33) <= 0; end_W(2, 34) <= 0; end_W(2, 35) <= 0; end_W(2, 36) <= 0; end_W(2, 37) <= 0; end_W(2, 38) <= 0; end_W(2, 39) <= 0; 
end_W(2, 40) <= 0; end_W(2, 41) <= 0; end_W(2, 42) <= 0; end_W(2, 43) <= 0; end_W(2, 44) <= 0; end_W(2, 45) <= 0; end_W(2, 46) <= 0; end_W(2, 47) <= 0; 
end_W(2, 48) <= 1; end_W(2, 49) <= 1; end_W(2, 50) <= 1; end_W(2, 51) <= 1; end_W(2, 52) <= 0; end_W(2, 53) <= 0; end_W(2, 54) <= 0; end_W(2, 55) <= 0; 
end_W(2, 56) <= 0; end_W(2, 57) <= 0; end_W(2, 58) <= 0; end_W(2, 59) <= 0; end_W(2, 60) <= 0; end_W(2, 61) <= 0; end_W(2, 62) <= 0; end_W(2, 63) <= 0; 
end_W(2, 64) <= 0; end_W(2, 65) <= 0; end_W(2, 66) <= 0; end_W(2, 67) <= 0; end_W(2, 68) <= 0; end_W(2, 69) <= 0; end_W(2, 70) <= 0; end_W(2, 71) <= 0; 
end_W(2, 72) <= 1; end_W(2, 73) <= 1; end_W(2, 74) <= 1; end_W(2, 75) <= 1; end_W(2, 76) <= 1; end_W(2, 77) <= 1; end_W(2, 78) <= 1; end_W(2, 79) <= 1; 
end_W(2, 80) <= 0; end_W(2, 81) <= 0; end_W(2, 82) <= 0; end_W(2, 83) <= 0; end_W(2, 84) <= 0; end_W(2, 85) <= 0; end_W(2, 86) <= 0; end_W(2, 87) <= 0; 
end_W(2, 88) <= 0; end_W(2, 89) <= 0; end_W(2, 90) <= 0; end_W(2, 91) <= 0; end_W(2, 92) <= 0; end_W(2, 93) <= 0; end_W(2, 94) <= 0; end_W(2, 95) <= 0; 
end_W(2, 96) <= 1; end_W(2, 97) <= 1; end_W(2, 98) <= 1; end_W(2, 99) <= 1; end_W(2, 100) <= 1; end_W(2, 101) <= 1; end_W(2, 102) <= 1; end_W(2, 103) <= 1; 
end_W(2, 104) <= 0; end_W(2, 105) <= 0; end_W(2, 106) <= 0; end_W(2, 107) <= 0; end_W(2, 108) <= 1; end_W(2, 109) <= 1; end_W(2, 110) <= 1; end_W(2, 111) <= 1; 
end_W(2, 112) <= 1; end_W(2, 113) <= 1; end_W(2, 114) <= 1; end_W(2, 115) <= 1; end_W(2, 116) <= 1; end_W(2, 117) <= 1; end_W(2, 118) <= 1; end_W(2, 119) <= 1; 
end_W(2, 120) <= 1; end_W(2, 121) <= 1; end_W(2, 122) <= 1; end_W(2, 123) <= 1; end_W(2, 124) <= 1; end_W(2, 125) <= 1; end_W(2, 126) <= 1; end_W(2, 127) <= 1; 
end_W(2, 128) <= 1; end_W(2, 129) <= 1; end_W(2, 130) <= 1; end_W(2, 131) <= 1; end_W(2, 132) <= 1; end_W(2, 133) <= 1; end_W(2, 134) <= 1; end_W(2, 135) <= 1; 
end_W(2, 136) <= 0; end_W(2, 137) <= 0; end_W(2, 138) <= 0; end_W(2, 139) <= 0; end_W(2, 140) <= 0; end_W(2, 141) <= 0; end_W(2, 142) <= 0; end_W(2, 143) <= 0; 
end_W(2, 144) <= 0; end_W(2, 145) <= 0; end_W(2, 146) <= 0; end_W(2, 147) <= 0; end_W(2, 148) <= 0; end_W(2, 149) <= 0; end_W(2, 150) <= 0; end_W(2, 151) <= 0; 
end_W(2, 152) <= 0; end_W(2, 153) <= 0; end_W(2, 154) <= 0; end_W(2, 155) <= 0; end_W(2, 156) <= 0; end_W(2, 157) <= 0; end_W(2, 158) <= 0; end_W(2, 159) <= 0; 
end_W(2, 160) <= 0; end_W(2, 161) <= 0; end_W(2, 162) <= 0; end_W(2, 163) <= 0; end_W(2, 164) <= 0; end_W(2, 165) <= 0; end_W(2, 166) <= 0; end_W(2, 167) <= 0; 
end_W(2, 168) <= 0; end_W(2, 169) <= 0; end_W(2, 170) <= 0; end_W(2, 171) <= 0; end_W(2, 172) <= 0; end_W(2, 173) <= 0; end_W(2, 174) <= 0; end_W(2, 175) <= 0; 
end_W(2, 176) <= 0; end_W(2, 177) <= 0; end_W(2, 178) <= 0; end_W(2, 179) <= 0; end_W(2, 180) <= 0; end_W(2, 181) <= 0; end_W(2, 182) <= 0; end_W(2, 183) <= 0; 
end_W(2, 184) <= 1; end_W(2, 185) <= 1; end_W(2, 186) <= 1; end_W(2, 187) <= 1; end_W(2, 188) <= 1; end_W(2, 189) <= 1; end_W(2, 190) <= 1; end_W(2, 191) <= 1; 
end_W(2, 192) <= 1; end_W(2, 193) <= 1; end_W(2, 194) <= 1; end_W(2, 195) <= 1; end_W(2, 196) <= 1; end_W(2, 197) <= 1; end_W(2, 198) <= 1; end_W(2, 199) <= 1; 
end_W(2, 200) <= 1; end_W(2, 201) <= 1; end_W(2, 202) <= 1; end_W(2, 203) <= 1; end_W(2, 204) <= 0; end_W(2, 205) <= 0; end_W(2, 206) <= 0; end_W(2, 207) <= 0; 
end_W(2, 208) <= 0; end_W(2, 209) <= 0; end_W(2, 210) <= 0; end_W(2, 211) <= 0; end_W(2, 212) <= 0; end_W(2, 213) <= 0; end_W(2, 214) <= 0; end_W(2, 215) <= 0; 
end_W(2, 216) <= 1; end_W(2, 217) <= 1; end_W(2, 218) <= 1; end_W(2, 219) <= 1; end_W(2, 220) <= 1; end_W(2, 221) <= 1; end_W(2, 222) <= 1; end_W(2, 223) <= 1; 
end_W(2, 224) <= 0; end_W(2, 225) <= 0; end_W(2, 226) <= 0; end_W(2, 227) <= 0; end_W(2, 228) <= 0; end_W(2, 229) <= 0; end_W(2, 230) <= 0; end_W(2, 231) <= 0; 
end_W(2, 232) <= 0; end_W(2, 233) <= 0; end_W(2, 234) <= 0; end_W(2, 235) <= 0; end_W(2, 236) <= 0; end_W(2, 237) <= 0; end_W(2, 238) <= 0; end_W(2, 239) <= 0; 
end_W(2, 240) <= 1; end_W(2, 241) <= 1; end_W(2, 242) <= 1; end_W(2, 243) <= 1; end_W(2, 244) <= 1; end_W(2, 245) <= 1; end_W(2, 246) <= 1; end_W(2, 247) <= 1; 
end_W(2, 248) <= 0; end_W(2, 249) <= 0; end_W(2, 250) <= 0; end_W(2, 251) <= 0; end_W(2, 252) <= 1; end_W(2, 253) <= 1; end_W(2, 254) <= 1; end_W(2, 255) <= 1; 
end_W(2, 256) <= 1; end_W(2, 257) <= 1; end_W(2, 258) <= 1; end_W(2, 259) <= 1; end_W(2, 260) <= 1; end_W(2, 261) <= 1; end_W(2, 262) <= 1; end_W(2, 263) <= 1; 
end_W(2, 264) <= 1; end_W(2, 265) <= 1; end_W(2, 266) <= 1; end_W(2, 267) <= 1; end_W(2, 268) <= 1; end_W(2, 269) <= 1; end_W(2, 270) <= 1; end_W(2, 271) <= 1; 
end_W(2, 272) <= 1; end_W(2, 273) <= 1; end_W(2, 274) <= 1; end_W(2, 275) <= 1; end_W(2, 276) <= 1; end_W(2, 277) <= 1; end_W(2, 278) <= 1; end_W(2, 279) <= 1; 
end_W(2, 280) <= 0; end_W(2, 281) <= 0; end_W(2, 282) <= 0; end_W(2, 283) <= 0; end_W(2, 284) <= 0; end_W(2, 285) <= 0; end_W(2, 286) <= 0; end_W(2, 287) <= 0; 
end_W(2, 288) <= 1; end_W(2, 289) <= 1; end_W(2, 290) <= 1; end_W(2, 291) <= 1; end_W(2, 292) <= 1; end_W(2, 293) <= 1; end_W(2, 294) <= 1; end_W(2, 295) <= 1; 
end_W(2, 296) <= 1; end_W(2, 297) <= 1; end_W(2, 298) <= 1; end_W(2, 299) <= 1; end_W(2, 300) <= 1; end_W(2, 301) <= 1; end_W(2, 302) <= 1; end_W(2, 303) <= 1; 
end_W(2, 304) <= 1; end_W(2, 305) <= 1; end_W(2, 306) <= 1; end_W(2, 307) <= 1; end_W(2, 308) <= 1; end_W(2, 309) <= 1; end_W(2, 310) <= 1; end_W(2, 311) <= 1; 
end_W(2, 312) <= 0; end_W(2, 313) <= 0; end_W(2, 314) <= 0; end_W(2, 315) <= 0; end_W(2, 316) <= 0; end_W(2, 317) <= 0; end_W(2, 318) <= 0; end_W(2, 319) <= 0; 
end_W(2, 320) <= 0; end_W(2, 321) <= 0; end_W(2, 322) <= 0; end_W(2, 323) <= 0; end_W(3, 0) <= 0; end_W(3, 1) <= 0; end_W(3, 2) <= 0; end_W(3, 3) <= 0; end_W(3, 4) <= 0; end_W(3, 5) <= 0; end_W(3, 6) <= 0; end_W(3, 7) <= 0; 
end_W(3, 8) <= 1; end_W(3, 9) <= 1; end_W(3, 10) <= 1; end_W(3, 11) <= 1; end_W(3, 12) <= 1; end_W(3, 13) <= 1; end_W(3, 14) <= 1; end_W(3, 15) <= 1; 
end_W(3, 16) <= 1; end_W(3, 17) <= 1; end_W(3, 18) <= 1; end_W(3, 19) <= 1; end_W(3, 20) <= 1; end_W(3, 21) <= 1; end_W(3, 22) <= 1; end_W(3, 23) <= 1; 
end_W(3, 24) <= 0; end_W(3, 25) <= 0; end_W(3, 26) <= 0; end_W(3, 27) <= 0; end_W(3, 28) <= 0; end_W(3, 29) <= 0; end_W(3, 30) <= 0; end_W(3, 31) <= 0; 
end_W(3, 32) <= 0; end_W(3, 33) <= 0; end_W(3, 34) <= 0; end_W(3, 35) <= 0; end_W(3, 36) <= 0; end_W(3, 37) <= 0; end_W(3, 38) <= 0; end_W(3, 39) <= 0; 
end_W(3, 40) <= 0; end_W(3, 41) <= 0; end_W(3, 42) <= 0; end_W(3, 43) <= 0; end_W(3, 44) <= 0; end_W(3, 45) <= 0; end_W(3, 46) <= 0; end_W(3, 47) <= 0; 
end_W(3, 48) <= 1; end_W(3, 49) <= 1; end_W(3, 50) <= 1; end_W(3, 51) <= 1; end_W(3, 52) <= 0; end_W(3, 53) <= 0; end_W(3, 54) <= 0; end_W(3, 55) <= 0; 
end_W(3, 56) <= 0; end_W(3, 57) <= 0; end_W(3, 58) <= 0; end_W(3, 59) <= 0; end_W(3, 60) <= 0; end_W(3, 61) <= 0; end_W(3, 62) <= 0; end_W(3, 63) <= 0; 
end_W(3, 64) <= 0; end_W(3, 65) <= 0; end_W(3, 66) <= 0; end_W(3, 67) <= 0; end_W(3, 68) <= 0; end_W(3, 69) <= 0; end_W(3, 70) <= 0; end_W(3, 71) <= 0; 
end_W(3, 72) <= 1; end_W(3, 73) <= 1; end_W(3, 74) <= 1; end_W(3, 75) <= 1; end_W(3, 76) <= 1; end_W(3, 77) <= 1; end_W(3, 78) <= 1; end_W(3, 79) <= 1; 
end_W(3, 80) <= 0; end_W(3, 81) <= 0; end_W(3, 82) <= 0; end_W(3, 83) <= 0; end_W(3, 84) <= 0; end_W(3, 85) <= 0; end_W(3, 86) <= 0; end_W(3, 87) <= 0; 
end_W(3, 88) <= 0; end_W(3, 89) <= 0; end_W(3, 90) <= 0; end_W(3, 91) <= 0; end_W(3, 92) <= 0; end_W(3, 93) <= 0; end_W(3, 94) <= 0; end_W(3, 95) <= 0; 
end_W(3, 96) <= 1; end_W(3, 97) <= 1; end_W(3, 98) <= 1; end_W(3, 99) <= 1; end_W(3, 100) <= 1; end_W(3, 101) <= 1; end_W(3, 102) <= 1; end_W(3, 103) <= 1; 
end_W(3, 104) <= 0; end_W(3, 105) <= 0; end_W(3, 106) <= 0; end_W(3, 107) <= 0; end_W(3, 108) <= 1; end_W(3, 109) <= 1; end_W(3, 110) <= 1; end_W(3, 111) <= 1; 
end_W(3, 112) <= 1; end_W(3, 113) <= 1; end_W(3, 114) <= 1; end_W(3, 115) <= 1; end_W(3, 116) <= 1; end_W(3, 117) <= 1; end_W(3, 118) <= 1; end_W(3, 119) <= 1; 
end_W(3, 120) <= 1; end_W(3, 121) <= 1; end_W(3, 122) <= 1; end_W(3, 123) <= 1; end_W(3, 124) <= 1; end_W(3, 125) <= 1; end_W(3, 126) <= 1; end_W(3, 127) <= 1; 
end_W(3, 128) <= 1; end_W(3, 129) <= 1; end_W(3, 130) <= 1; end_W(3, 131) <= 1; end_W(3, 132) <= 1; end_W(3, 133) <= 1; end_W(3, 134) <= 1; end_W(3, 135) <= 1; 
end_W(3, 136) <= 0; end_W(3, 137) <= 0; end_W(3, 138) <= 0; end_W(3, 139) <= 0; end_W(3, 140) <= 0; end_W(3, 141) <= 0; end_W(3, 142) <= 0; end_W(3, 143) <= 0; 
end_W(3, 144) <= 0; end_W(3, 145) <= 0; end_W(3, 146) <= 0; end_W(3, 147) <= 0; end_W(3, 148) <= 0; end_W(3, 149) <= 0; end_W(3, 150) <= 0; end_W(3, 151) <= 0; 
end_W(3, 152) <= 0; end_W(3, 153) <= 0; end_W(3, 154) <= 0; end_W(3, 155) <= 0; end_W(3, 156) <= 0; end_W(3, 157) <= 0; end_W(3, 158) <= 0; end_W(3, 159) <= 0; 
end_W(3, 160) <= 0; end_W(3, 161) <= 0; end_W(3, 162) <= 0; end_W(3, 163) <= 0; end_W(3, 164) <= 0; end_W(3, 165) <= 0; end_W(3, 166) <= 0; end_W(3, 167) <= 0; 
end_W(3, 168) <= 0; end_W(3, 169) <= 0; end_W(3, 170) <= 0; end_W(3, 171) <= 0; end_W(3, 172) <= 0; end_W(3, 173) <= 0; end_W(3, 174) <= 0; end_W(3, 175) <= 0; 
end_W(3, 176) <= 0; end_W(3, 177) <= 0; end_W(3, 178) <= 0; end_W(3, 179) <= 0; end_W(3, 180) <= 0; end_W(3, 181) <= 0; end_W(3, 182) <= 0; end_W(3, 183) <= 0; 
end_W(3, 184) <= 1; end_W(3, 185) <= 1; end_W(3, 186) <= 1; end_W(3, 187) <= 1; end_W(3, 188) <= 1; end_W(3, 189) <= 1; end_W(3, 190) <= 1; end_W(3, 191) <= 1; 
end_W(3, 192) <= 1; end_W(3, 193) <= 1; end_W(3, 194) <= 1; end_W(3, 195) <= 1; end_W(3, 196) <= 1; end_W(3, 197) <= 1; end_W(3, 198) <= 1; end_W(3, 199) <= 1; 
end_W(3, 200) <= 1; end_W(3, 201) <= 1; end_W(3, 202) <= 1; end_W(3, 203) <= 1; end_W(3, 204) <= 0; end_W(3, 205) <= 0; end_W(3, 206) <= 0; end_W(3, 207) <= 0; 
end_W(3, 208) <= 0; end_W(3, 209) <= 0; end_W(3, 210) <= 0; end_W(3, 211) <= 0; end_W(3, 212) <= 0; end_W(3, 213) <= 0; end_W(3, 214) <= 0; end_W(3, 215) <= 0; 
end_W(3, 216) <= 1; end_W(3, 217) <= 1; end_W(3, 218) <= 1; end_W(3, 219) <= 1; end_W(3, 220) <= 1; end_W(3, 221) <= 1; end_W(3, 222) <= 1; end_W(3, 223) <= 1; 
end_W(3, 224) <= 0; end_W(3, 225) <= 0; end_W(3, 226) <= 0; end_W(3, 227) <= 0; end_W(3, 228) <= 0; end_W(3, 229) <= 0; end_W(3, 230) <= 0; end_W(3, 231) <= 0; 
end_W(3, 232) <= 0; end_W(3, 233) <= 0; end_W(3, 234) <= 0; end_W(3, 235) <= 0; end_W(3, 236) <= 0; end_W(3, 237) <= 0; end_W(3, 238) <= 0; end_W(3, 239) <= 0; 
end_W(3, 240) <= 1; end_W(3, 241) <= 1; end_W(3, 242) <= 1; end_W(3, 243) <= 1; end_W(3, 244) <= 1; end_W(3, 245) <= 1; end_W(3, 246) <= 1; end_W(3, 247) <= 1; 
end_W(3, 248) <= 0; end_W(3, 249) <= 0; end_W(3, 250) <= 0; end_W(3, 251) <= 0; end_W(3, 252) <= 1; end_W(3, 253) <= 1; end_W(3, 254) <= 1; end_W(3, 255) <= 1; 
end_W(3, 256) <= 1; end_W(3, 257) <= 1; end_W(3, 258) <= 1; end_W(3, 259) <= 1; end_W(3, 260) <= 1; end_W(3, 261) <= 1; end_W(3, 262) <= 1; end_W(3, 263) <= 1; 
end_W(3, 264) <= 1; end_W(3, 265) <= 1; end_W(3, 266) <= 1; end_W(3, 267) <= 1; end_W(3, 268) <= 1; end_W(3, 269) <= 1; end_W(3, 270) <= 1; end_W(3, 271) <= 1; 
end_W(3, 272) <= 1; end_W(3, 273) <= 1; end_W(3, 274) <= 1; end_W(3, 275) <= 1; end_W(3, 276) <= 1; end_W(3, 277) <= 1; end_W(3, 278) <= 1; end_W(3, 279) <= 1; 
end_W(3, 280) <= 0; end_W(3, 281) <= 0; end_W(3, 282) <= 0; end_W(3, 283) <= 0; end_W(3, 284) <= 0; end_W(3, 285) <= 0; end_W(3, 286) <= 0; end_W(3, 287) <= 0; 
end_W(3, 288) <= 1; end_W(3, 289) <= 1; end_W(3, 290) <= 1; end_W(3, 291) <= 1; end_W(3, 292) <= 1; end_W(3, 293) <= 1; end_W(3, 294) <= 1; end_W(3, 295) <= 1; 
end_W(3, 296) <= 1; end_W(3, 297) <= 1; end_W(3, 298) <= 1; end_W(3, 299) <= 1; end_W(3, 300) <= 1; end_W(3, 301) <= 1; end_W(3, 302) <= 1; end_W(3, 303) <= 1; 
end_W(3, 304) <= 1; end_W(3, 305) <= 1; end_W(3, 306) <= 1; end_W(3, 307) <= 1; end_W(3, 308) <= 1; end_W(3, 309) <= 1; end_W(3, 310) <= 1; end_W(3, 311) <= 1; 
end_W(3, 312) <= 0; end_W(3, 313) <= 0; end_W(3, 314) <= 0; end_W(3, 315) <= 0; end_W(3, 316) <= 0; end_W(3, 317) <= 0; end_W(3, 318) <= 0; end_W(3, 319) <= 0; 
end_W(3, 320) <= 0; end_W(3, 321) <= 0; end_W(3, 322) <= 0; end_W(3, 323) <= 0; end_W(4, 0) <= 0; end_W(4, 1) <= 0; end_W(4, 2) <= 0; end_W(4, 3) <= 0; end_W(4, 4) <= 1; end_W(4, 5) <= 1; end_W(4, 6) <= 1; end_W(4, 7) <= 1; 
end_W(4, 8) <= 1; end_W(4, 9) <= 1; end_W(4, 10) <= 1; end_W(4, 11) <= 1; end_W(4, 12) <= 0; end_W(4, 13) <= 0; end_W(4, 14) <= 0; end_W(4, 15) <= 0; 
end_W(4, 16) <= 0; end_W(4, 17) <= 0; end_W(4, 18) <= 0; end_W(4, 19) <= 0; end_W(4, 20) <= 1; end_W(4, 21) <= 1; end_W(4, 22) <= 1; end_W(4, 23) <= 1; 
end_W(4, 24) <= 1; end_W(4, 25) <= 1; end_W(4, 26) <= 1; end_W(4, 27) <= 1; end_W(4, 28) <= 0; end_W(4, 29) <= 0; end_W(4, 30) <= 0; end_W(4, 31) <= 0; 
end_W(4, 32) <= 0; end_W(4, 33) <= 0; end_W(4, 34) <= 0; end_W(4, 35) <= 0; end_W(4, 36) <= 0; end_W(4, 37) <= 0; end_W(4, 38) <= 0; end_W(4, 39) <= 0; 
end_W(4, 40) <= 0; end_W(4, 41) <= 0; end_W(4, 42) <= 0; end_W(4, 43) <= 0; end_W(4, 44) <= 1; end_W(4, 45) <= 1; end_W(4, 46) <= 1; end_W(4, 47) <= 1; 
end_W(4, 48) <= 1; end_W(4, 49) <= 1; end_W(4, 50) <= 1; end_W(4, 51) <= 1; end_W(4, 52) <= 1; end_W(4, 53) <= 1; end_W(4, 54) <= 1; end_W(4, 55) <= 1; 
end_W(4, 56) <= 0; end_W(4, 57) <= 0; end_W(4, 58) <= 0; end_W(4, 59) <= 0; end_W(4, 60) <= 0; end_W(4, 61) <= 0; end_W(4, 62) <= 0; end_W(4, 63) <= 0; 
end_W(4, 64) <= 0; end_W(4, 65) <= 0; end_W(4, 66) <= 0; end_W(4, 67) <= 0; end_W(4, 68) <= 0; end_W(4, 69) <= 0; end_W(4, 70) <= 0; end_W(4, 71) <= 0; 
end_W(4, 72) <= 1; end_W(4, 73) <= 1; end_W(4, 74) <= 1; end_W(4, 75) <= 1; end_W(4, 76) <= 1; end_W(4, 77) <= 1; end_W(4, 78) <= 1; end_W(4, 79) <= 1; 
end_W(4, 80) <= 1; end_W(4, 81) <= 1; end_W(4, 82) <= 1; end_W(4, 83) <= 1; end_W(4, 84) <= 0; end_W(4, 85) <= 0; end_W(4, 86) <= 0; end_W(4, 87) <= 0; 
end_W(4, 88) <= 0; end_W(4, 89) <= 0; end_W(4, 90) <= 0; end_W(4, 91) <= 0; end_W(4, 92) <= 1; end_W(4, 93) <= 1; end_W(4, 94) <= 1; end_W(4, 95) <= 1; 
end_W(4, 96) <= 1; end_W(4, 97) <= 1; end_W(4, 98) <= 1; end_W(4, 99) <= 1; end_W(4, 100) <= 1; end_W(4, 101) <= 1; end_W(4, 102) <= 1; end_W(4, 103) <= 1; 
end_W(4, 104) <= 0; end_W(4, 105) <= 0; end_W(4, 106) <= 0; end_W(4, 107) <= 0; end_W(4, 108) <= 0; end_W(4, 109) <= 0; end_W(4, 110) <= 0; end_W(4, 111) <= 0; 
end_W(4, 112) <= 1; end_W(4, 113) <= 1; end_W(4, 114) <= 1; end_W(4, 115) <= 1; end_W(4, 116) <= 1; end_W(4, 117) <= 1; end_W(4, 118) <= 1; end_W(4, 119) <= 1; 
end_W(4, 120) <= 0; end_W(4, 121) <= 0; end_W(4, 122) <= 0; end_W(4, 123) <= 0; end_W(4, 124) <= 0; end_W(4, 125) <= 0; end_W(4, 126) <= 0; end_W(4, 127) <= 0; 
end_W(4, 128) <= 1; end_W(4, 129) <= 1; end_W(4, 130) <= 1; end_W(4, 131) <= 1; end_W(4, 132) <= 1; end_W(4, 133) <= 1; end_W(4, 134) <= 1; end_W(4, 135) <= 1; 
end_W(4, 136) <= 0; end_W(4, 137) <= 0; end_W(4, 138) <= 0; end_W(4, 139) <= 0; end_W(4, 140) <= 0; end_W(4, 141) <= 0; end_W(4, 142) <= 0; end_W(4, 143) <= 0; 
end_W(4, 144) <= 0; end_W(4, 145) <= 0; end_W(4, 146) <= 0; end_W(4, 147) <= 0; end_W(4, 148) <= 0; end_W(4, 149) <= 0; end_W(4, 150) <= 0; end_W(4, 151) <= 0; 
end_W(4, 152) <= 0; end_W(4, 153) <= 0; end_W(4, 154) <= 0; end_W(4, 155) <= 0; end_W(4, 156) <= 0; end_W(4, 157) <= 0; end_W(4, 158) <= 0; end_W(4, 159) <= 0; 
end_W(4, 160) <= 0; end_W(4, 161) <= 0; end_W(4, 162) <= 0; end_W(4, 163) <= 0; end_W(4, 164) <= 0; end_W(4, 165) <= 0; end_W(4, 166) <= 0; end_W(4, 167) <= 0; 
end_W(4, 168) <= 0; end_W(4, 169) <= 0; end_W(4, 170) <= 0; end_W(4, 171) <= 0; end_W(4, 172) <= 0; end_W(4, 173) <= 0; end_W(4, 174) <= 0; end_W(4, 175) <= 0; 
end_W(4, 176) <= 0; end_W(4, 177) <= 0; end_W(4, 178) <= 0; end_W(4, 179) <= 0; end_W(4, 180) <= 1; end_W(4, 181) <= 1; end_W(4, 182) <= 1; end_W(4, 183) <= 1; 
end_W(4, 184) <= 1; end_W(4, 185) <= 1; end_W(4, 186) <= 1; end_W(4, 187) <= 1; end_W(4, 188) <= 0; end_W(4, 189) <= 0; end_W(4, 190) <= 0; end_W(4, 191) <= 0; 
end_W(4, 192) <= 0; end_W(4, 193) <= 0; end_W(4, 194) <= 0; end_W(4, 195) <= 0; end_W(4, 196) <= 0; end_W(4, 197) <= 0; end_W(4, 198) <= 0; end_W(4, 199) <= 0; 
end_W(4, 200) <= 1; end_W(4, 201) <= 1; end_W(4, 202) <= 1; end_W(4, 203) <= 1; end_W(4, 204) <= 1; end_W(4, 205) <= 1; end_W(4, 206) <= 1; end_W(4, 207) <= 1; 
end_W(4, 208) <= 0; end_W(4, 209) <= 0; end_W(4, 210) <= 0; end_W(4, 211) <= 0; end_W(4, 212) <= 0; end_W(4, 213) <= 0; end_W(4, 214) <= 0; end_W(4, 215) <= 0; 
end_W(4, 216) <= 1; end_W(4, 217) <= 1; end_W(4, 218) <= 1; end_W(4, 219) <= 1; end_W(4, 220) <= 1; end_W(4, 221) <= 1; end_W(4, 222) <= 1; end_W(4, 223) <= 1; 
end_W(4, 224) <= 0; end_W(4, 225) <= 0; end_W(4, 226) <= 0; end_W(4, 227) <= 0; end_W(4, 228) <= 0; end_W(4, 229) <= 0; end_W(4, 230) <= 0; end_W(4, 231) <= 0; 
end_W(4, 232) <= 0; end_W(4, 233) <= 0; end_W(4, 234) <= 0; end_W(4, 235) <= 0; end_W(4, 236) <= 0; end_W(4, 237) <= 0; end_W(4, 238) <= 0; end_W(4, 239) <= 0; 
end_W(4, 240) <= 1; end_W(4, 241) <= 1; end_W(4, 242) <= 1; end_W(4, 243) <= 1; end_W(4, 244) <= 1; end_W(4, 245) <= 1; end_W(4, 246) <= 1; end_W(4, 247) <= 1; 
end_W(4, 248) <= 0; end_W(4, 249) <= 0; end_W(4, 250) <= 0; end_W(4, 251) <= 0; end_W(4, 252) <= 0; end_W(4, 253) <= 0; end_W(4, 254) <= 0; end_W(4, 255) <= 0; 
end_W(4, 256) <= 1; end_W(4, 257) <= 1; end_W(4, 258) <= 1; end_W(4, 259) <= 1; end_W(4, 260) <= 1; end_W(4, 261) <= 1; end_W(4, 262) <= 1; end_W(4, 263) <= 1; 
end_W(4, 264) <= 0; end_W(4, 265) <= 0; end_W(4, 266) <= 0; end_W(4, 267) <= 0; end_W(4, 268) <= 0; end_W(4, 269) <= 0; end_W(4, 270) <= 0; end_W(4, 271) <= 0; 
end_W(4, 272) <= 1; end_W(4, 273) <= 1; end_W(4, 274) <= 1; end_W(4, 275) <= 1; end_W(4, 276) <= 1; end_W(4, 277) <= 1; end_W(4, 278) <= 1; end_W(4, 279) <= 1; 
end_W(4, 280) <= 0; end_W(4, 281) <= 0; end_W(4, 282) <= 0; end_W(4, 283) <= 0; end_W(4, 284) <= 0; end_W(4, 285) <= 0; end_W(4, 286) <= 0; end_W(4, 287) <= 0; 
end_W(4, 288) <= 0; end_W(4, 289) <= 0; end_W(4, 290) <= 0; end_W(4, 291) <= 0; end_W(4, 292) <= 1; end_W(4, 293) <= 1; end_W(4, 294) <= 1; end_W(4, 295) <= 1; 
end_W(4, 296) <= 1; end_W(4, 297) <= 1; end_W(4, 298) <= 1; end_W(4, 299) <= 1; end_W(4, 300) <= 0; end_W(4, 301) <= 0; end_W(4, 302) <= 0; end_W(4, 303) <= 0; 
end_W(4, 304) <= 0; end_W(4, 305) <= 0; end_W(4, 306) <= 0; end_W(4, 307) <= 0; end_W(4, 308) <= 1; end_W(4, 309) <= 1; end_W(4, 310) <= 1; end_W(4, 311) <= 1; 
end_W(4, 312) <= 1; end_W(4, 313) <= 1; end_W(4, 314) <= 1; end_W(4, 315) <= 1; end_W(4, 316) <= 0; end_W(4, 317) <= 0; end_W(4, 318) <= 0; end_W(4, 319) <= 0; 
end_W(4, 320) <= 0; end_W(4, 321) <= 0; end_W(4, 322) <= 0; end_W(4, 323) <= 0; end_W(5, 0) <= 0; end_W(5, 1) <= 0; end_W(5, 2) <= 0; end_W(5, 3) <= 0; end_W(5, 4) <= 1; end_W(5, 5) <= 1; end_W(5, 6) <= 1; end_W(5, 7) <= 1; 
end_W(5, 8) <= 1; end_W(5, 9) <= 1; end_W(5, 10) <= 1; end_W(5, 11) <= 1; end_W(5, 12) <= 0; end_W(5, 13) <= 0; end_W(5, 14) <= 0; end_W(5, 15) <= 0; 
end_W(5, 16) <= 0; end_W(5, 17) <= 0; end_W(5, 18) <= 0; end_W(5, 19) <= 0; end_W(5, 20) <= 1; end_W(5, 21) <= 1; end_W(5, 22) <= 1; end_W(5, 23) <= 1; 
end_W(5, 24) <= 1; end_W(5, 25) <= 1; end_W(5, 26) <= 1; end_W(5, 27) <= 1; end_W(5, 28) <= 0; end_W(5, 29) <= 0; end_W(5, 30) <= 0; end_W(5, 31) <= 0; 
end_W(5, 32) <= 0; end_W(5, 33) <= 0; end_W(5, 34) <= 0; end_W(5, 35) <= 0; end_W(5, 36) <= 0; end_W(5, 37) <= 0; end_W(5, 38) <= 0; end_W(5, 39) <= 0; 
end_W(5, 40) <= 0; end_W(5, 41) <= 0; end_W(5, 42) <= 0; end_W(5, 43) <= 0; end_W(5, 44) <= 1; end_W(5, 45) <= 1; end_W(5, 46) <= 1; end_W(5, 47) <= 1; 
end_W(5, 48) <= 1; end_W(5, 49) <= 1; end_W(5, 50) <= 1; end_W(5, 51) <= 1; end_W(5, 52) <= 1; end_W(5, 53) <= 1; end_W(5, 54) <= 1; end_W(5, 55) <= 1; 
end_W(5, 56) <= 0; end_W(5, 57) <= 0; end_W(5, 58) <= 0; end_W(5, 59) <= 0; end_W(5, 60) <= 0; end_W(5, 61) <= 0; end_W(5, 62) <= 0; end_W(5, 63) <= 0; 
end_W(5, 64) <= 0; end_W(5, 65) <= 0; end_W(5, 66) <= 0; end_W(5, 67) <= 0; end_W(5, 68) <= 0; end_W(5, 69) <= 0; end_W(5, 70) <= 0; end_W(5, 71) <= 0; 
end_W(5, 72) <= 1; end_W(5, 73) <= 1; end_W(5, 74) <= 1; end_W(5, 75) <= 1; end_W(5, 76) <= 1; end_W(5, 77) <= 1; end_W(5, 78) <= 1; end_W(5, 79) <= 1; 
end_W(5, 80) <= 1; end_W(5, 81) <= 1; end_W(5, 82) <= 1; end_W(5, 83) <= 1; end_W(5, 84) <= 0; end_W(5, 85) <= 0; end_W(5, 86) <= 0; end_W(5, 87) <= 0; 
end_W(5, 88) <= 0; end_W(5, 89) <= 0; end_W(5, 90) <= 0; end_W(5, 91) <= 0; end_W(5, 92) <= 1; end_W(5, 93) <= 1; end_W(5, 94) <= 1; end_W(5, 95) <= 1; 
end_W(5, 96) <= 1; end_W(5, 97) <= 1; end_W(5, 98) <= 1; end_W(5, 99) <= 1; end_W(5, 100) <= 1; end_W(5, 101) <= 1; end_W(5, 102) <= 1; end_W(5, 103) <= 1; 
end_W(5, 104) <= 0; end_W(5, 105) <= 0; end_W(5, 106) <= 0; end_W(5, 107) <= 0; end_W(5, 108) <= 0; end_W(5, 109) <= 0; end_W(5, 110) <= 0; end_W(5, 111) <= 0; 
end_W(5, 112) <= 1; end_W(5, 113) <= 1; end_W(5, 114) <= 1; end_W(5, 115) <= 1; end_W(5, 116) <= 1; end_W(5, 117) <= 1; end_W(5, 118) <= 1; end_W(5, 119) <= 1; 
end_W(5, 120) <= 0; end_W(5, 121) <= 0; end_W(5, 122) <= 0; end_W(5, 123) <= 0; end_W(5, 124) <= 0; end_W(5, 125) <= 0; end_W(5, 126) <= 0; end_W(5, 127) <= 0; 
end_W(5, 128) <= 1; end_W(5, 129) <= 1; end_W(5, 130) <= 1; end_W(5, 131) <= 1; end_W(5, 132) <= 1; end_W(5, 133) <= 1; end_W(5, 134) <= 1; end_W(5, 135) <= 1; 
end_W(5, 136) <= 0; end_W(5, 137) <= 0; end_W(5, 138) <= 0; end_W(5, 139) <= 0; end_W(5, 140) <= 0; end_W(5, 141) <= 0; end_W(5, 142) <= 0; end_W(5, 143) <= 0; 
end_W(5, 144) <= 0; end_W(5, 145) <= 0; end_W(5, 146) <= 0; end_W(5, 147) <= 0; end_W(5, 148) <= 0; end_W(5, 149) <= 0; end_W(5, 150) <= 0; end_W(5, 151) <= 0; 
end_W(5, 152) <= 0; end_W(5, 153) <= 0; end_W(5, 154) <= 0; end_W(5, 155) <= 0; end_W(5, 156) <= 0; end_W(5, 157) <= 0; end_W(5, 158) <= 0; end_W(5, 159) <= 0; 
end_W(5, 160) <= 0; end_W(5, 161) <= 0; end_W(5, 162) <= 0; end_W(5, 163) <= 0; end_W(5, 164) <= 0; end_W(5, 165) <= 0; end_W(5, 166) <= 0; end_W(5, 167) <= 0; 
end_W(5, 168) <= 0; end_W(5, 169) <= 0; end_W(5, 170) <= 0; end_W(5, 171) <= 0; end_W(5, 172) <= 0; end_W(5, 173) <= 0; end_W(5, 174) <= 0; end_W(5, 175) <= 0; 
end_W(5, 176) <= 0; end_W(5, 177) <= 0; end_W(5, 178) <= 0; end_W(5, 179) <= 0; end_W(5, 180) <= 1; end_W(5, 181) <= 1; end_W(5, 182) <= 1; end_W(5, 183) <= 1; 
end_W(5, 184) <= 1; end_W(5, 185) <= 1; end_W(5, 186) <= 1; end_W(5, 187) <= 1; end_W(5, 188) <= 0; end_W(5, 189) <= 0; end_W(5, 190) <= 0; end_W(5, 191) <= 0; 
end_W(5, 192) <= 0; end_W(5, 193) <= 0; end_W(5, 194) <= 0; end_W(5, 195) <= 0; end_W(5, 196) <= 0; end_W(5, 197) <= 0; end_W(5, 198) <= 0; end_W(5, 199) <= 0; 
end_W(5, 200) <= 1; end_W(5, 201) <= 1; end_W(5, 202) <= 1; end_W(5, 203) <= 1; end_W(5, 204) <= 1; end_W(5, 205) <= 1; end_W(5, 206) <= 1; end_W(5, 207) <= 1; 
end_W(5, 208) <= 0; end_W(5, 209) <= 0; end_W(5, 210) <= 0; end_W(5, 211) <= 0; end_W(5, 212) <= 0; end_W(5, 213) <= 0; end_W(5, 214) <= 0; end_W(5, 215) <= 0; 
end_W(5, 216) <= 1; end_W(5, 217) <= 1; end_W(5, 218) <= 1; end_W(5, 219) <= 1; end_W(5, 220) <= 1; end_W(5, 221) <= 1; end_W(5, 222) <= 1; end_W(5, 223) <= 1; 
end_W(5, 224) <= 0; end_W(5, 225) <= 0; end_W(5, 226) <= 0; end_W(5, 227) <= 0; end_W(5, 228) <= 0; end_W(5, 229) <= 0; end_W(5, 230) <= 0; end_W(5, 231) <= 0; 
end_W(5, 232) <= 0; end_W(5, 233) <= 0; end_W(5, 234) <= 0; end_W(5, 235) <= 0; end_W(5, 236) <= 0; end_W(5, 237) <= 0; end_W(5, 238) <= 0; end_W(5, 239) <= 0; 
end_W(5, 240) <= 1; end_W(5, 241) <= 1; end_W(5, 242) <= 1; end_W(5, 243) <= 1; end_W(5, 244) <= 1; end_W(5, 245) <= 1; end_W(5, 246) <= 1; end_W(5, 247) <= 1; 
end_W(5, 248) <= 0; end_W(5, 249) <= 0; end_W(5, 250) <= 0; end_W(5, 251) <= 0; end_W(5, 252) <= 0; end_W(5, 253) <= 0; end_W(5, 254) <= 0; end_W(5, 255) <= 0; 
end_W(5, 256) <= 1; end_W(5, 257) <= 1; end_W(5, 258) <= 1; end_W(5, 259) <= 1; end_W(5, 260) <= 1; end_W(5, 261) <= 1; end_W(5, 262) <= 1; end_W(5, 263) <= 1; 
end_W(5, 264) <= 0; end_W(5, 265) <= 0; end_W(5, 266) <= 0; end_W(5, 267) <= 0; end_W(5, 268) <= 0; end_W(5, 269) <= 0; end_W(5, 270) <= 0; end_W(5, 271) <= 0; 
end_W(5, 272) <= 1; end_W(5, 273) <= 1; end_W(5, 274) <= 1; end_W(5, 275) <= 1; end_W(5, 276) <= 1; end_W(5, 277) <= 1; end_W(5, 278) <= 1; end_W(5, 279) <= 1; 
end_W(5, 280) <= 0; end_W(5, 281) <= 0; end_W(5, 282) <= 0; end_W(5, 283) <= 0; end_W(5, 284) <= 0; end_W(5, 285) <= 0; end_W(5, 286) <= 0; end_W(5, 287) <= 0; 
end_W(5, 288) <= 0; end_W(5, 289) <= 0; end_W(5, 290) <= 0; end_W(5, 291) <= 0; end_W(5, 292) <= 1; end_W(5, 293) <= 1; end_W(5, 294) <= 1; end_W(5, 295) <= 1; 
end_W(5, 296) <= 1; end_W(5, 297) <= 1; end_W(5, 298) <= 1; end_W(5, 299) <= 1; end_W(5, 300) <= 0; end_W(5, 301) <= 0; end_W(5, 302) <= 0; end_W(5, 303) <= 0; 
end_W(5, 304) <= 0; end_W(5, 305) <= 0; end_W(5, 306) <= 0; end_W(5, 307) <= 0; end_W(5, 308) <= 1; end_W(5, 309) <= 1; end_W(5, 310) <= 1; end_W(5, 311) <= 1; 
end_W(5, 312) <= 1; end_W(5, 313) <= 1; end_W(5, 314) <= 1; end_W(5, 315) <= 1; end_W(5, 316) <= 0; end_W(5, 317) <= 0; end_W(5, 318) <= 0; end_W(5, 319) <= 0; 
end_W(5, 320) <= 0; end_W(5, 321) <= 0; end_W(5, 322) <= 0; end_W(5, 323) <= 0; end_W(6, 0) <= 0; end_W(6, 1) <= 0; end_W(6, 2) <= 0; end_W(6, 3) <= 0; end_W(6, 4) <= 1; end_W(6, 5) <= 1; end_W(6, 6) <= 1; end_W(6, 7) <= 1; 
end_W(6, 8) <= 1; end_W(6, 9) <= 1; end_W(6, 10) <= 1; end_W(6, 11) <= 1; end_W(6, 12) <= 0; end_W(6, 13) <= 0; end_W(6, 14) <= 0; end_W(6, 15) <= 0; 
end_W(6, 16) <= 0; end_W(6, 17) <= 0; end_W(6, 18) <= 0; end_W(6, 19) <= 0; end_W(6, 20) <= 1; end_W(6, 21) <= 1; end_W(6, 22) <= 1; end_W(6, 23) <= 1; 
end_W(6, 24) <= 1; end_W(6, 25) <= 1; end_W(6, 26) <= 1; end_W(6, 27) <= 1; end_W(6, 28) <= 0; end_W(6, 29) <= 0; end_W(6, 30) <= 0; end_W(6, 31) <= 0; 
end_W(6, 32) <= 0; end_W(6, 33) <= 0; end_W(6, 34) <= 0; end_W(6, 35) <= 0; end_W(6, 36) <= 0; end_W(6, 37) <= 0; end_W(6, 38) <= 0; end_W(6, 39) <= 0; 
end_W(6, 40) <= 0; end_W(6, 41) <= 0; end_W(6, 42) <= 0; end_W(6, 43) <= 0; end_W(6, 44) <= 1; end_W(6, 45) <= 1; end_W(6, 46) <= 1; end_W(6, 47) <= 1; 
end_W(6, 48) <= 1; end_W(6, 49) <= 1; end_W(6, 50) <= 1; end_W(6, 51) <= 1; end_W(6, 52) <= 1; end_W(6, 53) <= 1; end_W(6, 54) <= 1; end_W(6, 55) <= 1; 
end_W(6, 56) <= 0; end_W(6, 57) <= 0; end_W(6, 58) <= 0; end_W(6, 59) <= 0; end_W(6, 60) <= 0; end_W(6, 61) <= 0; end_W(6, 62) <= 0; end_W(6, 63) <= 0; 
end_W(6, 64) <= 0; end_W(6, 65) <= 0; end_W(6, 66) <= 0; end_W(6, 67) <= 0; end_W(6, 68) <= 0; end_W(6, 69) <= 0; end_W(6, 70) <= 0; end_W(6, 71) <= 0; 
end_W(6, 72) <= 1; end_W(6, 73) <= 1; end_W(6, 74) <= 1; end_W(6, 75) <= 1; end_W(6, 76) <= 1; end_W(6, 77) <= 1; end_W(6, 78) <= 1; end_W(6, 79) <= 1; 
end_W(6, 80) <= 1; end_W(6, 81) <= 1; end_W(6, 82) <= 1; end_W(6, 83) <= 1; end_W(6, 84) <= 0; end_W(6, 85) <= 0; end_W(6, 86) <= 0; end_W(6, 87) <= 0; 
end_W(6, 88) <= 0; end_W(6, 89) <= 0; end_W(6, 90) <= 0; end_W(6, 91) <= 0; end_W(6, 92) <= 1; end_W(6, 93) <= 1; end_W(6, 94) <= 1; end_W(6, 95) <= 1; 
end_W(6, 96) <= 1; end_W(6, 97) <= 1; end_W(6, 98) <= 1; end_W(6, 99) <= 1; end_W(6, 100) <= 1; end_W(6, 101) <= 1; end_W(6, 102) <= 1; end_W(6, 103) <= 1; 
end_W(6, 104) <= 0; end_W(6, 105) <= 0; end_W(6, 106) <= 0; end_W(6, 107) <= 0; end_W(6, 108) <= 0; end_W(6, 109) <= 0; end_W(6, 110) <= 0; end_W(6, 111) <= 0; 
end_W(6, 112) <= 1; end_W(6, 113) <= 1; end_W(6, 114) <= 1; end_W(6, 115) <= 1; end_W(6, 116) <= 1; end_W(6, 117) <= 1; end_W(6, 118) <= 1; end_W(6, 119) <= 1; 
end_W(6, 120) <= 0; end_W(6, 121) <= 0; end_W(6, 122) <= 0; end_W(6, 123) <= 0; end_W(6, 124) <= 0; end_W(6, 125) <= 0; end_W(6, 126) <= 0; end_W(6, 127) <= 0; 
end_W(6, 128) <= 1; end_W(6, 129) <= 1; end_W(6, 130) <= 1; end_W(6, 131) <= 1; end_W(6, 132) <= 1; end_W(6, 133) <= 1; end_W(6, 134) <= 1; end_W(6, 135) <= 1; 
end_W(6, 136) <= 0; end_W(6, 137) <= 0; end_W(6, 138) <= 0; end_W(6, 139) <= 0; end_W(6, 140) <= 0; end_W(6, 141) <= 0; end_W(6, 142) <= 0; end_W(6, 143) <= 0; 
end_W(6, 144) <= 0; end_W(6, 145) <= 0; end_W(6, 146) <= 0; end_W(6, 147) <= 0; end_W(6, 148) <= 0; end_W(6, 149) <= 0; end_W(6, 150) <= 0; end_W(6, 151) <= 0; 
end_W(6, 152) <= 0; end_W(6, 153) <= 0; end_W(6, 154) <= 0; end_W(6, 155) <= 0; end_W(6, 156) <= 0; end_W(6, 157) <= 0; end_W(6, 158) <= 0; end_W(6, 159) <= 0; 
end_W(6, 160) <= 0; end_W(6, 161) <= 0; end_W(6, 162) <= 0; end_W(6, 163) <= 0; end_W(6, 164) <= 0; end_W(6, 165) <= 0; end_W(6, 166) <= 0; end_W(6, 167) <= 0; 
end_W(6, 168) <= 0; end_W(6, 169) <= 0; end_W(6, 170) <= 0; end_W(6, 171) <= 0; end_W(6, 172) <= 0; end_W(6, 173) <= 0; end_W(6, 174) <= 0; end_W(6, 175) <= 0; 
end_W(6, 176) <= 0; end_W(6, 177) <= 0; end_W(6, 178) <= 0; end_W(6, 179) <= 0; end_W(6, 180) <= 1; end_W(6, 181) <= 1; end_W(6, 182) <= 1; end_W(6, 183) <= 1; 
end_W(6, 184) <= 1; end_W(6, 185) <= 1; end_W(6, 186) <= 1; end_W(6, 187) <= 1; end_W(6, 188) <= 0; end_W(6, 189) <= 0; end_W(6, 190) <= 0; end_W(6, 191) <= 0; 
end_W(6, 192) <= 0; end_W(6, 193) <= 0; end_W(6, 194) <= 0; end_W(6, 195) <= 0; end_W(6, 196) <= 0; end_W(6, 197) <= 0; end_W(6, 198) <= 0; end_W(6, 199) <= 0; 
end_W(6, 200) <= 1; end_W(6, 201) <= 1; end_W(6, 202) <= 1; end_W(6, 203) <= 1; end_W(6, 204) <= 1; end_W(6, 205) <= 1; end_W(6, 206) <= 1; end_W(6, 207) <= 1; 
end_W(6, 208) <= 0; end_W(6, 209) <= 0; end_W(6, 210) <= 0; end_W(6, 211) <= 0; end_W(6, 212) <= 0; end_W(6, 213) <= 0; end_W(6, 214) <= 0; end_W(6, 215) <= 0; 
end_W(6, 216) <= 1; end_W(6, 217) <= 1; end_W(6, 218) <= 1; end_W(6, 219) <= 1; end_W(6, 220) <= 1; end_W(6, 221) <= 1; end_W(6, 222) <= 1; end_W(6, 223) <= 1; 
end_W(6, 224) <= 0; end_W(6, 225) <= 0; end_W(6, 226) <= 0; end_W(6, 227) <= 0; end_W(6, 228) <= 0; end_W(6, 229) <= 0; end_W(6, 230) <= 0; end_W(6, 231) <= 0; 
end_W(6, 232) <= 0; end_W(6, 233) <= 0; end_W(6, 234) <= 0; end_W(6, 235) <= 0; end_W(6, 236) <= 0; end_W(6, 237) <= 0; end_W(6, 238) <= 0; end_W(6, 239) <= 0; 
end_W(6, 240) <= 1; end_W(6, 241) <= 1; end_W(6, 242) <= 1; end_W(6, 243) <= 1; end_W(6, 244) <= 1; end_W(6, 245) <= 1; end_W(6, 246) <= 1; end_W(6, 247) <= 1; 
end_W(6, 248) <= 0; end_W(6, 249) <= 0; end_W(6, 250) <= 0; end_W(6, 251) <= 0; end_W(6, 252) <= 0; end_W(6, 253) <= 0; end_W(6, 254) <= 0; end_W(6, 255) <= 0; 
end_W(6, 256) <= 1; end_W(6, 257) <= 1; end_W(6, 258) <= 1; end_W(6, 259) <= 1; end_W(6, 260) <= 1; end_W(6, 261) <= 1; end_W(6, 262) <= 1; end_W(6, 263) <= 1; 
end_W(6, 264) <= 0; end_W(6, 265) <= 0; end_W(6, 266) <= 0; end_W(6, 267) <= 0; end_W(6, 268) <= 0; end_W(6, 269) <= 0; end_W(6, 270) <= 0; end_W(6, 271) <= 0; 
end_W(6, 272) <= 1; end_W(6, 273) <= 1; end_W(6, 274) <= 1; end_W(6, 275) <= 1; end_W(6, 276) <= 1; end_W(6, 277) <= 1; end_W(6, 278) <= 1; end_W(6, 279) <= 1; 
end_W(6, 280) <= 0; end_W(6, 281) <= 0; end_W(6, 282) <= 0; end_W(6, 283) <= 0; end_W(6, 284) <= 0; end_W(6, 285) <= 0; end_W(6, 286) <= 0; end_W(6, 287) <= 0; 
end_W(6, 288) <= 0; end_W(6, 289) <= 0; end_W(6, 290) <= 0; end_W(6, 291) <= 0; end_W(6, 292) <= 1; end_W(6, 293) <= 1; end_W(6, 294) <= 1; end_W(6, 295) <= 1; 
end_W(6, 296) <= 1; end_W(6, 297) <= 1; end_W(6, 298) <= 1; end_W(6, 299) <= 1; end_W(6, 300) <= 0; end_W(6, 301) <= 0; end_W(6, 302) <= 0; end_W(6, 303) <= 0; 
end_W(6, 304) <= 0; end_W(6, 305) <= 0; end_W(6, 306) <= 0; end_W(6, 307) <= 0; end_W(6, 308) <= 1; end_W(6, 309) <= 1; end_W(6, 310) <= 1; end_W(6, 311) <= 1; 
end_W(6, 312) <= 1; end_W(6, 313) <= 1; end_W(6, 314) <= 1; end_W(6, 315) <= 1; end_W(6, 316) <= 0; end_W(6, 317) <= 0; end_W(6, 318) <= 0; end_W(6, 319) <= 0; 
end_W(6, 320) <= 0; end_W(6, 321) <= 0; end_W(6, 322) <= 0; end_W(6, 323) <= 0; end_W(7, 0) <= 0; end_W(7, 1) <= 0; end_W(7, 2) <= 0; end_W(7, 3) <= 0; end_W(7, 4) <= 1; end_W(7, 5) <= 1; end_W(7, 6) <= 1; end_W(7, 7) <= 1; 
end_W(7, 8) <= 1; end_W(7, 9) <= 1; end_W(7, 10) <= 1; end_W(7, 11) <= 1; end_W(7, 12) <= 0; end_W(7, 13) <= 0; end_W(7, 14) <= 0; end_W(7, 15) <= 0; 
end_W(7, 16) <= 0; end_W(7, 17) <= 0; end_W(7, 18) <= 0; end_W(7, 19) <= 0; end_W(7, 20) <= 1; end_W(7, 21) <= 1; end_W(7, 22) <= 1; end_W(7, 23) <= 1; 
end_W(7, 24) <= 1; end_W(7, 25) <= 1; end_W(7, 26) <= 1; end_W(7, 27) <= 1; end_W(7, 28) <= 0; end_W(7, 29) <= 0; end_W(7, 30) <= 0; end_W(7, 31) <= 0; 
end_W(7, 32) <= 0; end_W(7, 33) <= 0; end_W(7, 34) <= 0; end_W(7, 35) <= 0; end_W(7, 36) <= 0; end_W(7, 37) <= 0; end_W(7, 38) <= 0; end_W(7, 39) <= 0; 
end_W(7, 40) <= 0; end_W(7, 41) <= 0; end_W(7, 42) <= 0; end_W(7, 43) <= 0; end_W(7, 44) <= 1; end_W(7, 45) <= 1; end_W(7, 46) <= 1; end_W(7, 47) <= 1; 
end_W(7, 48) <= 1; end_W(7, 49) <= 1; end_W(7, 50) <= 1; end_W(7, 51) <= 1; end_W(7, 52) <= 1; end_W(7, 53) <= 1; end_W(7, 54) <= 1; end_W(7, 55) <= 1; 
end_W(7, 56) <= 0; end_W(7, 57) <= 0; end_W(7, 58) <= 0; end_W(7, 59) <= 0; end_W(7, 60) <= 0; end_W(7, 61) <= 0; end_W(7, 62) <= 0; end_W(7, 63) <= 0; 
end_W(7, 64) <= 0; end_W(7, 65) <= 0; end_W(7, 66) <= 0; end_W(7, 67) <= 0; end_W(7, 68) <= 0; end_W(7, 69) <= 0; end_W(7, 70) <= 0; end_W(7, 71) <= 0; 
end_W(7, 72) <= 1; end_W(7, 73) <= 1; end_W(7, 74) <= 1; end_W(7, 75) <= 1; end_W(7, 76) <= 1; end_W(7, 77) <= 1; end_W(7, 78) <= 1; end_W(7, 79) <= 1; 
end_W(7, 80) <= 1; end_W(7, 81) <= 1; end_W(7, 82) <= 1; end_W(7, 83) <= 1; end_W(7, 84) <= 0; end_W(7, 85) <= 0; end_W(7, 86) <= 0; end_W(7, 87) <= 0; 
end_W(7, 88) <= 0; end_W(7, 89) <= 0; end_W(7, 90) <= 0; end_W(7, 91) <= 0; end_W(7, 92) <= 1; end_W(7, 93) <= 1; end_W(7, 94) <= 1; end_W(7, 95) <= 1; 
end_W(7, 96) <= 1; end_W(7, 97) <= 1; end_W(7, 98) <= 1; end_W(7, 99) <= 1; end_W(7, 100) <= 1; end_W(7, 101) <= 1; end_W(7, 102) <= 1; end_W(7, 103) <= 1; 
end_W(7, 104) <= 0; end_W(7, 105) <= 0; end_W(7, 106) <= 0; end_W(7, 107) <= 0; end_W(7, 108) <= 0; end_W(7, 109) <= 0; end_W(7, 110) <= 0; end_W(7, 111) <= 0; 
end_W(7, 112) <= 1; end_W(7, 113) <= 1; end_W(7, 114) <= 1; end_W(7, 115) <= 1; end_W(7, 116) <= 1; end_W(7, 117) <= 1; end_W(7, 118) <= 1; end_W(7, 119) <= 1; 
end_W(7, 120) <= 0; end_W(7, 121) <= 0; end_W(7, 122) <= 0; end_W(7, 123) <= 0; end_W(7, 124) <= 0; end_W(7, 125) <= 0; end_W(7, 126) <= 0; end_W(7, 127) <= 0; 
end_W(7, 128) <= 1; end_W(7, 129) <= 1; end_W(7, 130) <= 1; end_W(7, 131) <= 1; end_W(7, 132) <= 1; end_W(7, 133) <= 1; end_W(7, 134) <= 1; end_W(7, 135) <= 1; 
end_W(7, 136) <= 0; end_W(7, 137) <= 0; end_W(7, 138) <= 0; end_W(7, 139) <= 0; end_W(7, 140) <= 0; end_W(7, 141) <= 0; end_W(7, 142) <= 0; end_W(7, 143) <= 0; 
end_W(7, 144) <= 0; end_W(7, 145) <= 0; end_W(7, 146) <= 0; end_W(7, 147) <= 0; end_W(7, 148) <= 0; end_W(7, 149) <= 0; end_W(7, 150) <= 0; end_W(7, 151) <= 0; 
end_W(7, 152) <= 0; end_W(7, 153) <= 0; end_W(7, 154) <= 0; end_W(7, 155) <= 0; end_W(7, 156) <= 0; end_W(7, 157) <= 0; end_W(7, 158) <= 0; end_W(7, 159) <= 0; 
end_W(7, 160) <= 0; end_W(7, 161) <= 0; end_W(7, 162) <= 0; end_W(7, 163) <= 0; end_W(7, 164) <= 0; end_W(7, 165) <= 0; end_W(7, 166) <= 0; end_W(7, 167) <= 0; 
end_W(7, 168) <= 0; end_W(7, 169) <= 0; end_W(7, 170) <= 0; end_W(7, 171) <= 0; end_W(7, 172) <= 0; end_W(7, 173) <= 0; end_W(7, 174) <= 0; end_W(7, 175) <= 0; 
end_W(7, 176) <= 0; end_W(7, 177) <= 0; end_W(7, 178) <= 0; end_W(7, 179) <= 0; end_W(7, 180) <= 1; end_W(7, 181) <= 1; end_W(7, 182) <= 1; end_W(7, 183) <= 1; 
end_W(7, 184) <= 1; end_W(7, 185) <= 1; end_W(7, 186) <= 1; end_W(7, 187) <= 1; end_W(7, 188) <= 0; end_W(7, 189) <= 0; end_W(7, 190) <= 0; end_W(7, 191) <= 0; 
end_W(7, 192) <= 0; end_W(7, 193) <= 0; end_W(7, 194) <= 0; end_W(7, 195) <= 0; end_W(7, 196) <= 0; end_W(7, 197) <= 0; end_W(7, 198) <= 0; end_W(7, 199) <= 0; 
end_W(7, 200) <= 1; end_W(7, 201) <= 1; end_W(7, 202) <= 1; end_W(7, 203) <= 1; end_W(7, 204) <= 1; end_W(7, 205) <= 1; end_W(7, 206) <= 1; end_W(7, 207) <= 1; 
end_W(7, 208) <= 0; end_W(7, 209) <= 0; end_W(7, 210) <= 0; end_W(7, 211) <= 0; end_W(7, 212) <= 0; end_W(7, 213) <= 0; end_W(7, 214) <= 0; end_W(7, 215) <= 0; 
end_W(7, 216) <= 1; end_W(7, 217) <= 1; end_W(7, 218) <= 1; end_W(7, 219) <= 1; end_W(7, 220) <= 1; end_W(7, 221) <= 1; end_W(7, 222) <= 1; end_W(7, 223) <= 1; 
end_W(7, 224) <= 0; end_W(7, 225) <= 0; end_W(7, 226) <= 0; end_W(7, 227) <= 0; end_W(7, 228) <= 0; end_W(7, 229) <= 0; end_W(7, 230) <= 0; end_W(7, 231) <= 0; 
end_W(7, 232) <= 0; end_W(7, 233) <= 0; end_W(7, 234) <= 0; end_W(7, 235) <= 0; end_W(7, 236) <= 0; end_W(7, 237) <= 0; end_W(7, 238) <= 0; end_W(7, 239) <= 0; 
end_W(7, 240) <= 1; end_W(7, 241) <= 1; end_W(7, 242) <= 1; end_W(7, 243) <= 1; end_W(7, 244) <= 1; end_W(7, 245) <= 1; end_W(7, 246) <= 1; end_W(7, 247) <= 1; 
end_W(7, 248) <= 0; end_W(7, 249) <= 0; end_W(7, 250) <= 0; end_W(7, 251) <= 0; end_W(7, 252) <= 0; end_W(7, 253) <= 0; end_W(7, 254) <= 0; end_W(7, 255) <= 0; 
end_W(7, 256) <= 1; end_W(7, 257) <= 1; end_W(7, 258) <= 1; end_W(7, 259) <= 1; end_W(7, 260) <= 1; end_W(7, 261) <= 1; end_W(7, 262) <= 1; end_W(7, 263) <= 1; 
end_W(7, 264) <= 0; end_W(7, 265) <= 0; end_W(7, 266) <= 0; end_W(7, 267) <= 0; end_W(7, 268) <= 0; end_W(7, 269) <= 0; end_W(7, 270) <= 0; end_W(7, 271) <= 0; 
end_W(7, 272) <= 1; end_W(7, 273) <= 1; end_W(7, 274) <= 1; end_W(7, 275) <= 1; end_W(7, 276) <= 1; end_W(7, 277) <= 1; end_W(7, 278) <= 1; end_W(7, 279) <= 1; 
end_W(7, 280) <= 0; end_W(7, 281) <= 0; end_W(7, 282) <= 0; end_W(7, 283) <= 0; end_W(7, 284) <= 0; end_W(7, 285) <= 0; end_W(7, 286) <= 0; end_W(7, 287) <= 0; 
end_W(7, 288) <= 0; end_W(7, 289) <= 0; end_W(7, 290) <= 0; end_W(7, 291) <= 0; end_W(7, 292) <= 1; end_W(7, 293) <= 1; end_W(7, 294) <= 1; end_W(7, 295) <= 1; 
end_W(7, 296) <= 1; end_W(7, 297) <= 1; end_W(7, 298) <= 1; end_W(7, 299) <= 1; end_W(7, 300) <= 0; end_W(7, 301) <= 0; end_W(7, 302) <= 0; end_W(7, 303) <= 0; 
end_W(7, 304) <= 0; end_W(7, 305) <= 0; end_W(7, 306) <= 0; end_W(7, 307) <= 0; end_W(7, 308) <= 1; end_W(7, 309) <= 1; end_W(7, 310) <= 1; end_W(7, 311) <= 1; 
end_W(7, 312) <= 1; end_W(7, 313) <= 1; end_W(7, 314) <= 1; end_W(7, 315) <= 1; end_W(7, 316) <= 0; end_W(7, 317) <= 0; end_W(7, 318) <= 0; end_W(7, 319) <= 0; 
end_W(7, 320) <= 0; end_W(7, 321) <= 0; end_W(7, 322) <= 0; end_W(7, 323) <= 0; end_W(8, 0) <= 1; end_W(8, 1) <= 1; end_W(8, 2) <= 1; end_W(8, 3) <= 1; end_W(8, 4) <= 1; end_W(8, 5) <= 1; end_W(8, 6) <= 1; end_W(8, 7) <= 1; 
end_W(8, 8) <= 0; end_W(8, 9) <= 0; end_W(8, 10) <= 0; end_W(8, 11) <= 0; end_W(8, 12) <= 0; end_W(8, 13) <= 0; end_W(8, 14) <= 0; end_W(8, 15) <= 0; 
end_W(8, 16) <= 0; end_W(8, 17) <= 0; end_W(8, 18) <= 0; end_W(8, 19) <= 0; end_W(8, 20) <= 0; end_W(8, 21) <= 0; end_W(8, 22) <= 0; end_W(8, 23) <= 0; 
end_W(8, 24) <= 1; end_W(8, 25) <= 1; end_W(8, 26) <= 1; end_W(8, 27) <= 1; end_W(8, 28) <= 0; end_W(8, 29) <= 0; end_W(8, 30) <= 0; end_W(8, 31) <= 0; 
end_W(8, 32) <= 0; end_W(8, 33) <= 0; end_W(8, 34) <= 0; end_W(8, 35) <= 0; end_W(8, 36) <= 0; end_W(8, 37) <= 0; end_W(8, 38) <= 0; end_W(8, 39) <= 0; 
end_W(8, 40) <= 1; end_W(8, 41) <= 1; end_W(8, 42) <= 1; end_W(8, 43) <= 1; end_W(8, 44) <= 1; end_W(8, 45) <= 1; end_W(8, 46) <= 1; end_W(8, 47) <= 1; 
end_W(8, 48) <= 0; end_W(8, 49) <= 0; end_W(8, 50) <= 0; end_W(8, 51) <= 0; end_W(8, 52) <= 1; end_W(8, 53) <= 1; end_W(8, 54) <= 1; end_W(8, 55) <= 1; 
end_W(8, 56) <= 1; end_W(8, 57) <= 1; end_W(8, 58) <= 1; end_W(8, 59) <= 1; end_W(8, 60) <= 0; end_W(8, 61) <= 0; end_W(8, 62) <= 0; end_W(8, 63) <= 0; 
end_W(8, 64) <= 0; end_W(8, 65) <= 0; end_W(8, 66) <= 0; end_W(8, 67) <= 0; end_W(8, 68) <= 0; end_W(8, 69) <= 0; end_W(8, 70) <= 0; end_W(8, 71) <= 0; 
end_W(8, 72) <= 1; end_W(8, 73) <= 1; end_W(8, 74) <= 1; end_W(8, 75) <= 1; end_W(8, 76) <= 1; end_W(8, 77) <= 1; end_W(8, 78) <= 1; end_W(8, 79) <= 1; 
end_W(8, 80) <= 1; end_W(8, 81) <= 1; end_W(8, 82) <= 1; end_W(8, 83) <= 1; end_W(8, 84) <= 1; end_W(8, 85) <= 1; end_W(8, 86) <= 1; end_W(8, 87) <= 1; 
end_W(8, 88) <= 1; end_W(8, 89) <= 1; end_W(8, 90) <= 1; end_W(8, 91) <= 1; end_W(8, 92) <= 1; end_W(8, 93) <= 1; end_W(8, 94) <= 1; end_W(8, 95) <= 1; 
end_W(8, 96) <= 1; end_W(8, 97) <= 1; end_W(8, 98) <= 1; end_W(8, 99) <= 1; end_W(8, 100) <= 1; end_W(8, 101) <= 1; end_W(8, 102) <= 1; end_W(8, 103) <= 1; 
end_W(8, 104) <= 0; end_W(8, 105) <= 0; end_W(8, 106) <= 0; end_W(8, 107) <= 0; end_W(8, 108) <= 0; end_W(8, 109) <= 0; end_W(8, 110) <= 0; end_W(8, 111) <= 0; 
end_W(8, 112) <= 1; end_W(8, 113) <= 1; end_W(8, 114) <= 1; end_W(8, 115) <= 1; end_W(8, 116) <= 1; end_W(8, 117) <= 1; end_W(8, 118) <= 1; end_W(8, 119) <= 1; 
end_W(8, 120) <= 0; end_W(8, 121) <= 0; end_W(8, 122) <= 0; end_W(8, 123) <= 0; end_W(8, 124) <= 0; end_W(8, 125) <= 0; end_W(8, 126) <= 0; end_W(8, 127) <= 0; 
end_W(8, 128) <= 0; end_W(8, 129) <= 0; end_W(8, 130) <= 0; end_W(8, 131) <= 0; end_W(8, 132) <= 1; end_W(8, 133) <= 1; end_W(8, 134) <= 1; end_W(8, 135) <= 1; 
end_W(8, 136) <= 0; end_W(8, 137) <= 0; end_W(8, 138) <= 0; end_W(8, 139) <= 0; end_W(8, 140) <= 0; end_W(8, 141) <= 0; end_W(8, 142) <= 0; end_W(8, 143) <= 0; 
end_W(8, 144) <= 0; end_W(8, 145) <= 0; end_W(8, 146) <= 0; end_W(8, 147) <= 0; end_W(8, 148) <= 0; end_W(8, 149) <= 0; end_W(8, 150) <= 0; end_W(8, 151) <= 0; 
end_W(8, 152) <= 0; end_W(8, 153) <= 0; end_W(8, 154) <= 0; end_W(8, 155) <= 0; end_W(8, 156) <= 0; end_W(8, 157) <= 0; end_W(8, 158) <= 0; end_W(8, 159) <= 0; 
end_W(8, 160) <= 0; end_W(8, 161) <= 0; end_W(8, 162) <= 0; end_W(8, 163) <= 0; end_W(8, 164) <= 0; end_W(8, 165) <= 0; end_W(8, 166) <= 0; end_W(8, 167) <= 0; 
end_W(8, 168) <= 0; end_W(8, 169) <= 0; end_W(8, 170) <= 0; end_W(8, 171) <= 0; end_W(8, 172) <= 0; end_W(8, 173) <= 0; end_W(8, 174) <= 0; end_W(8, 175) <= 0; 
end_W(8, 176) <= 0; end_W(8, 177) <= 0; end_W(8, 178) <= 0; end_W(8, 179) <= 0; end_W(8, 180) <= 1; end_W(8, 181) <= 1; end_W(8, 182) <= 1; end_W(8, 183) <= 1; 
end_W(8, 184) <= 1; end_W(8, 185) <= 1; end_W(8, 186) <= 1; end_W(8, 187) <= 1; end_W(8, 188) <= 0; end_W(8, 189) <= 0; end_W(8, 190) <= 0; end_W(8, 191) <= 0; 
end_W(8, 192) <= 0; end_W(8, 193) <= 0; end_W(8, 194) <= 0; end_W(8, 195) <= 0; end_W(8, 196) <= 0; end_W(8, 197) <= 0; end_W(8, 198) <= 0; end_W(8, 199) <= 0; 
end_W(8, 200) <= 1; end_W(8, 201) <= 1; end_W(8, 202) <= 1; end_W(8, 203) <= 1; end_W(8, 204) <= 1; end_W(8, 205) <= 1; end_W(8, 206) <= 1; end_W(8, 207) <= 1; 
end_W(8, 208) <= 0; end_W(8, 209) <= 0; end_W(8, 210) <= 0; end_W(8, 211) <= 0; end_W(8, 212) <= 0; end_W(8, 213) <= 0; end_W(8, 214) <= 0; end_W(8, 215) <= 0; 
end_W(8, 216) <= 1; end_W(8, 217) <= 1; end_W(8, 218) <= 1; end_W(8, 219) <= 1; end_W(8, 220) <= 1; end_W(8, 221) <= 1; end_W(8, 222) <= 1; end_W(8, 223) <= 1; 
end_W(8, 224) <= 0; end_W(8, 225) <= 0; end_W(8, 226) <= 0; end_W(8, 227) <= 0; end_W(8, 228) <= 0; end_W(8, 229) <= 0; end_W(8, 230) <= 0; end_W(8, 231) <= 0; 
end_W(8, 232) <= 0; end_W(8, 233) <= 0; end_W(8, 234) <= 0; end_W(8, 235) <= 0; end_W(8, 236) <= 0; end_W(8, 237) <= 0; end_W(8, 238) <= 0; end_W(8, 239) <= 0; 
end_W(8, 240) <= 1; end_W(8, 241) <= 1; end_W(8, 242) <= 1; end_W(8, 243) <= 1; end_W(8, 244) <= 1; end_W(8, 245) <= 1; end_W(8, 246) <= 1; end_W(8, 247) <= 1; 
end_W(8, 248) <= 0; end_W(8, 249) <= 0; end_W(8, 250) <= 0; end_W(8, 251) <= 0; end_W(8, 252) <= 0; end_W(8, 253) <= 0; end_W(8, 254) <= 0; end_W(8, 255) <= 0; 
end_W(8, 256) <= 1; end_W(8, 257) <= 1; end_W(8, 258) <= 1; end_W(8, 259) <= 1; end_W(8, 260) <= 1; end_W(8, 261) <= 1; end_W(8, 262) <= 1; end_W(8, 263) <= 1; 
end_W(8, 264) <= 0; end_W(8, 265) <= 0; end_W(8, 266) <= 0; end_W(8, 267) <= 0; end_W(8, 268) <= 0; end_W(8, 269) <= 0; end_W(8, 270) <= 0; end_W(8, 271) <= 0; 
end_W(8, 272) <= 0; end_W(8, 273) <= 0; end_W(8, 274) <= 0; end_W(8, 275) <= 0; end_W(8, 276) <= 1; end_W(8, 277) <= 1; end_W(8, 278) <= 1; end_W(8, 279) <= 1; 
end_W(8, 280) <= 0; end_W(8, 281) <= 0; end_W(8, 282) <= 0; end_W(8, 283) <= 0; end_W(8, 284) <= 0; end_W(8, 285) <= 0; end_W(8, 286) <= 0; end_W(8, 287) <= 0; 
end_W(8, 288) <= 0; end_W(8, 289) <= 0; end_W(8, 290) <= 0; end_W(8, 291) <= 0; end_W(8, 292) <= 1; end_W(8, 293) <= 1; end_W(8, 294) <= 1; end_W(8, 295) <= 1; 
end_W(8, 296) <= 1; end_W(8, 297) <= 1; end_W(8, 298) <= 1; end_W(8, 299) <= 1; end_W(8, 300) <= 0; end_W(8, 301) <= 0; end_W(8, 302) <= 0; end_W(8, 303) <= 0; 
end_W(8, 304) <= 0; end_W(8, 305) <= 0; end_W(8, 306) <= 0; end_W(8, 307) <= 0; end_W(8, 308) <= 1; end_W(8, 309) <= 1; end_W(8, 310) <= 1; end_W(8, 311) <= 1; 
end_W(8, 312) <= 1; end_W(8, 313) <= 1; end_W(8, 314) <= 1; end_W(8, 315) <= 1; end_W(8, 316) <= 0; end_W(8, 317) <= 0; end_W(8, 318) <= 0; end_W(8, 319) <= 0; 
end_W(8, 320) <= 0; end_W(8, 321) <= 0; end_W(8, 322) <= 0; end_W(8, 323) <= 0; end_W(9, 0) <= 1; end_W(9, 1) <= 1; end_W(9, 2) <= 1; end_W(9, 3) <= 1; end_W(9, 4) <= 1; end_W(9, 5) <= 1; end_W(9, 6) <= 1; end_W(9, 7) <= 1; 
end_W(9, 8) <= 0; end_W(9, 9) <= 0; end_W(9, 10) <= 0; end_W(9, 11) <= 0; end_W(9, 12) <= 0; end_W(9, 13) <= 0; end_W(9, 14) <= 0; end_W(9, 15) <= 0; 
end_W(9, 16) <= 0; end_W(9, 17) <= 0; end_W(9, 18) <= 0; end_W(9, 19) <= 0; end_W(9, 20) <= 0; end_W(9, 21) <= 0; end_W(9, 22) <= 0; end_W(9, 23) <= 0; 
end_W(9, 24) <= 1; end_W(9, 25) <= 1; end_W(9, 26) <= 1; end_W(9, 27) <= 1; end_W(9, 28) <= 0; end_W(9, 29) <= 0; end_W(9, 30) <= 0; end_W(9, 31) <= 0; 
end_W(9, 32) <= 0; end_W(9, 33) <= 0; end_W(9, 34) <= 0; end_W(9, 35) <= 0; end_W(9, 36) <= 0; end_W(9, 37) <= 0; end_W(9, 38) <= 0; end_W(9, 39) <= 0; 
end_W(9, 40) <= 1; end_W(9, 41) <= 1; end_W(9, 42) <= 1; end_W(9, 43) <= 1; end_W(9, 44) <= 1; end_W(9, 45) <= 1; end_W(9, 46) <= 1; end_W(9, 47) <= 1; 
end_W(9, 48) <= 0; end_W(9, 49) <= 0; end_W(9, 50) <= 0; end_W(9, 51) <= 0; end_W(9, 52) <= 1; end_W(9, 53) <= 1; end_W(9, 54) <= 1; end_W(9, 55) <= 1; 
end_W(9, 56) <= 1; end_W(9, 57) <= 1; end_W(9, 58) <= 1; end_W(9, 59) <= 1; end_W(9, 60) <= 0; end_W(9, 61) <= 0; end_W(9, 62) <= 0; end_W(9, 63) <= 0; 
end_W(9, 64) <= 0; end_W(9, 65) <= 0; end_W(9, 66) <= 0; end_W(9, 67) <= 0; end_W(9, 68) <= 0; end_W(9, 69) <= 0; end_W(9, 70) <= 0; end_W(9, 71) <= 0; 
end_W(9, 72) <= 1; end_W(9, 73) <= 1; end_W(9, 74) <= 1; end_W(9, 75) <= 1; end_W(9, 76) <= 1; end_W(9, 77) <= 1; end_W(9, 78) <= 1; end_W(9, 79) <= 1; 
end_W(9, 80) <= 1; end_W(9, 81) <= 1; end_W(9, 82) <= 1; end_W(9, 83) <= 1; end_W(9, 84) <= 1; end_W(9, 85) <= 1; end_W(9, 86) <= 1; end_W(9, 87) <= 1; 
end_W(9, 88) <= 1; end_W(9, 89) <= 1; end_W(9, 90) <= 1; end_W(9, 91) <= 1; end_W(9, 92) <= 1; end_W(9, 93) <= 1; end_W(9, 94) <= 1; end_W(9, 95) <= 1; 
end_W(9, 96) <= 1; end_W(9, 97) <= 1; end_W(9, 98) <= 1; end_W(9, 99) <= 1; end_W(9, 100) <= 1; end_W(9, 101) <= 1; end_W(9, 102) <= 1; end_W(9, 103) <= 1; 
end_W(9, 104) <= 0; end_W(9, 105) <= 0; end_W(9, 106) <= 0; end_W(9, 107) <= 0; end_W(9, 108) <= 0; end_W(9, 109) <= 0; end_W(9, 110) <= 0; end_W(9, 111) <= 0; 
end_W(9, 112) <= 1; end_W(9, 113) <= 1; end_W(9, 114) <= 1; end_W(9, 115) <= 1; end_W(9, 116) <= 1; end_W(9, 117) <= 1; end_W(9, 118) <= 1; end_W(9, 119) <= 1; 
end_W(9, 120) <= 0; end_W(9, 121) <= 0; end_W(9, 122) <= 0; end_W(9, 123) <= 0; end_W(9, 124) <= 0; end_W(9, 125) <= 0; end_W(9, 126) <= 0; end_W(9, 127) <= 0; 
end_W(9, 128) <= 0; end_W(9, 129) <= 0; end_W(9, 130) <= 0; end_W(9, 131) <= 0; end_W(9, 132) <= 1; end_W(9, 133) <= 1; end_W(9, 134) <= 1; end_W(9, 135) <= 1; 
end_W(9, 136) <= 0; end_W(9, 137) <= 0; end_W(9, 138) <= 0; end_W(9, 139) <= 0; end_W(9, 140) <= 0; end_W(9, 141) <= 0; end_W(9, 142) <= 0; end_W(9, 143) <= 0; 
end_W(9, 144) <= 0; end_W(9, 145) <= 0; end_W(9, 146) <= 0; end_W(9, 147) <= 0; end_W(9, 148) <= 0; end_W(9, 149) <= 0; end_W(9, 150) <= 0; end_W(9, 151) <= 0; 
end_W(9, 152) <= 0; end_W(9, 153) <= 0; end_W(9, 154) <= 0; end_W(9, 155) <= 0; end_W(9, 156) <= 0; end_W(9, 157) <= 0; end_W(9, 158) <= 0; end_W(9, 159) <= 0; 
end_W(9, 160) <= 0; end_W(9, 161) <= 0; end_W(9, 162) <= 0; end_W(9, 163) <= 0; end_W(9, 164) <= 0; end_W(9, 165) <= 0; end_W(9, 166) <= 0; end_W(9, 167) <= 0; 
end_W(9, 168) <= 0; end_W(9, 169) <= 0; end_W(9, 170) <= 0; end_W(9, 171) <= 0; end_W(9, 172) <= 0; end_W(9, 173) <= 0; end_W(9, 174) <= 0; end_W(9, 175) <= 0; 
end_W(9, 176) <= 0; end_W(9, 177) <= 0; end_W(9, 178) <= 0; end_W(9, 179) <= 0; end_W(9, 180) <= 1; end_W(9, 181) <= 1; end_W(9, 182) <= 1; end_W(9, 183) <= 1; 
end_W(9, 184) <= 1; end_W(9, 185) <= 1; end_W(9, 186) <= 1; end_W(9, 187) <= 1; end_W(9, 188) <= 0; end_W(9, 189) <= 0; end_W(9, 190) <= 0; end_W(9, 191) <= 0; 
end_W(9, 192) <= 0; end_W(9, 193) <= 0; end_W(9, 194) <= 0; end_W(9, 195) <= 0; end_W(9, 196) <= 0; end_W(9, 197) <= 0; end_W(9, 198) <= 0; end_W(9, 199) <= 0; 
end_W(9, 200) <= 1; end_W(9, 201) <= 1; end_W(9, 202) <= 1; end_W(9, 203) <= 1; end_W(9, 204) <= 1; end_W(9, 205) <= 1; end_W(9, 206) <= 1; end_W(9, 207) <= 1; 
end_W(9, 208) <= 0; end_W(9, 209) <= 0; end_W(9, 210) <= 0; end_W(9, 211) <= 0; end_W(9, 212) <= 0; end_W(9, 213) <= 0; end_W(9, 214) <= 0; end_W(9, 215) <= 0; 
end_W(9, 216) <= 1; end_W(9, 217) <= 1; end_W(9, 218) <= 1; end_W(9, 219) <= 1; end_W(9, 220) <= 1; end_W(9, 221) <= 1; end_W(9, 222) <= 1; end_W(9, 223) <= 1; 
end_W(9, 224) <= 0; end_W(9, 225) <= 0; end_W(9, 226) <= 0; end_W(9, 227) <= 0; end_W(9, 228) <= 0; end_W(9, 229) <= 0; end_W(9, 230) <= 0; end_W(9, 231) <= 0; 
end_W(9, 232) <= 0; end_W(9, 233) <= 0; end_W(9, 234) <= 0; end_W(9, 235) <= 0; end_W(9, 236) <= 0; end_W(9, 237) <= 0; end_W(9, 238) <= 0; end_W(9, 239) <= 0; 
end_W(9, 240) <= 1; end_W(9, 241) <= 1; end_W(9, 242) <= 1; end_W(9, 243) <= 1; end_W(9, 244) <= 1; end_W(9, 245) <= 1; end_W(9, 246) <= 1; end_W(9, 247) <= 1; 
end_W(9, 248) <= 0; end_W(9, 249) <= 0; end_W(9, 250) <= 0; end_W(9, 251) <= 0; end_W(9, 252) <= 0; end_W(9, 253) <= 0; end_W(9, 254) <= 0; end_W(9, 255) <= 0; 
end_W(9, 256) <= 1; end_W(9, 257) <= 1; end_W(9, 258) <= 1; end_W(9, 259) <= 1; end_W(9, 260) <= 1; end_W(9, 261) <= 1; end_W(9, 262) <= 1; end_W(9, 263) <= 1; 
end_W(9, 264) <= 0; end_W(9, 265) <= 0; end_W(9, 266) <= 0; end_W(9, 267) <= 0; end_W(9, 268) <= 0; end_W(9, 269) <= 0; end_W(9, 270) <= 0; end_W(9, 271) <= 0; 
end_W(9, 272) <= 0; end_W(9, 273) <= 0; end_W(9, 274) <= 0; end_W(9, 275) <= 0; end_W(9, 276) <= 1; end_W(9, 277) <= 1; end_W(9, 278) <= 1; end_W(9, 279) <= 1; 
end_W(9, 280) <= 0; end_W(9, 281) <= 0; end_W(9, 282) <= 0; end_W(9, 283) <= 0; end_W(9, 284) <= 0; end_W(9, 285) <= 0; end_W(9, 286) <= 0; end_W(9, 287) <= 0; 
end_W(9, 288) <= 0; end_W(9, 289) <= 0; end_W(9, 290) <= 0; end_W(9, 291) <= 0; end_W(9, 292) <= 1; end_W(9, 293) <= 1; end_W(9, 294) <= 1; end_W(9, 295) <= 1; 
end_W(9, 296) <= 1; end_W(9, 297) <= 1; end_W(9, 298) <= 1; end_W(9, 299) <= 1; end_W(9, 300) <= 0; end_W(9, 301) <= 0; end_W(9, 302) <= 0; end_W(9, 303) <= 0; 
end_W(9, 304) <= 0; end_W(9, 305) <= 0; end_W(9, 306) <= 0; end_W(9, 307) <= 0; end_W(9, 308) <= 1; end_W(9, 309) <= 1; end_W(9, 310) <= 1; end_W(9, 311) <= 1; 
end_W(9, 312) <= 1; end_W(9, 313) <= 1; end_W(9, 314) <= 1; end_W(9, 315) <= 1; end_W(9, 316) <= 0; end_W(9, 317) <= 0; end_W(9, 318) <= 0; end_W(9, 319) <= 0; 
end_W(9, 320) <= 0; end_W(9, 321) <= 0; end_W(9, 322) <= 0; end_W(9, 323) <= 0; end_W(10, 0) <= 1; end_W(10, 1) <= 1; end_W(10, 2) <= 1; end_W(10, 3) <= 1; end_W(10, 4) <= 1; end_W(10, 5) <= 1; end_W(10, 6) <= 1; end_W(10, 7) <= 1; 
end_W(10, 8) <= 0; end_W(10, 9) <= 0; end_W(10, 10) <= 0; end_W(10, 11) <= 0; end_W(10, 12) <= 0; end_W(10, 13) <= 0; end_W(10, 14) <= 0; end_W(10, 15) <= 0; 
end_W(10, 16) <= 0; end_W(10, 17) <= 0; end_W(10, 18) <= 0; end_W(10, 19) <= 0; end_W(10, 20) <= 0; end_W(10, 21) <= 0; end_W(10, 22) <= 0; end_W(10, 23) <= 0; 
end_W(10, 24) <= 1; end_W(10, 25) <= 1; end_W(10, 26) <= 1; end_W(10, 27) <= 1; end_W(10, 28) <= 0; end_W(10, 29) <= 0; end_W(10, 30) <= 0; end_W(10, 31) <= 0; 
end_W(10, 32) <= 0; end_W(10, 33) <= 0; end_W(10, 34) <= 0; end_W(10, 35) <= 0; end_W(10, 36) <= 0; end_W(10, 37) <= 0; end_W(10, 38) <= 0; end_W(10, 39) <= 0; 
end_W(10, 40) <= 1; end_W(10, 41) <= 1; end_W(10, 42) <= 1; end_W(10, 43) <= 1; end_W(10, 44) <= 1; end_W(10, 45) <= 1; end_W(10, 46) <= 1; end_W(10, 47) <= 1; 
end_W(10, 48) <= 0; end_W(10, 49) <= 0; end_W(10, 50) <= 0; end_W(10, 51) <= 0; end_W(10, 52) <= 1; end_W(10, 53) <= 1; end_W(10, 54) <= 1; end_W(10, 55) <= 1; 
end_W(10, 56) <= 1; end_W(10, 57) <= 1; end_W(10, 58) <= 1; end_W(10, 59) <= 1; end_W(10, 60) <= 0; end_W(10, 61) <= 0; end_W(10, 62) <= 0; end_W(10, 63) <= 0; 
end_W(10, 64) <= 0; end_W(10, 65) <= 0; end_W(10, 66) <= 0; end_W(10, 67) <= 0; end_W(10, 68) <= 0; end_W(10, 69) <= 0; end_W(10, 70) <= 0; end_W(10, 71) <= 0; 
end_W(10, 72) <= 1; end_W(10, 73) <= 1; end_W(10, 74) <= 1; end_W(10, 75) <= 1; end_W(10, 76) <= 1; end_W(10, 77) <= 1; end_W(10, 78) <= 1; end_W(10, 79) <= 1; 
end_W(10, 80) <= 1; end_W(10, 81) <= 1; end_W(10, 82) <= 1; end_W(10, 83) <= 1; end_W(10, 84) <= 1; end_W(10, 85) <= 1; end_W(10, 86) <= 1; end_W(10, 87) <= 1; 
end_W(10, 88) <= 1; end_W(10, 89) <= 1; end_W(10, 90) <= 1; end_W(10, 91) <= 1; end_W(10, 92) <= 1; end_W(10, 93) <= 1; end_W(10, 94) <= 1; end_W(10, 95) <= 1; 
end_W(10, 96) <= 1; end_W(10, 97) <= 1; end_W(10, 98) <= 1; end_W(10, 99) <= 1; end_W(10, 100) <= 1; end_W(10, 101) <= 1; end_W(10, 102) <= 1; end_W(10, 103) <= 1; 
end_W(10, 104) <= 0; end_W(10, 105) <= 0; end_W(10, 106) <= 0; end_W(10, 107) <= 0; end_W(10, 108) <= 0; end_W(10, 109) <= 0; end_W(10, 110) <= 0; end_W(10, 111) <= 0; 
end_W(10, 112) <= 1; end_W(10, 113) <= 1; end_W(10, 114) <= 1; end_W(10, 115) <= 1; end_W(10, 116) <= 1; end_W(10, 117) <= 1; end_W(10, 118) <= 1; end_W(10, 119) <= 1; 
end_W(10, 120) <= 0; end_W(10, 121) <= 0; end_W(10, 122) <= 0; end_W(10, 123) <= 0; end_W(10, 124) <= 0; end_W(10, 125) <= 0; end_W(10, 126) <= 0; end_W(10, 127) <= 0; 
end_W(10, 128) <= 0; end_W(10, 129) <= 0; end_W(10, 130) <= 0; end_W(10, 131) <= 0; end_W(10, 132) <= 1; end_W(10, 133) <= 1; end_W(10, 134) <= 1; end_W(10, 135) <= 1; 
end_W(10, 136) <= 0; end_W(10, 137) <= 0; end_W(10, 138) <= 0; end_W(10, 139) <= 0; end_W(10, 140) <= 0; end_W(10, 141) <= 0; end_W(10, 142) <= 0; end_W(10, 143) <= 0; 
end_W(10, 144) <= 0; end_W(10, 145) <= 0; end_W(10, 146) <= 0; end_W(10, 147) <= 0; end_W(10, 148) <= 0; end_W(10, 149) <= 0; end_W(10, 150) <= 0; end_W(10, 151) <= 0; 
end_W(10, 152) <= 0; end_W(10, 153) <= 0; end_W(10, 154) <= 0; end_W(10, 155) <= 0; end_W(10, 156) <= 0; end_W(10, 157) <= 0; end_W(10, 158) <= 0; end_W(10, 159) <= 0; 
end_W(10, 160) <= 0; end_W(10, 161) <= 0; end_W(10, 162) <= 0; end_W(10, 163) <= 0; end_W(10, 164) <= 0; end_W(10, 165) <= 0; end_W(10, 166) <= 0; end_W(10, 167) <= 0; 
end_W(10, 168) <= 0; end_W(10, 169) <= 0; end_W(10, 170) <= 0; end_W(10, 171) <= 0; end_W(10, 172) <= 0; end_W(10, 173) <= 0; end_W(10, 174) <= 0; end_W(10, 175) <= 0; 
end_W(10, 176) <= 0; end_W(10, 177) <= 0; end_W(10, 178) <= 0; end_W(10, 179) <= 0; end_W(10, 180) <= 1; end_W(10, 181) <= 1; end_W(10, 182) <= 1; end_W(10, 183) <= 1; 
end_W(10, 184) <= 1; end_W(10, 185) <= 1; end_W(10, 186) <= 1; end_W(10, 187) <= 1; end_W(10, 188) <= 0; end_W(10, 189) <= 0; end_W(10, 190) <= 0; end_W(10, 191) <= 0; 
end_W(10, 192) <= 0; end_W(10, 193) <= 0; end_W(10, 194) <= 0; end_W(10, 195) <= 0; end_W(10, 196) <= 0; end_W(10, 197) <= 0; end_W(10, 198) <= 0; end_W(10, 199) <= 0; 
end_W(10, 200) <= 1; end_W(10, 201) <= 1; end_W(10, 202) <= 1; end_W(10, 203) <= 1; end_W(10, 204) <= 1; end_W(10, 205) <= 1; end_W(10, 206) <= 1; end_W(10, 207) <= 1; 
end_W(10, 208) <= 0; end_W(10, 209) <= 0; end_W(10, 210) <= 0; end_W(10, 211) <= 0; end_W(10, 212) <= 0; end_W(10, 213) <= 0; end_W(10, 214) <= 0; end_W(10, 215) <= 0; 
end_W(10, 216) <= 1; end_W(10, 217) <= 1; end_W(10, 218) <= 1; end_W(10, 219) <= 1; end_W(10, 220) <= 1; end_W(10, 221) <= 1; end_W(10, 222) <= 1; end_W(10, 223) <= 1; 
end_W(10, 224) <= 0; end_W(10, 225) <= 0; end_W(10, 226) <= 0; end_W(10, 227) <= 0; end_W(10, 228) <= 0; end_W(10, 229) <= 0; end_W(10, 230) <= 0; end_W(10, 231) <= 0; 
end_W(10, 232) <= 0; end_W(10, 233) <= 0; end_W(10, 234) <= 0; end_W(10, 235) <= 0; end_W(10, 236) <= 0; end_W(10, 237) <= 0; end_W(10, 238) <= 0; end_W(10, 239) <= 0; 
end_W(10, 240) <= 1; end_W(10, 241) <= 1; end_W(10, 242) <= 1; end_W(10, 243) <= 1; end_W(10, 244) <= 1; end_W(10, 245) <= 1; end_W(10, 246) <= 1; end_W(10, 247) <= 1; 
end_W(10, 248) <= 0; end_W(10, 249) <= 0; end_W(10, 250) <= 0; end_W(10, 251) <= 0; end_W(10, 252) <= 0; end_W(10, 253) <= 0; end_W(10, 254) <= 0; end_W(10, 255) <= 0; 
end_W(10, 256) <= 1; end_W(10, 257) <= 1; end_W(10, 258) <= 1; end_W(10, 259) <= 1; end_W(10, 260) <= 1; end_W(10, 261) <= 1; end_W(10, 262) <= 1; end_W(10, 263) <= 1; 
end_W(10, 264) <= 0; end_W(10, 265) <= 0; end_W(10, 266) <= 0; end_W(10, 267) <= 0; end_W(10, 268) <= 0; end_W(10, 269) <= 0; end_W(10, 270) <= 0; end_W(10, 271) <= 0; 
end_W(10, 272) <= 0; end_W(10, 273) <= 0; end_W(10, 274) <= 0; end_W(10, 275) <= 0; end_W(10, 276) <= 1; end_W(10, 277) <= 1; end_W(10, 278) <= 1; end_W(10, 279) <= 1; 
end_W(10, 280) <= 0; end_W(10, 281) <= 0; end_W(10, 282) <= 0; end_W(10, 283) <= 0; end_W(10, 284) <= 0; end_W(10, 285) <= 0; end_W(10, 286) <= 0; end_W(10, 287) <= 0; 
end_W(10, 288) <= 0; end_W(10, 289) <= 0; end_W(10, 290) <= 0; end_W(10, 291) <= 0; end_W(10, 292) <= 1; end_W(10, 293) <= 1; end_W(10, 294) <= 1; end_W(10, 295) <= 1; 
end_W(10, 296) <= 1; end_W(10, 297) <= 1; end_W(10, 298) <= 1; end_W(10, 299) <= 1; end_W(10, 300) <= 0; end_W(10, 301) <= 0; end_W(10, 302) <= 0; end_W(10, 303) <= 0; 
end_W(10, 304) <= 0; end_W(10, 305) <= 0; end_W(10, 306) <= 0; end_W(10, 307) <= 0; end_W(10, 308) <= 1; end_W(10, 309) <= 1; end_W(10, 310) <= 1; end_W(10, 311) <= 1; 
end_W(10, 312) <= 1; end_W(10, 313) <= 1; end_W(10, 314) <= 1; end_W(10, 315) <= 1; end_W(10, 316) <= 0; end_W(10, 317) <= 0; end_W(10, 318) <= 0; end_W(10, 319) <= 0; 
end_W(10, 320) <= 0; end_W(10, 321) <= 0; end_W(10, 322) <= 0; end_W(10, 323) <= 0; end_W(11, 0) <= 1; end_W(11, 1) <= 1; end_W(11, 2) <= 1; end_W(11, 3) <= 1; end_W(11, 4) <= 1; end_W(11, 5) <= 1; end_W(11, 6) <= 1; end_W(11, 7) <= 1; 
end_W(11, 8) <= 0; end_W(11, 9) <= 0; end_W(11, 10) <= 0; end_W(11, 11) <= 0; end_W(11, 12) <= 0; end_W(11, 13) <= 0; end_W(11, 14) <= 0; end_W(11, 15) <= 0; 
end_W(11, 16) <= 0; end_W(11, 17) <= 0; end_W(11, 18) <= 0; end_W(11, 19) <= 0; end_W(11, 20) <= 0; end_W(11, 21) <= 0; end_W(11, 22) <= 0; end_W(11, 23) <= 0; 
end_W(11, 24) <= 1; end_W(11, 25) <= 1; end_W(11, 26) <= 1; end_W(11, 27) <= 1; end_W(11, 28) <= 0; end_W(11, 29) <= 0; end_W(11, 30) <= 0; end_W(11, 31) <= 0; 
end_W(11, 32) <= 0; end_W(11, 33) <= 0; end_W(11, 34) <= 0; end_W(11, 35) <= 0; end_W(11, 36) <= 0; end_W(11, 37) <= 0; end_W(11, 38) <= 0; end_W(11, 39) <= 0; 
end_W(11, 40) <= 1; end_W(11, 41) <= 1; end_W(11, 42) <= 1; end_W(11, 43) <= 1; end_W(11, 44) <= 1; end_W(11, 45) <= 1; end_W(11, 46) <= 1; end_W(11, 47) <= 1; 
end_W(11, 48) <= 0; end_W(11, 49) <= 0; end_W(11, 50) <= 0; end_W(11, 51) <= 0; end_W(11, 52) <= 1; end_W(11, 53) <= 1; end_W(11, 54) <= 1; end_W(11, 55) <= 1; 
end_W(11, 56) <= 1; end_W(11, 57) <= 1; end_W(11, 58) <= 1; end_W(11, 59) <= 1; end_W(11, 60) <= 0; end_W(11, 61) <= 0; end_W(11, 62) <= 0; end_W(11, 63) <= 0; 
end_W(11, 64) <= 0; end_W(11, 65) <= 0; end_W(11, 66) <= 0; end_W(11, 67) <= 0; end_W(11, 68) <= 0; end_W(11, 69) <= 0; end_W(11, 70) <= 0; end_W(11, 71) <= 0; 
end_W(11, 72) <= 1; end_W(11, 73) <= 1; end_W(11, 74) <= 1; end_W(11, 75) <= 1; end_W(11, 76) <= 1; end_W(11, 77) <= 1; end_W(11, 78) <= 1; end_W(11, 79) <= 1; 
end_W(11, 80) <= 1; end_W(11, 81) <= 1; end_W(11, 82) <= 1; end_W(11, 83) <= 1; end_W(11, 84) <= 1; end_W(11, 85) <= 1; end_W(11, 86) <= 1; end_W(11, 87) <= 1; 
end_W(11, 88) <= 1; end_W(11, 89) <= 1; end_W(11, 90) <= 1; end_W(11, 91) <= 1; end_W(11, 92) <= 1; end_W(11, 93) <= 1; end_W(11, 94) <= 1; end_W(11, 95) <= 1; 
end_W(11, 96) <= 1; end_W(11, 97) <= 1; end_W(11, 98) <= 1; end_W(11, 99) <= 1; end_W(11, 100) <= 1; end_W(11, 101) <= 1; end_W(11, 102) <= 1; end_W(11, 103) <= 1; 
end_W(11, 104) <= 0; end_W(11, 105) <= 0; end_W(11, 106) <= 0; end_W(11, 107) <= 0; end_W(11, 108) <= 0; end_W(11, 109) <= 0; end_W(11, 110) <= 0; end_W(11, 111) <= 0; 
end_W(11, 112) <= 1; end_W(11, 113) <= 1; end_W(11, 114) <= 1; end_W(11, 115) <= 1; end_W(11, 116) <= 1; end_W(11, 117) <= 1; end_W(11, 118) <= 1; end_W(11, 119) <= 1; 
end_W(11, 120) <= 0; end_W(11, 121) <= 0; end_W(11, 122) <= 0; end_W(11, 123) <= 0; end_W(11, 124) <= 0; end_W(11, 125) <= 0; end_W(11, 126) <= 0; end_W(11, 127) <= 0; 
end_W(11, 128) <= 0; end_W(11, 129) <= 0; end_W(11, 130) <= 0; end_W(11, 131) <= 0; end_W(11, 132) <= 1; end_W(11, 133) <= 1; end_W(11, 134) <= 1; end_W(11, 135) <= 1; 
end_W(11, 136) <= 0; end_W(11, 137) <= 0; end_W(11, 138) <= 0; end_W(11, 139) <= 0; end_W(11, 140) <= 0; end_W(11, 141) <= 0; end_W(11, 142) <= 0; end_W(11, 143) <= 0; 
end_W(11, 144) <= 0; end_W(11, 145) <= 0; end_W(11, 146) <= 0; end_W(11, 147) <= 0; end_W(11, 148) <= 0; end_W(11, 149) <= 0; end_W(11, 150) <= 0; end_W(11, 151) <= 0; 
end_W(11, 152) <= 0; end_W(11, 153) <= 0; end_W(11, 154) <= 0; end_W(11, 155) <= 0; end_W(11, 156) <= 0; end_W(11, 157) <= 0; end_W(11, 158) <= 0; end_W(11, 159) <= 0; 
end_W(11, 160) <= 0; end_W(11, 161) <= 0; end_W(11, 162) <= 0; end_W(11, 163) <= 0; end_W(11, 164) <= 0; end_W(11, 165) <= 0; end_W(11, 166) <= 0; end_W(11, 167) <= 0; 
end_W(11, 168) <= 0; end_W(11, 169) <= 0; end_W(11, 170) <= 0; end_W(11, 171) <= 0; end_W(11, 172) <= 0; end_W(11, 173) <= 0; end_W(11, 174) <= 0; end_W(11, 175) <= 0; 
end_W(11, 176) <= 0; end_W(11, 177) <= 0; end_W(11, 178) <= 0; end_W(11, 179) <= 0; end_W(11, 180) <= 1; end_W(11, 181) <= 1; end_W(11, 182) <= 1; end_W(11, 183) <= 1; 
end_W(11, 184) <= 1; end_W(11, 185) <= 1; end_W(11, 186) <= 1; end_W(11, 187) <= 1; end_W(11, 188) <= 0; end_W(11, 189) <= 0; end_W(11, 190) <= 0; end_W(11, 191) <= 0; 
end_W(11, 192) <= 0; end_W(11, 193) <= 0; end_W(11, 194) <= 0; end_W(11, 195) <= 0; end_W(11, 196) <= 0; end_W(11, 197) <= 0; end_W(11, 198) <= 0; end_W(11, 199) <= 0; 
end_W(11, 200) <= 1; end_W(11, 201) <= 1; end_W(11, 202) <= 1; end_W(11, 203) <= 1; end_W(11, 204) <= 1; end_W(11, 205) <= 1; end_W(11, 206) <= 1; end_W(11, 207) <= 1; 
end_W(11, 208) <= 0; end_W(11, 209) <= 0; end_W(11, 210) <= 0; end_W(11, 211) <= 0; end_W(11, 212) <= 0; end_W(11, 213) <= 0; end_W(11, 214) <= 0; end_W(11, 215) <= 0; 
end_W(11, 216) <= 1; end_W(11, 217) <= 1; end_W(11, 218) <= 1; end_W(11, 219) <= 1; end_W(11, 220) <= 1; end_W(11, 221) <= 1; end_W(11, 222) <= 1; end_W(11, 223) <= 1; 
end_W(11, 224) <= 0; end_W(11, 225) <= 0; end_W(11, 226) <= 0; end_W(11, 227) <= 0; end_W(11, 228) <= 0; end_W(11, 229) <= 0; end_W(11, 230) <= 0; end_W(11, 231) <= 0; 
end_W(11, 232) <= 0; end_W(11, 233) <= 0; end_W(11, 234) <= 0; end_W(11, 235) <= 0; end_W(11, 236) <= 0; end_W(11, 237) <= 0; end_W(11, 238) <= 0; end_W(11, 239) <= 0; 
end_W(11, 240) <= 1; end_W(11, 241) <= 1; end_W(11, 242) <= 1; end_W(11, 243) <= 1; end_W(11, 244) <= 1; end_W(11, 245) <= 1; end_W(11, 246) <= 1; end_W(11, 247) <= 1; 
end_W(11, 248) <= 0; end_W(11, 249) <= 0; end_W(11, 250) <= 0; end_W(11, 251) <= 0; end_W(11, 252) <= 0; end_W(11, 253) <= 0; end_W(11, 254) <= 0; end_W(11, 255) <= 0; 
end_W(11, 256) <= 1; end_W(11, 257) <= 1; end_W(11, 258) <= 1; end_W(11, 259) <= 1; end_W(11, 260) <= 1; end_W(11, 261) <= 1; end_W(11, 262) <= 1; end_W(11, 263) <= 1; 
end_W(11, 264) <= 0; end_W(11, 265) <= 0; end_W(11, 266) <= 0; end_W(11, 267) <= 0; end_W(11, 268) <= 0; end_W(11, 269) <= 0; end_W(11, 270) <= 0; end_W(11, 271) <= 0; 
end_W(11, 272) <= 0; end_W(11, 273) <= 0; end_W(11, 274) <= 0; end_W(11, 275) <= 0; end_W(11, 276) <= 1; end_W(11, 277) <= 1; end_W(11, 278) <= 1; end_W(11, 279) <= 1; 
end_W(11, 280) <= 0; end_W(11, 281) <= 0; end_W(11, 282) <= 0; end_W(11, 283) <= 0; end_W(11, 284) <= 0; end_W(11, 285) <= 0; end_W(11, 286) <= 0; end_W(11, 287) <= 0; 
end_W(11, 288) <= 0; end_W(11, 289) <= 0; end_W(11, 290) <= 0; end_W(11, 291) <= 0; end_W(11, 292) <= 1; end_W(11, 293) <= 1; end_W(11, 294) <= 1; end_W(11, 295) <= 1; 
end_W(11, 296) <= 1; end_W(11, 297) <= 1; end_W(11, 298) <= 1; end_W(11, 299) <= 1; end_W(11, 300) <= 0; end_W(11, 301) <= 0; end_W(11, 302) <= 0; end_W(11, 303) <= 0; 
end_W(11, 304) <= 0; end_W(11, 305) <= 0; end_W(11, 306) <= 0; end_W(11, 307) <= 0; end_W(11, 308) <= 1; end_W(11, 309) <= 1; end_W(11, 310) <= 1; end_W(11, 311) <= 1; 
end_W(11, 312) <= 1; end_W(11, 313) <= 1; end_W(11, 314) <= 1; end_W(11, 315) <= 1; end_W(11, 316) <= 0; end_W(11, 317) <= 0; end_W(11, 318) <= 0; end_W(11, 319) <= 0; 
end_W(11, 320) <= 0; end_W(11, 321) <= 0; end_W(11, 322) <= 0; end_W(11, 323) <= 0; end_W(12, 0) <= 1; end_W(12, 1) <= 1; end_W(12, 2) <= 1; end_W(12, 3) <= 1; end_W(12, 4) <= 1; end_W(12, 5) <= 1; end_W(12, 6) <= 1; end_W(12, 7) <= 1; 
end_W(12, 8) <= 0; end_W(12, 9) <= 0; end_W(12, 10) <= 0; end_W(12, 11) <= 0; end_W(12, 12) <= 0; end_W(12, 13) <= 0; end_W(12, 14) <= 0; end_W(12, 15) <= 0; 
end_W(12, 16) <= 0; end_W(12, 17) <= 0; end_W(12, 18) <= 0; end_W(12, 19) <= 0; end_W(12, 20) <= 0; end_W(12, 21) <= 0; end_W(12, 22) <= 0; end_W(12, 23) <= 0; 
end_W(12, 24) <= 0; end_W(12, 25) <= 0; end_W(12, 26) <= 0; end_W(12, 27) <= 0; end_W(12, 28) <= 0; end_W(12, 29) <= 0; end_W(12, 30) <= 0; end_W(12, 31) <= 0; 
end_W(12, 32) <= 0; end_W(12, 33) <= 0; end_W(12, 34) <= 0; end_W(12, 35) <= 0; end_W(12, 36) <= 1; end_W(12, 37) <= 1; end_W(12, 38) <= 1; end_W(12, 39) <= 1; 
end_W(12, 40) <= 1; end_W(12, 41) <= 1; end_W(12, 42) <= 1; end_W(12, 43) <= 1; end_W(12, 44) <= 0; end_W(12, 45) <= 0; end_W(12, 46) <= 0; end_W(12, 47) <= 0; 
end_W(12, 48) <= 0; end_W(12, 49) <= 0; end_W(12, 50) <= 0; end_W(12, 51) <= 0; end_W(12, 52) <= 0; end_W(12, 53) <= 0; end_W(12, 54) <= 0; end_W(12, 55) <= 0; 
end_W(12, 56) <= 1; end_W(12, 57) <= 1; end_W(12, 58) <= 1; end_W(12, 59) <= 1; end_W(12, 60) <= 1; end_W(12, 61) <= 1; end_W(12, 62) <= 1; end_W(12, 63) <= 1; 
end_W(12, 64) <= 0; end_W(12, 65) <= 0; end_W(12, 66) <= 0; end_W(12, 67) <= 0; end_W(12, 68) <= 0; end_W(12, 69) <= 0; end_W(12, 70) <= 0; end_W(12, 71) <= 0; 
end_W(12, 72) <= 1; end_W(12, 73) <= 1; end_W(12, 74) <= 1; end_W(12, 75) <= 1; end_W(12, 76) <= 1; end_W(12, 77) <= 1; end_W(12, 78) <= 1; end_W(12, 79) <= 1; 
end_W(12, 80) <= 1; end_W(12, 81) <= 1; end_W(12, 82) <= 1; end_W(12, 83) <= 1; end_W(12, 84) <= 1; end_W(12, 85) <= 1; end_W(12, 86) <= 1; end_W(12, 87) <= 1; 
end_W(12, 88) <= 1; end_W(12, 89) <= 1; end_W(12, 90) <= 1; end_W(12, 91) <= 1; end_W(12, 92) <= 1; end_W(12, 93) <= 1; end_W(12, 94) <= 1; end_W(12, 95) <= 1; 
end_W(12, 96) <= 1; end_W(12, 97) <= 1; end_W(12, 98) <= 1; end_W(12, 99) <= 1; end_W(12, 100) <= 1; end_W(12, 101) <= 1; end_W(12, 102) <= 1; end_W(12, 103) <= 1; 
end_W(12, 104) <= 0; end_W(12, 105) <= 0; end_W(12, 106) <= 0; end_W(12, 107) <= 0; end_W(12, 108) <= 0; end_W(12, 109) <= 0; end_W(12, 110) <= 0; end_W(12, 111) <= 0; 
end_W(12, 112) <= 1; end_W(12, 113) <= 1; end_W(12, 114) <= 1; end_W(12, 115) <= 1; end_W(12, 116) <= 1; end_W(12, 117) <= 1; end_W(12, 118) <= 1; end_W(12, 119) <= 1; 
end_W(12, 120) <= 0; end_W(12, 121) <= 0; end_W(12, 122) <= 0; end_W(12, 123) <= 0; end_W(12, 124) <= 1; end_W(12, 125) <= 1; end_W(12, 126) <= 1; end_W(12, 127) <= 1; 
end_W(12, 128) <= 0; end_W(12, 129) <= 0; end_W(12, 130) <= 0; end_W(12, 131) <= 0; end_W(12, 132) <= 0; end_W(12, 133) <= 0; end_W(12, 134) <= 0; end_W(12, 135) <= 0; 
end_W(12, 136) <= 0; end_W(12, 137) <= 0; end_W(12, 138) <= 0; end_W(12, 139) <= 0; end_W(12, 140) <= 0; end_W(12, 141) <= 0; end_W(12, 142) <= 0; end_W(12, 143) <= 0; 
end_W(12, 144) <= 0; end_W(12, 145) <= 0; end_W(12, 146) <= 0; end_W(12, 147) <= 0; end_W(12, 148) <= 0; end_W(12, 149) <= 0; end_W(12, 150) <= 0; end_W(12, 151) <= 0; 
end_W(12, 152) <= 0; end_W(12, 153) <= 0; end_W(12, 154) <= 0; end_W(12, 155) <= 0; end_W(12, 156) <= 0; end_W(12, 157) <= 0; end_W(12, 158) <= 0; end_W(12, 159) <= 0; 
end_W(12, 160) <= 0; end_W(12, 161) <= 0; end_W(12, 162) <= 0; end_W(12, 163) <= 0; end_W(12, 164) <= 0; end_W(12, 165) <= 0; end_W(12, 166) <= 0; end_W(12, 167) <= 0; 
end_W(12, 168) <= 0; end_W(12, 169) <= 0; end_W(12, 170) <= 0; end_W(12, 171) <= 0; end_W(12, 172) <= 0; end_W(12, 173) <= 0; end_W(12, 174) <= 0; end_W(12, 175) <= 0; 
end_W(12, 176) <= 0; end_W(12, 177) <= 0; end_W(12, 178) <= 0; end_W(12, 179) <= 0; end_W(12, 180) <= 1; end_W(12, 181) <= 1; end_W(12, 182) <= 1; end_W(12, 183) <= 1; 
end_W(12, 184) <= 1; end_W(12, 185) <= 1; end_W(12, 186) <= 1; end_W(12, 187) <= 1; end_W(12, 188) <= 0; end_W(12, 189) <= 0; end_W(12, 190) <= 0; end_W(12, 191) <= 0; 
end_W(12, 192) <= 0; end_W(12, 193) <= 0; end_W(12, 194) <= 0; end_W(12, 195) <= 0; end_W(12, 196) <= 0; end_W(12, 197) <= 0; end_W(12, 198) <= 0; end_W(12, 199) <= 0; 
end_W(12, 200) <= 1; end_W(12, 201) <= 1; end_W(12, 202) <= 1; end_W(12, 203) <= 1; end_W(12, 204) <= 1; end_W(12, 205) <= 1; end_W(12, 206) <= 1; end_W(12, 207) <= 1; 
end_W(12, 208) <= 0; end_W(12, 209) <= 0; end_W(12, 210) <= 0; end_W(12, 211) <= 0; end_W(12, 212) <= 0; end_W(12, 213) <= 0; end_W(12, 214) <= 0; end_W(12, 215) <= 0; 
end_W(12, 216) <= 1; end_W(12, 217) <= 1; end_W(12, 218) <= 1; end_W(12, 219) <= 1; end_W(12, 220) <= 1; end_W(12, 221) <= 1; end_W(12, 222) <= 1; end_W(12, 223) <= 1; 
end_W(12, 224) <= 0; end_W(12, 225) <= 0; end_W(12, 226) <= 0; end_W(12, 227) <= 0; end_W(12, 228) <= 0; end_W(12, 229) <= 0; end_W(12, 230) <= 0; end_W(12, 231) <= 0; 
end_W(12, 232) <= 0; end_W(12, 233) <= 0; end_W(12, 234) <= 0; end_W(12, 235) <= 0; end_W(12, 236) <= 0; end_W(12, 237) <= 0; end_W(12, 238) <= 0; end_W(12, 239) <= 0; 
end_W(12, 240) <= 1; end_W(12, 241) <= 1; end_W(12, 242) <= 1; end_W(12, 243) <= 1; end_W(12, 244) <= 1; end_W(12, 245) <= 1; end_W(12, 246) <= 1; end_W(12, 247) <= 1; 
end_W(12, 248) <= 0; end_W(12, 249) <= 0; end_W(12, 250) <= 0; end_W(12, 251) <= 0; end_W(12, 252) <= 0; end_W(12, 253) <= 0; end_W(12, 254) <= 0; end_W(12, 255) <= 0; 
end_W(12, 256) <= 1; end_W(12, 257) <= 1; end_W(12, 258) <= 1; end_W(12, 259) <= 1; end_W(12, 260) <= 1; end_W(12, 261) <= 1; end_W(12, 262) <= 1; end_W(12, 263) <= 1; 
end_W(12, 264) <= 0; end_W(12, 265) <= 0; end_W(12, 266) <= 0; end_W(12, 267) <= 0; end_W(12, 268) <= 1; end_W(12, 269) <= 1; end_W(12, 270) <= 1; end_W(12, 271) <= 1; 
end_W(12, 272) <= 0; end_W(12, 273) <= 0; end_W(12, 274) <= 0; end_W(12, 275) <= 0; end_W(12, 276) <= 0; end_W(12, 277) <= 0; end_W(12, 278) <= 0; end_W(12, 279) <= 0; 
end_W(12, 280) <= 0; end_W(12, 281) <= 0; end_W(12, 282) <= 0; end_W(12, 283) <= 0; end_W(12, 284) <= 0; end_W(12, 285) <= 0; end_W(12, 286) <= 0; end_W(12, 287) <= 0; 
end_W(12, 288) <= 0; end_W(12, 289) <= 0; end_W(12, 290) <= 0; end_W(12, 291) <= 0; end_W(12, 292) <= 1; end_W(12, 293) <= 1; end_W(12, 294) <= 1; end_W(12, 295) <= 1; 
end_W(12, 296) <= 1; end_W(12, 297) <= 1; end_W(12, 298) <= 1; end_W(12, 299) <= 1; end_W(12, 300) <= 0; end_W(12, 301) <= 0; end_W(12, 302) <= 0; end_W(12, 303) <= 0; 
end_W(12, 304) <= 0; end_W(12, 305) <= 0; end_W(12, 306) <= 0; end_W(12, 307) <= 0; end_W(12, 308) <= 1; end_W(12, 309) <= 1; end_W(12, 310) <= 1; end_W(12, 311) <= 1; 
end_W(12, 312) <= 1; end_W(12, 313) <= 1; end_W(12, 314) <= 1; end_W(12, 315) <= 1; end_W(12, 316) <= 0; end_W(12, 317) <= 0; end_W(12, 318) <= 0; end_W(12, 319) <= 0; 
end_W(12, 320) <= 0; end_W(12, 321) <= 0; end_W(12, 322) <= 0; end_W(12, 323) <= 0; end_W(13, 0) <= 1; end_W(13, 1) <= 1; end_W(13, 2) <= 1; end_W(13, 3) <= 1; end_W(13, 4) <= 1; end_W(13, 5) <= 1; end_W(13, 6) <= 1; end_W(13, 7) <= 1; 
end_W(13, 8) <= 0; end_W(13, 9) <= 0; end_W(13, 10) <= 0; end_W(13, 11) <= 0; end_W(13, 12) <= 0; end_W(13, 13) <= 0; end_W(13, 14) <= 0; end_W(13, 15) <= 0; 
end_W(13, 16) <= 0; end_W(13, 17) <= 0; end_W(13, 18) <= 0; end_W(13, 19) <= 0; end_W(13, 20) <= 0; end_W(13, 21) <= 0; end_W(13, 22) <= 0; end_W(13, 23) <= 0; 
end_W(13, 24) <= 0; end_W(13, 25) <= 0; end_W(13, 26) <= 0; end_W(13, 27) <= 0; end_W(13, 28) <= 0; end_W(13, 29) <= 0; end_W(13, 30) <= 0; end_W(13, 31) <= 0; 
end_W(13, 32) <= 0; end_W(13, 33) <= 0; end_W(13, 34) <= 0; end_W(13, 35) <= 0; end_W(13, 36) <= 1; end_W(13, 37) <= 1; end_W(13, 38) <= 1; end_W(13, 39) <= 1; 
end_W(13, 40) <= 1; end_W(13, 41) <= 1; end_W(13, 42) <= 1; end_W(13, 43) <= 1; end_W(13, 44) <= 0; end_W(13, 45) <= 0; end_W(13, 46) <= 0; end_W(13, 47) <= 0; 
end_W(13, 48) <= 0; end_W(13, 49) <= 0; end_W(13, 50) <= 0; end_W(13, 51) <= 0; end_W(13, 52) <= 0; end_W(13, 53) <= 0; end_W(13, 54) <= 0; end_W(13, 55) <= 0; 
end_W(13, 56) <= 1; end_W(13, 57) <= 1; end_W(13, 58) <= 1; end_W(13, 59) <= 1; end_W(13, 60) <= 1; end_W(13, 61) <= 1; end_W(13, 62) <= 1; end_W(13, 63) <= 1; 
end_W(13, 64) <= 0; end_W(13, 65) <= 0; end_W(13, 66) <= 0; end_W(13, 67) <= 0; end_W(13, 68) <= 0; end_W(13, 69) <= 0; end_W(13, 70) <= 0; end_W(13, 71) <= 0; 
end_W(13, 72) <= 1; end_W(13, 73) <= 1; end_W(13, 74) <= 1; end_W(13, 75) <= 1; end_W(13, 76) <= 1; end_W(13, 77) <= 1; end_W(13, 78) <= 1; end_W(13, 79) <= 1; 
end_W(13, 80) <= 1; end_W(13, 81) <= 1; end_W(13, 82) <= 1; end_W(13, 83) <= 1; end_W(13, 84) <= 1; end_W(13, 85) <= 1; end_W(13, 86) <= 1; end_W(13, 87) <= 1; 
end_W(13, 88) <= 1; end_W(13, 89) <= 1; end_W(13, 90) <= 1; end_W(13, 91) <= 1; end_W(13, 92) <= 1; end_W(13, 93) <= 1; end_W(13, 94) <= 1; end_W(13, 95) <= 1; 
end_W(13, 96) <= 1; end_W(13, 97) <= 1; end_W(13, 98) <= 1; end_W(13, 99) <= 1; end_W(13, 100) <= 1; end_W(13, 101) <= 1; end_W(13, 102) <= 1; end_W(13, 103) <= 1; 
end_W(13, 104) <= 0; end_W(13, 105) <= 0; end_W(13, 106) <= 0; end_W(13, 107) <= 0; end_W(13, 108) <= 0; end_W(13, 109) <= 0; end_W(13, 110) <= 0; end_W(13, 111) <= 0; 
end_W(13, 112) <= 1; end_W(13, 113) <= 1; end_W(13, 114) <= 1; end_W(13, 115) <= 1; end_W(13, 116) <= 1; end_W(13, 117) <= 1; end_W(13, 118) <= 1; end_W(13, 119) <= 1; 
end_W(13, 120) <= 0; end_W(13, 121) <= 0; end_W(13, 122) <= 0; end_W(13, 123) <= 0; end_W(13, 124) <= 1; end_W(13, 125) <= 1; end_W(13, 126) <= 1; end_W(13, 127) <= 1; 
end_W(13, 128) <= 0; end_W(13, 129) <= 0; end_W(13, 130) <= 0; end_W(13, 131) <= 0; end_W(13, 132) <= 0; end_W(13, 133) <= 0; end_W(13, 134) <= 0; end_W(13, 135) <= 0; 
end_W(13, 136) <= 0; end_W(13, 137) <= 0; end_W(13, 138) <= 0; end_W(13, 139) <= 0; end_W(13, 140) <= 0; end_W(13, 141) <= 0; end_W(13, 142) <= 0; end_W(13, 143) <= 0; 
end_W(13, 144) <= 0; end_W(13, 145) <= 0; end_W(13, 146) <= 0; end_W(13, 147) <= 0; end_W(13, 148) <= 0; end_W(13, 149) <= 0; end_W(13, 150) <= 0; end_W(13, 151) <= 0; 
end_W(13, 152) <= 0; end_W(13, 153) <= 0; end_W(13, 154) <= 0; end_W(13, 155) <= 0; end_W(13, 156) <= 0; end_W(13, 157) <= 0; end_W(13, 158) <= 0; end_W(13, 159) <= 0; 
end_W(13, 160) <= 0; end_W(13, 161) <= 0; end_W(13, 162) <= 0; end_W(13, 163) <= 0; end_W(13, 164) <= 0; end_W(13, 165) <= 0; end_W(13, 166) <= 0; end_W(13, 167) <= 0; 
end_W(13, 168) <= 0; end_W(13, 169) <= 0; end_W(13, 170) <= 0; end_W(13, 171) <= 0; end_W(13, 172) <= 0; end_W(13, 173) <= 0; end_W(13, 174) <= 0; end_W(13, 175) <= 0; 
end_W(13, 176) <= 0; end_W(13, 177) <= 0; end_W(13, 178) <= 0; end_W(13, 179) <= 0; end_W(13, 180) <= 1; end_W(13, 181) <= 1; end_W(13, 182) <= 1; end_W(13, 183) <= 1; 
end_W(13, 184) <= 1; end_W(13, 185) <= 1; end_W(13, 186) <= 1; end_W(13, 187) <= 1; end_W(13, 188) <= 0; end_W(13, 189) <= 0; end_W(13, 190) <= 0; end_W(13, 191) <= 0; 
end_W(13, 192) <= 0; end_W(13, 193) <= 0; end_W(13, 194) <= 0; end_W(13, 195) <= 0; end_W(13, 196) <= 0; end_W(13, 197) <= 0; end_W(13, 198) <= 0; end_W(13, 199) <= 0; 
end_W(13, 200) <= 1; end_W(13, 201) <= 1; end_W(13, 202) <= 1; end_W(13, 203) <= 1; end_W(13, 204) <= 1; end_W(13, 205) <= 1; end_W(13, 206) <= 1; end_W(13, 207) <= 1; 
end_W(13, 208) <= 0; end_W(13, 209) <= 0; end_W(13, 210) <= 0; end_W(13, 211) <= 0; end_W(13, 212) <= 0; end_W(13, 213) <= 0; end_W(13, 214) <= 0; end_W(13, 215) <= 0; 
end_W(13, 216) <= 1; end_W(13, 217) <= 1; end_W(13, 218) <= 1; end_W(13, 219) <= 1; end_W(13, 220) <= 1; end_W(13, 221) <= 1; end_W(13, 222) <= 1; end_W(13, 223) <= 1; 
end_W(13, 224) <= 0; end_W(13, 225) <= 0; end_W(13, 226) <= 0; end_W(13, 227) <= 0; end_W(13, 228) <= 0; end_W(13, 229) <= 0; end_W(13, 230) <= 0; end_W(13, 231) <= 0; 
end_W(13, 232) <= 0; end_W(13, 233) <= 0; end_W(13, 234) <= 0; end_W(13, 235) <= 0; end_W(13, 236) <= 0; end_W(13, 237) <= 0; end_W(13, 238) <= 0; end_W(13, 239) <= 0; 
end_W(13, 240) <= 1; end_W(13, 241) <= 1; end_W(13, 242) <= 1; end_W(13, 243) <= 1; end_W(13, 244) <= 1; end_W(13, 245) <= 1; end_W(13, 246) <= 1; end_W(13, 247) <= 1; 
end_W(13, 248) <= 0; end_W(13, 249) <= 0; end_W(13, 250) <= 0; end_W(13, 251) <= 0; end_W(13, 252) <= 0; end_W(13, 253) <= 0; end_W(13, 254) <= 0; end_W(13, 255) <= 0; 
end_W(13, 256) <= 1; end_W(13, 257) <= 1; end_W(13, 258) <= 1; end_W(13, 259) <= 1; end_W(13, 260) <= 1; end_W(13, 261) <= 1; end_W(13, 262) <= 1; end_W(13, 263) <= 1; 
end_W(13, 264) <= 0; end_W(13, 265) <= 0; end_W(13, 266) <= 0; end_W(13, 267) <= 0; end_W(13, 268) <= 1; end_W(13, 269) <= 1; end_W(13, 270) <= 1; end_W(13, 271) <= 1; 
end_W(13, 272) <= 0; end_W(13, 273) <= 0; end_W(13, 274) <= 0; end_W(13, 275) <= 0; end_W(13, 276) <= 0; end_W(13, 277) <= 0; end_W(13, 278) <= 0; end_W(13, 279) <= 0; 
end_W(13, 280) <= 0; end_W(13, 281) <= 0; end_W(13, 282) <= 0; end_W(13, 283) <= 0; end_W(13, 284) <= 0; end_W(13, 285) <= 0; end_W(13, 286) <= 0; end_W(13, 287) <= 0; 
end_W(13, 288) <= 0; end_W(13, 289) <= 0; end_W(13, 290) <= 0; end_W(13, 291) <= 0; end_W(13, 292) <= 1; end_W(13, 293) <= 1; end_W(13, 294) <= 1; end_W(13, 295) <= 1; 
end_W(13, 296) <= 1; end_W(13, 297) <= 1; end_W(13, 298) <= 1; end_W(13, 299) <= 1; end_W(13, 300) <= 0; end_W(13, 301) <= 0; end_W(13, 302) <= 0; end_W(13, 303) <= 0; 
end_W(13, 304) <= 0; end_W(13, 305) <= 0; end_W(13, 306) <= 0; end_W(13, 307) <= 0; end_W(13, 308) <= 1; end_W(13, 309) <= 1; end_W(13, 310) <= 1; end_W(13, 311) <= 1; 
end_W(13, 312) <= 1; end_W(13, 313) <= 1; end_W(13, 314) <= 1; end_W(13, 315) <= 1; end_W(13, 316) <= 0; end_W(13, 317) <= 0; end_W(13, 318) <= 0; end_W(13, 319) <= 0; 
end_W(13, 320) <= 0; end_W(13, 321) <= 0; end_W(13, 322) <= 0; end_W(13, 323) <= 0; end_W(14, 0) <= 1; end_W(14, 1) <= 1; end_W(14, 2) <= 1; end_W(14, 3) <= 1; end_W(14, 4) <= 1; end_W(14, 5) <= 1; end_W(14, 6) <= 1; end_W(14, 7) <= 1; 
end_W(14, 8) <= 0; end_W(14, 9) <= 0; end_W(14, 10) <= 0; end_W(14, 11) <= 0; end_W(14, 12) <= 0; end_W(14, 13) <= 0; end_W(14, 14) <= 0; end_W(14, 15) <= 0; 
end_W(14, 16) <= 0; end_W(14, 17) <= 0; end_W(14, 18) <= 0; end_W(14, 19) <= 0; end_W(14, 20) <= 0; end_W(14, 21) <= 0; end_W(14, 22) <= 0; end_W(14, 23) <= 0; 
end_W(14, 24) <= 0; end_W(14, 25) <= 0; end_W(14, 26) <= 0; end_W(14, 27) <= 0; end_W(14, 28) <= 0; end_W(14, 29) <= 0; end_W(14, 30) <= 0; end_W(14, 31) <= 0; 
end_W(14, 32) <= 0; end_W(14, 33) <= 0; end_W(14, 34) <= 0; end_W(14, 35) <= 0; end_W(14, 36) <= 1; end_W(14, 37) <= 1; end_W(14, 38) <= 1; end_W(14, 39) <= 1; 
end_W(14, 40) <= 1; end_W(14, 41) <= 1; end_W(14, 42) <= 1; end_W(14, 43) <= 1; end_W(14, 44) <= 0; end_W(14, 45) <= 0; end_W(14, 46) <= 0; end_W(14, 47) <= 0; 
end_W(14, 48) <= 0; end_W(14, 49) <= 0; end_W(14, 50) <= 0; end_W(14, 51) <= 0; end_W(14, 52) <= 0; end_W(14, 53) <= 0; end_W(14, 54) <= 0; end_W(14, 55) <= 0; 
end_W(14, 56) <= 1; end_W(14, 57) <= 1; end_W(14, 58) <= 1; end_W(14, 59) <= 1; end_W(14, 60) <= 1; end_W(14, 61) <= 1; end_W(14, 62) <= 1; end_W(14, 63) <= 1; 
end_W(14, 64) <= 0; end_W(14, 65) <= 0; end_W(14, 66) <= 0; end_W(14, 67) <= 0; end_W(14, 68) <= 0; end_W(14, 69) <= 0; end_W(14, 70) <= 0; end_W(14, 71) <= 0; 
end_W(14, 72) <= 1; end_W(14, 73) <= 1; end_W(14, 74) <= 1; end_W(14, 75) <= 1; end_W(14, 76) <= 1; end_W(14, 77) <= 1; end_W(14, 78) <= 1; end_W(14, 79) <= 1; 
end_W(14, 80) <= 1; end_W(14, 81) <= 1; end_W(14, 82) <= 1; end_W(14, 83) <= 1; end_W(14, 84) <= 1; end_W(14, 85) <= 1; end_W(14, 86) <= 1; end_W(14, 87) <= 1; 
end_W(14, 88) <= 1; end_W(14, 89) <= 1; end_W(14, 90) <= 1; end_W(14, 91) <= 1; end_W(14, 92) <= 1; end_W(14, 93) <= 1; end_W(14, 94) <= 1; end_W(14, 95) <= 1; 
end_W(14, 96) <= 1; end_W(14, 97) <= 1; end_W(14, 98) <= 1; end_W(14, 99) <= 1; end_W(14, 100) <= 1; end_W(14, 101) <= 1; end_W(14, 102) <= 1; end_W(14, 103) <= 1; 
end_W(14, 104) <= 0; end_W(14, 105) <= 0; end_W(14, 106) <= 0; end_W(14, 107) <= 0; end_W(14, 108) <= 0; end_W(14, 109) <= 0; end_W(14, 110) <= 0; end_W(14, 111) <= 0; 
end_W(14, 112) <= 1; end_W(14, 113) <= 1; end_W(14, 114) <= 1; end_W(14, 115) <= 1; end_W(14, 116) <= 1; end_W(14, 117) <= 1; end_W(14, 118) <= 1; end_W(14, 119) <= 1; 
end_W(14, 120) <= 0; end_W(14, 121) <= 0; end_W(14, 122) <= 0; end_W(14, 123) <= 0; end_W(14, 124) <= 1; end_W(14, 125) <= 1; end_W(14, 126) <= 1; end_W(14, 127) <= 1; 
end_W(14, 128) <= 0; end_W(14, 129) <= 0; end_W(14, 130) <= 0; end_W(14, 131) <= 0; end_W(14, 132) <= 0; end_W(14, 133) <= 0; end_W(14, 134) <= 0; end_W(14, 135) <= 0; 
end_W(14, 136) <= 0; end_W(14, 137) <= 0; end_W(14, 138) <= 0; end_W(14, 139) <= 0; end_W(14, 140) <= 0; end_W(14, 141) <= 0; end_W(14, 142) <= 0; end_W(14, 143) <= 0; 
end_W(14, 144) <= 0; end_W(14, 145) <= 0; end_W(14, 146) <= 0; end_W(14, 147) <= 0; end_W(14, 148) <= 0; end_W(14, 149) <= 0; end_W(14, 150) <= 0; end_W(14, 151) <= 0; 
end_W(14, 152) <= 0; end_W(14, 153) <= 0; end_W(14, 154) <= 0; end_W(14, 155) <= 0; end_W(14, 156) <= 0; end_W(14, 157) <= 0; end_W(14, 158) <= 0; end_W(14, 159) <= 0; 
end_W(14, 160) <= 0; end_W(14, 161) <= 0; end_W(14, 162) <= 0; end_W(14, 163) <= 0; end_W(14, 164) <= 0; end_W(14, 165) <= 0; end_W(14, 166) <= 0; end_W(14, 167) <= 0; 
end_W(14, 168) <= 0; end_W(14, 169) <= 0; end_W(14, 170) <= 0; end_W(14, 171) <= 0; end_W(14, 172) <= 0; end_W(14, 173) <= 0; end_W(14, 174) <= 0; end_W(14, 175) <= 0; 
end_W(14, 176) <= 0; end_W(14, 177) <= 0; end_W(14, 178) <= 0; end_W(14, 179) <= 0; end_W(14, 180) <= 1; end_W(14, 181) <= 1; end_W(14, 182) <= 1; end_W(14, 183) <= 1; 
end_W(14, 184) <= 1; end_W(14, 185) <= 1; end_W(14, 186) <= 1; end_W(14, 187) <= 1; end_W(14, 188) <= 0; end_W(14, 189) <= 0; end_W(14, 190) <= 0; end_W(14, 191) <= 0; 
end_W(14, 192) <= 0; end_W(14, 193) <= 0; end_W(14, 194) <= 0; end_W(14, 195) <= 0; end_W(14, 196) <= 0; end_W(14, 197) <= 0; end_W(14, 198) <= 0; end_W(14, 199) <= 0; 
end_W(14, 200) <= 1; end_W(14, 201) <= 1; end_W(14, 202) <= 1; end_W(14, 203) <= 1; end_W(14, 204) <= 1; end_W(14, 205) <= 1; end_W(14, 206) <= 1; end_W(14, 207) <= 1; 
end_W(14, 208) <= 0; end_W(14, 209) <= 0; end_W(14, 210) <= 0; end_W(14, 211) <= 0; end_W(14, 212) <= 0; end_W(14, 213) <= 0; end_W(14, 214) <= 0; end_W(14, 215) <= 0; 
end_W(14, 216) <= 1; end_W(14, 217) <= 1; end_W(14, 218) <= 1; end_W(14, 219) <= 1; end_W(14, 220) <= 1; end_W(14, 221) <= 1; end_W(14, 222) <= 1; end_W(14, 223) <= 1; 
end_W(14, 224) <= 0; end_W(14, 225) <= 0; end_W(14, 226) <= 0; end_W(14, 227) <= 0; end_W(14, 228) <= 0; end_W(14, 229) <= 0; end_W(14, 230) <= 0; end_W(14, 231) <= 0; 
end_W(14, 232) <= 0; end_W(14, 233) <= 0; end_W(14, 234) <= 0; end_W(14, 235) <= 0; end_W(14, 236) <= 0; end_W(14, 237) <= 0; end_W(14, 238) <= 0; end_W(14, 239) <= 0; 
end_W(14, 240) <= 1; end_W(14, 241) <= 1; end_W(14, 242) <= 1; end_W(14, 243) <= 1; end_W(14, 244) <= 1; end_W(14, 245) <= 1; end_W(14, 246) <= 1; end_W(14, 247) <= 1; 
end_W(14, 248) <= 0; end_W(14, 249) <= 0; end_W(14, 250) <= 0; end_W(14, 251) <= 0; end_W(14, 252) <= 0; end_W(14, 253) <= 0; end_W(14, 254) <= 0; end_W(14, 255) <= 0; 
end_W(14, 256) <= 1; end_W(14, 257) <= 1; end_W(14, 258) <= 1; end_W(14, 259) <= 1; end_W(14, 260) <= 1; end_W(14, 261) <= 1; end_W(14, 262) <= 1; end_W(14, 263) <= 1; 
end_W(14, 264) <= 0; end_W(14, 265) <= 0; end_W(14, 266) <= 0; end_W(14, 267) <= 0; end_W(14, 268) <= 1; end_W(14, 269) <= 1; end_W(14, 270) <= 1; end_W(14, 271) <= 1; 
end_W(14, 272) <= 0; end_W(14, 273) <= 0; end_W(14, 274) <= 0; end_W(14, 275) <= 0; end_W(14, 276) <= 0; end_W(14, 277) <= 0; end_W(14, 278) <= 0; end_W(14, 279) <= 0; 
end_W(14, 280) <= 0; end_W(14, 281) <= 0; end_W(14, 282) <= 0; end_W(14, 283) <= 0; end_W(14, 284) <= 0; end_W(14, 285) <= 0; end_W(14, 286) <= 0; end_W(14, 287) <= 0; 
end_W(14, 288) <= 0; end_W(14, 289) <= 0; end_W(14, 290) <= 0; end_W(14, 291) <= 0; end_W(14, 292) <= 1; end_W(14, 293) <= 1; end_W(14, 294) <= 1; end_W(14, 295) <= 1; 
end_W(14, 296) <= 1; end_W(14, 297) <= 1; end_W(14, 298) <= 1; end_W(14, 299) <= 1; end_W(14, 300) <= 0; end_W(14, 301) <= 0; end_W(14, 302) <= 0; end_W(14, 303) <= 0; 
end_W(14, 304) <= 0; end_W(14, 305) <= 0; end_W(14, 306) <= 0; end_W(14, 307) <= 0; end_W(14, 308) <= 1; end_W(14, 309) <= 1; end_W(14, 310) <= 1; end_W(14, 311) <= 1; 
end_W(14, 312) <= 1; end_W(14, 313) <= 1; end_W(14, 314) <= 1; end_W(14, 315) <= 1; end_W(14, 316) <= 0; end_W(14, 317) <= 0; end_W(14, 318) <= 0; end_W(14, 319) <= 0; 
end_W(14, 320) <= 0; end_W(14, 321) <= 0; end_W(14, 322) <= 0; end_W(14, 323) <= 0; end_W(15, 0) <= 1; end_W(15, 1) <= 1; end_W(15, 2) <= 1; end_W(15, 3) <= 1; end_W(15, 4) <= 1; end_W(15, 5) <= 1; end_W(15, 6) <= 1; end_W(15, 7) <= 1; 
end_W(15, 8) <= 0; end_W(15, 9) <= 0; end_W(15, 10) <= 0; end_W(15, 11) <= 0; end_W(15, 12) <= 0; end_W(15, 13) <= 0; end_W(15, 14) <= 0; end_W(15, 15) <= 0; 
end_W(15, 16) <= 0; end_W(15, 17) <= 0; end_W(15, 18) <= 0; end_W(15, 19) <= 0; end_W(15, 20) <= 0; end_W(15, 21) <= 0; end_W(15, 22) <= 0; end_W(15, 23) <= 0; 
end_W(15, 24) <= 0; end_W(15, 25) <= 0; end_W(15, 26) <= 0; end_W(15, 27) <= 0; end_W(15, 28) <= 0; end_W(15, 29) <= 0; end_W(15, 30) <= 0; end_W(15, 31) <= 0; 
end_W(15, 32) <= 0; end_W(15, 33) <= 0; end_W(15, 34) <= 0; end_W(15, 35) <= 0; end_W(15, 36) <= 1; end_W(15, 37) <= 1; end_W(15, 38) <= 1; end_W(15, 39) <= 1; 
end_W(15, 40) <= 1; end_W(15, 41) <= 1; end_W(15, 42) <= 1; end_W(15, 43) <= 1; end_W(15, 44) <= 0; end_W(15, 45) <= 0; end_W(15, 46) <= 0; end_W(15, 47) <= 0; 
end_W(15, 48) <= 0; end_W(15, 49) <= 0; end_W(15, 50) <= 0; end_W(15, 51) <= 0; end_W(15, 52) <= 0; end_W(15, 53) <= 0; end_W(15, 54) <= 0; end_W(15, 55) <= 0; 
end_W(15, 56) <= 1; end_W(15, 57) <= 1; end_W(15, 58) <= 1; end_W(15, 59) <= 1; end_W(15, 60) <= 1; end_W(15, 61) <= 1; end_W(15, 62) <= 1; end_W(15, 63) <= 1; 
end_W(15, 64) <= 0; end_W(15, 65) <= 0; end_W(15, 66) <= 0; end_W(15, 67) <= 0; end_W(15, 68) <= 0; end_W(15, 69) <= 0; end_W(15, 70) <= 0; end_W(15, 71) <= 0; 
end_W(15, 72) <= 1; end_W(15, 73) <= 1; end_W(15, 74) <= 1; end_W(15, 75) <= 1; end_W(15, 76) <= 1; end_W(15, 77) <= 1; end_W(15, 78) <= 1; end_W(15, 79) <= 1; 
end_W(15, 80) <= 1; end_W(15, 81) <= 1; end_W(15, 82) <= 1; end_W(15, 83) <= 1; end_W(15, 84) <= 1; end_W(15, 85) <= 1; end_W(15, 86) <= 1; end_W(15, 87) <= 1; 
end_W(15, 88) <= 1; end_W(15, 89) <= 1; end_W(15, 90) <= 1; end_W(15, 91) <= 1; end_W(15, 92) <= 1; end_W(15, 93) <= 1; end_W(15, 94) <= 1; end_W(15, 95) <= 1; 
end_W(15, 96) <= 1; end_W(15, 97) <= 1; end_W(15, 98) <= 1; end_W(15, 99) <= 1; end_W(15, 100) <= 1; end_W(15, 101) <= 1; end_W(15, 102) <= 1; end_W(15, 103) <= 1; 
end_W(15, 104) <= 0; end_W(15, 105) <= 0; end_W(15, 106) <= 0; end_W(15, 107) <= 0; end_W(15, 108) <= 0; end_W(15, 109) <= 0; end_W(15, 110) <= 0; end_W(15, 111) <= 0; 
end_W(15, 112) <= 1; end_W(15, 113) <= 1; end_W(15, 114) <= 1; end_W(15, 115) <= 1; end_W(15, 116) <= 1; end_W(15, 117) <= 1; end_W(15, 118) <= 1; end_W(15, 119) <= 1; 
end_W(15, 120) <= 0; end_W(15, 121) <= 0; end_W(15, 122) <= 0; end_W(15, 123) <= 0; end_W(15, 124) <= 1; end_W(15, 125) <= 1; end_W(15, 126) <= 1; end_W(15, 127) <= 1; 
end_W(15, 128) <= 0; end_W(15, 129) <= 0; end_W(15, 130) <= 0; end_W(15, 131) <= 0; end_W(15, 132) <= 0; end_W(15, 133) <= 0; end_W(15, 134) <= 0; end_W(15, 135) <= 0; 
end_W(15, 136) <= 0; end_W(15, 137) <= 0; end_W(15, 138) <= 0; end_W(15, 139) <= 0; end_W(15, 140) <= 0; end_W(15, 141) <= 0; end_W(15, 142) <= 0; end_W(15, 143) <= 0; 
end_W(15, 144) <= 0; end_W(15, 145) <= 0; end_W(15, 146) <= 0; end_W(15, 147) <= 0; end_W(15, 148) <= 0; end_W(15, 149) <= 0; end_W(15, 150) <= 0; end_W(15, 151) <= 0; 
end_W(15, 152) <= 0; end_W(15, 153) <= 0; end_W(15, 154) <= 0; end_W(15, 155) <= 0; end_W(15, 156) <= 0; end_W(15, 157) <= 0; end_W(15, 158) <= 0; end_W(15, 159) <= 0; 
end_W(15, 160) <= 0; end_W(15, 161) <= 0; end_W(15, 162) <= 0; end_W(15, 163) <= 0; end_W(15, 164) <= 0; end_W(15, 165) <= 0; end_W(15, 166) <= 0; end_W(15, 167) <= 0; 
end_W(15, 168) <= 0; end_W(15, 169) <= 0; end_W(15, 170) <= 0; end_W(15, 171) <= 0; end_W(15, 172) <= 0; end_W(15, 173) <= 0; end_W(15, 174) <= 0; end_W(15, 175) <= 0; 
end_W(15, 176) <= 0; end_W(15, 177) <= 0; end_W(15, 178) <= 0; end_W(15, 179) <= 0; end_W(15, 180) <= 1; end_W(15, 181) <= 1; end_W(15, 182) <= 1; end_W(15, 183) <= 1; 
end_W(15, 184) <= 1; end_W(15, 185) <= 1; end_W(15, 186) <= 1; end_W(15, 187) <= 1; end_W(15, 188) <= 0; end_W(15, 189) <= 0; end_W(15, 190) <= 0; end_W(15, 191) <= 0; 
end_W(15, 192) <= 0; end_W(15, 193) <= 0; end_W(15, 194) <= 0; end_W(15, 195) <= 0; end_W(15, 196) <= 0; end_W(15, 197) <= 0; end_W(15, 198) <= 0; end_W(15, 199) <= 0; 
end_W(15, 200) <= 1; end_W(15, 201) <= 1; end_W(15, 202) <= 1; end_W(15, 203) <= 1; end_W(15, 204) <= 1; end_W(15, 205) <= 1; end_W(15, 206) <= 1; end_W(15, 207) <= 1; 
end_W(15, 208) <= 0; end_W(15, 209) <= 0; end_W(15, 210) <= 0; end_W(15, 211) <= 0; end_W(15, 212) <= 0; end_W(15, 213) <= 0; end_W(15, 214) <= 0; end_W(15, 215) <= 0; 
end_W(15, 216) <= 1; end_W(15, 217) <= 1; end_W(15, 218) <= 1; end_W(15, 219) <= 1; end_W(15, 220) <= 1; end_W(15, 221) <= 1; end_W(15, 222) <= 1; end_W(15, 223) <= 1; 
end_W(15, 224) <= 0; end_W(15, 225) <= 0; end_W(15, 226) <= 0; end_W(15, 227) <= 0; end_W(15, 228) <= 0; end_W(15, 229) <= 0; end_W(15, 230) <= 0; end_W(15, 231) <= 0; 
end_W(15, 232) <= 0; end_W(15, 233) <= 0; end_W(15, 234) <= 0; end_W(15, 235) <= 0; end_W(15, 236) <= 0; end_W(15, 237) <= 0; end_W(15, 238) <= 0; end_W(15, 239) <= 0; 
end_W(15, 240) <= 1; end_W(15, 241) <= 1; end_W(15, 242) <= 1; end_W(15, 243) <= 1; end_W(15, 244) <= 1; end_W(15, 245) <= 1; end_W(15, 246) <= 1; end_W(15, 247) <= 1; 
end_W(15, 248) <= 0; end_W(15, 249) <= 0; end_W(15, 250) <= 0; end_W(15, 251) <= 0; end_W(15, 252) <= 0; end_W(15, 253) <= 0; end_W(15, 254) <= 0; end_W(15, 255) <= 0; 
end_W(15, 256) <= 1; end_W(15, 257) <= 1; end_W(15, 258) <= 1; end_W(15, 259) <= 1; end_W(15, 260) <= 1; end_W(15, 261) <= 1; end_W(15, 262) <= 1; end_W(15, 263) <= 1; 
end_W(15, 264) <= 0; end_W(15, 265) <= 0; end_W(15, 266) <= 0; end_W(15, 267) <= 0; end_W(15, 268) <= 1; end_W(15, 269) <= 1; end_W(15, 270) <= 1; end_W(15, 271) <= 1; 
end_W(15, 272) <= 0; end_W(15, 273) <= 0; end_W(15, 274) <= 0; end_W(15, 275) <= 0; end_W(15, 276) <= 0; end_W(15, 277) <= 0; end_W(15, 278) <= 0; end_W(15, 279) <= 0; 
end_W(15, 280) <= 0; end_W(15, 281) <= 0; end_W(15, 282) <= 0; end_W(15, 283) <= 0; end_W(15, 284) <= 0; end_W(15, 285) <= 0; end_W(15, 286) <= 0; end_W(15, 287) <= 0; 
end_W(15, 288) <= 0; end_W(15, 289) <= 0; end_W(15, 290) <= 0; end_W(15, 291) <= 0; end_W(15, 292) <= 1; end_W(15, 293) <= 1; end_W(15, 294) <= 1; end_W(15, 295) <= 1; 
end_W(15, 296) <= 1; end_W(15, 297) <= 1; end_W(15, 298) <= 1; end_W(15, 299) <= 1; end_W(15, 300) <= 0; end_W(15, 301) <= 0; end_W(15, 302) <= 0; end_W(15, 303) <= 0; 
end_W(15, 304) <= 0; end_W(15, 305) <= 0; end_W(15, 306) <= 0; end_W(15, 307) <= 0; end_W(15, 308) <= 1; end_W(15, 309) <= 1; end_W(15, 310) <= 1; end_W(15, 311) <= 1; 
end_W(15, 312) <= 1; end_W(15, 313) <= 1; end_W(15, 314) <= 1; end_W(15, 315) <= 1; end_W(15, 316) <= 0; end_W(15, 317) <= 0; end_W(15, 318) <= 0; end_W(15, 319) <= 0; 
end_W(15, 320) <= 0; end_W(15, 321) <= 0; end_W(15, 322) <= 0; end_W(15, 323) <= 0; end_W(16, 0) <= 1; end_W(16, 1) <= 1; end_W(16, 2) <= 1; end_W(16, 3) <= 1; end_W(16, 4) <= 1; end_W(16, 5) <= 1; end_W(16, 6) <= 1; end_W(16, 7) <= 1; 
end_W(16, 8) <= 0; end_W(16, 9) <= 0; end_W(16, 10) <= 0; end_W(16, 11) <= 0; end_W(16, 12) <= 0; end_W(16, 13) <= 0; end_W(16, 14) <= 0; end_W(16, 15) <= 0; 
end_W(16, 16) <= 0; end_W(16, 17) <= 0; end_W(16, 18) <= 0; end_W(16, 19) <= 0; end_W(16, 20) <= 0; end_W(16, 21) <= 0; end_W(16, 22) <= 0; end_W(16, 23) <= 0; 
end_W(16, 24) <= 0; end_W(16, 25) <= 0; end_W(16, 26) <= 0; end_W(16, 27) <= 0; end_W(16, 28) <= 0; end_W(16, 29) <= 0; end_W(16, 30) <= 0; end_W(16, 31) <= 0; 
end_W(16, 32) <= 0; end_W(16, 33) <= 0; end_W(16, 34) <= 0; end_W(16, 35) <= 0; end_W(16, 36) <= 1; end_W(16, 37) <= 1; end_W(16, 38) <= 1; end_W(16, 39) <= 1; 
end_W(16, 40) <= 1; end_W(16, 41) <= 1; end_W(16, 42) <= 1; end_W(16, 43) <= 1; end_W(16, 44) <= 0; end_W(16, 45) <= 0; end_W(16, 46) <= 0; end_W(16, 47) <= 0; 
end_W(16, 48) <= 0; end_W(16, 49) <= 0; end_W(16, 50) <= 0; end_W(16, 51) <= 0; end_W(16, 52) <= 0; end_W(16, 53) <= 0; end_W(16, 54) <= 0; end_W(16, 55) <= 0; 
end_W(16, 56) <= 1; end_W(16, 57) <= 1; end_W(16, 58) <= 1; end_W(16, 59) <= 1; end_W(16, 60) <= 1; end_W(16, 61) <= 1; end_W(16, 62) <= 1; end_W(16, 63) <= 1; 
end_W(16, 64) <= 0; end_W(16, 65) <= 0; end_W(16, 66) <= 0; end_W(16, 67) <= 0; end_W(16, 68) <= 0; end_W(16, 69) <= 0; end_W(16, 70) <= 0; end_W(16, 71) <= 0; 
end_W(16, 72) <= 1; end_W(16, 73) <= 1; end_W(16, 74) <= 1; end_W(16, 75) <= 1; end_W(16, 76) <= 1; end_W(16, 77) <= 1; end_W(16, 78) <= 1; end_W(16, 79) <= 1; 
end_W(16, 80) <= 0; end_W(16, 81) <= 0; end_W(16, 82) <= 0; end_W(16, 83) <= 0; end_W(16, 84) <= 1; end_W(16, 85) <= 1; end_W(16, 86) <= 1; end_W(16, 87) <= 1; 
end_W(16, 88) <= 1; end_W(16, 89) <= 1; end_W(16, 90) <= 1; end_W(16, 91) <= 1; end_W(16, 92) <= 0; end_W(16, 93) <= 0; end_W(16, 94) <= 0; end_W(16, 95) <= 0; 
end_W(16, 96) <= 1; end_W(16, 97) <= 1; end_W(16, 98) <= 1; end_W(16, 99) <= 1; end_W(16, 100) <= 1; end_W(16, 101) <= 1; end_W(16, 102) <= 1; end_W(16, 103) <= 1; 
end_W(16, 104) <= 0; end_W(16, 105) <= 0; end_W(16, 106) <= 0; end_W(16, 107) <= 0; end_W(16, 108) <= 0; end_W(16, 109) <= 0; end_W(16, 110) <= 0; end_W(16, 111) <= 0; 
end_W(16, 112) <= 1; end_W(16, 113) <= 1; end_W(16, 114) <= 1; end_W(16, 115) <= 1; end_W(16, 116) <= 1; end_W(16, 117) <= 1; end_W(16, 118) <= 1; end_W(16, 119) <= 1; 
end_W(16, 120) <= 1; end_W(16, 121) <= 1; end_W(16, 122) <= 1; end_W(16, 123) <= 1; end_W(16, 124) <= 1; end_W(16, 125) <= 1; end_W(16, 126) <= 1; end_W(16, 127) <= 1; 
end_W(16, 128) <= 0; end_W(16, 129) <= 0; end_W(16, 130) <= 0; end_W(16, 131) <= 0; end_W(16, 132) <= 0; end_W(16, 133) <= 0; end_W(16, 134) <= 0; end_W(16, 135) <= 0; 
end_W(16, 136) <= 0; end_W(16, 137) <= 0; end_W(16, 138) <= 0; end_W(16, 139) <= 0; end_W(16, 140) <= 0; end_W(16, 141) <= 0; end_W(16, 142) <= 0; end_W(16, 143) <= 0; 
end_W(16, 144) <= 0; end_W(16, 145) <= 0; end_W(16, 146) <= 0; end_W(16, 147) <= 0; end_W(16, 148) <= 0; end_W(16, 149) <= 0; end_W(16, 150) <= 0; end_W(16, 151) <= 0; 
end_W(16, 152) <= 0; end_W(16, 153) <= 0; end_W(16, 154) <= 0; end_W(16, 155) <= 0; end_W(16, 156) <= 0; end_W(16, 157) <= 0; end_W(16, 158) <= 0; end_W(16, 159) <= 0; 
end_W(16, 160) <= 0; end_W(16, 161) <= 0; end_W(16, 162) <= 0; end_W(16, 163) <= 0; end_W(16, 164) <= 0; end_W(16, 165) <= 0; end_W(16, 166) <= 0; end_W(16, 167) <= 0; 
end_W(16, 168) <= 0; end_W(16, 169) <= 0; end_W(16, 170) <= 0; end_W(16, 171) <= 0; end_W(16, 172) <= 0; end_W(16, 173) <= 0; end_W(16, 174) <= 0; end_W(16, 175) <= 0; 
end_W(16, 176) <= 0; end_W(16, 177) <= 0; end_W(16, 178) <= 0; end_W(16, 179) <= 0; end_W(16, 180) <= 1; end_W(16, 181) <= 1; end_W(16, 182) <= 1; end_W(16, 183) <= 1; 
end_W(16, 184) <= 1; end_W(16, 185) <= 1; end_W(16, 186) <= 1; end_W(16, 187) <= 1; end_W(16, 188) <= 0; end_W(16, 189) <= 0; end_W(16, 190) <= 0; end_W(16, 191) <= 0; 
end_W(16, 192) <= 0; end_W(16, 193) <= 0; end_W(16, 194) <= 0; end_W(16, 195) <= 0; end_W(16, 196) <= 0; end_W(16, 197) <= 0; end_W(16, 198) <= 0; end_W(16, 199) <= 0; 
end_W(16, 200) <= 1; end_W(16, 201) <= 1; end_W(16, 202) <= 1; end_W(16, 203) <= 1; end_W(16, 204) <= 1; end_W(16, 205) <= 1; end_W(16, 206) <= 1; end_W(16, 207) <= 1; 
end_W(16, 208) <= 0; end_W(16, 209) <= 0; end_W(16, 210) <= 0; end_W(16, 211) <= 0; end_W(16, 212) <= 0; end_W(16, 213) <= 0; end_W(16, 214) <= 0; end_W(16, 215) <= 0; 
end_W(16, 216) <= 1; end_W(16, 217) <= 1; end_W(16, 218) <= 1; end_W(16, 219) <= 1; end_W(16, 220) <= 1; end_W(16, 221) <= 1; end_W(16, 222) <= 1; end_W(16, 223) <= 1; 
end_W(16, 224) <= 0; end_W(16, 225) <= 0; end_W(16, 226) <= 0; end_W(16, 227) <= 0; end_W(16, 228) <= 0; end_W(16, 229) <= 0; end_W(16, 230) <= 0; end_W(16, 231) <= 0; 
end_W(16, 232) <= 0; end_W(16, 233) <= 0; end_W(16, 234) <= 0; end_W(16, 235) <= 0; end_W(16, 236) <= 0; end_W(16, 237) <= 0; end_W(16, 238) <= 0; end_W(16, 239) <= 0; 
end_W(16, 240) <= 1; end_W(16, 241) <= 1; end_W(16, 242) <= 1; end_W(16, 243) <= 1; end_W(16, 244) <= 1; end_W(16, 245) <= 1; end_W(16, 246) <= 1; end_W(16, 247) <= 1; 
end_W(16, 248) <= 0; end_W(16, 249) <= 0; end_W(16, 250) <= 0; end_W(16, 251) <= 0; end_W(16, 252) <= 0; end_W(16, 253) <= 0; end_W(16, 254) <= 0; end_W(16, 255) <= 0; 
end_W(16, 256) <= 1; end_W(16, 257) <= 1; end_W(16, 258) <= 1; end_W(16, 259) <= 1; end_W(16, 260) <= 1; end_W(16, 261) <= 1; end_W(16, 262) <= 1; end_W(16, 263) <= 1; 
end_W(16, 264) <= 1; end_W(16, 265) <= 1; end_W(16, 266) <= 1; end_W(16, 267) <= 1; end_W(16, 268) <= 1; end_W(16, 269) <= 1; end_W(16, 270) <= 1; end_W(16, 271) <= 1; 
end_W(16, 272) <= 0; end_W(16, 273) <= 0; end_W(16, 274) <= 0; end_W(16, 275) <= 0; end_W(16, 276) <= 0; end_W(16, 277) <= 0; end_W(16, 278) <= 0; end_W(16, 279) <= 0; 
end_W(16, 280) <= 0; end_W(16, 281) <= 0; end_W(16, 282) <= 0; end_W(16, 283) <= 0; end_W(16, 284) <= 0; end_W(16, 285) <= 0; end_W(16, 286) <= 0; end_W(16, 287) <= 0; 
end_W(16, 288) <= 0; end_W(16, 289) <= 0; end_W(16, 290) <= 0; end_W(16, 291) <= 0; end_W(16, 292) <= 1; end_W(16, 293) <= 1; end_W(16, 294) <= 1; end_W(16, 295) <= 1; 
end_W(16, 296) <= 1; end_W(16, 297) <= 1; end_W(16, 298) <= 1; end_W(16, 299) <= 1; end_W(16, 300) <= 1; end_W(16, 301) <= 1; end_W(16, 302) <= 1; end_W(16, 303) <= 1; 
end_W(16, 304) <= 1; end_W(16, 305) <= 1; end_W(16, 306) <= 1; end_W(16, 307) <= 1; end_W(16, 308) <= 1; end_W(16, 309) <= 1; end_W(16, 310) <= 1; end_W(16, 311) <= 1; 
end_W(16, 312) <= 0; end_W(16, 313) <= 0; end_W(16, 314) <= 0; end_W(16, 315) <= 0; end_W(16, 316) <= 0; end_W(16, 317) <= 0; end_W(16, 318) <= 0; end_W(16, 319) <= 0; 
end_W(16, 320) <= 0; end_W(16, 321) <= 0; end_W(16, 322) <= 0; end_W(16, 323) <= 0; end_W(17, 0) <= 1; end_W(17, 1) <= 1; end_W(17, 2) <= 1; end_W(17, 3) <= 1; end_W(17, 4) <= 1; end_W(17, 5) <= 1; end_W(17, 6) <= 1; end_W(17, 7) <= 1; 
end_W(17, 8) <= 0; end_W(17, 9) <= 0; end_W(17, 10) <= 0; end_W(17, 11) <= 0; end_W(17, 12) <= 0; end_W(17, 13) <= 0; end_W(17, 14) <= 0; end_W(17, 15) <= 0; 
end_W(17, 16) <= 0; end_W(17, 17) <= 0; end_W(17, 18) <= 0; end_W(17, 19) <= 0; end_W(17, 20) <= 0; end_W(17, 21) <= 0; end_W(17, 22) <= 0; end_W(17, 23) <= 0; 
end_W(17, 24) <= 0; end_W(17, 25) <= 0; end_W(17, 26) <= 0; end_W(17, 27) <= 0; end_W(17, 28) <= 0; end_W(17, 29) <= 0; end_W(17, 30) <= 0; end_W(17, 31) <= 0; 
end_W(17, 32) <= 0; end_W(17, 33) <= 0; end_W(17, 34) <= 0; end_W(17, 35) <= 0; end_W(17, 36) <= 1; end_W(17, 37) <= 1; end_W(17, 38) <= 1; end_W(17, 39) <= 1; 
end_W(17, 40) <= 1; end_W(17, 41) <= 1; end_W(17, 42) <= 1; end_W(17, 43) <= 1; end_W(17, 44) <= 0; end_W(17, 45) <= 0; end_W(17, 46) <= 0; end_W(17, 47) <= 0; 
end_W(17, 48) <= 0; end_W(17, 49) <= 0; end_W(17, 50) <= 0; end_W(17, 51) <= 0; end_W(17, 52) <= 0; end_W(17, 53) <= 0; end_W(17, 54) <= 0; end_W(17, 55) <= 0; 
end_W(17, 56) <= 1; end_W(17, 57) <= 1; end_W(17, 58) <= 1; end_W(17, 59) <= 1; end_W(17, 60) <= 1; end_W(17, 61) <= 1; end_W(17, 62) <= 1; end_W(17, 63) <= 1; 
end_W(17, 64) <= 0; end_W(17, 65) <= 0; end_W(17, 66) <= 0; end_W(17, 67) <= 0; end_W(17, 68) <= 0; end_W(17, 69) <= 0; end_W(17, 70) <= 0; end_W(17, 71) <= 0; 
end_W(17, 72) <= 1; end_W(17, 73) <= 1; end_W(17, 74) <= 1; end_W(17, 75) <= 1; end_W(17, 76) <= 1; end_W(17, 77) <= 1; end_W(17, 78) <= 1; end_W(17, 79) <= 1; 
end_W(17, 80) <= 0; end_W(17, 81) <= 0; end_W(17, 82) <= 0; end_W(17, 83) <= 0; end_W(17, 84) <= 1; end_W(17, 85) <= 1; end_W(17, 86) <= 1; end_W(17, 87) <= 1; 
end_W(17, 88) <= 1; end_W(17, 89) <= 1; end_W(17, 90) <= 1; end_W(17, 91) <= 1; end_W(17, 92) <= 0; end_W(17, 93) <= 0; end_W(17, 94) <= 0; end_W(17, 95) <= 0; 
end_W(17, 96) <= 1; end_W(17, 97) <= 1; end_W(17, 98) <= 1; end_W(17, 99) <= 1; end_W(17, 100) <= 1; end_W(17, 101) <= 1; end_W(17, 102) <= 1; end_W(17, 103) <= 1; 
end_W(17, 104) <= 0; end_W(17, 105) <= 0; end_W(17, 106) <= 0; end_W(17, 107) <= 0; end_W(17, 108) <= 0; end_W(17, 109) <= 0; end_W(17, 110) <= 0; end_W(17, 111) <= 0; 
end_W(17, 112) <= 1; end_W(17, 113) <= 1; end_W(17, 114) <= 1; end_W(17, 115) <= 1; end_W(17, 116) <= 1; end_W(17, 117) <= 1; end_W(17, 118) <= 1; end_W(17, 119) <= 1; 
end_W(17, 120) <= 1; end_W(17, 121) <= 1; end_W(17, 122) <= 1; end_W(17, 123) <= 1; end_W(17, 124) <= 1; end_W(17, 125) <= 1; end_W(17, 126) <= 1; end_W(17, 127) <= 1; 
end_W(17, 128) <= 0; end_W(17, 129) <= 0; end_W(17, 130) <= 0; end_W(17, 131) <= 0; end_W(17, 132) <= 0; end_W(17, 133) <= 0; end_W(17, 134) <= 0; end_W(17, 135) <= 0; 
end_W(17, 136) <= 0; end_W(17, 137) <= 0; end_W(17, 138) <= 0; end_W(17, 139) <= 0; end_W(17, 140) <= 0; end_W(17, 141) <= 0; end_W(17, 142) <= 0; end_W(17, 143) <= 0; 
end_W(17, 144) <= 0; end_W(17, 145) <= 0; end_W(17, 146) <= 0; end_W(17, 147) <= 0; end_W(17, 148) <= 0; end_W(17, 149) <= 0; end_W(17, 150) <= 0; end_W(17, 151) <= 0; 
end_W(17, 152) <= 0; end_W(17, 153) <= 0; end_W(17, 154) <= 0; end_W(17, 155) <= 0; end_W(17, 156) <= 0; end_W(17, 157) <= 0; end_W(17, 158) <= 0; end_W(17, 159) <= 0; 
end_W(17, 160) <= 0; end_W(17, 161) <= 0; end_W(17, 162) <= 0; end_W(17, 163) <= 0; end_W(17, 164) <= 0; end_W(17, 165) <= 0; end_W(17, 166) <= 0; end_W(17, 167) <= 0; 
end_W(17, 168) <= 0; end_W(17, 169) <= 0; end_W(17, 170) <= 0; end_W(17, 171) <= 0; end_W(17, 172) <= 0; end_W(17, 173) <= 0; end_W(17, 174) <= 0; end_W(17, 175) <= 0; 
end_W(17, 176) <= 0; end_W(17, 177) <= 0; end_W(17, 178) <= 0; end_W(17, 179) <= 0; end_W(17, 180) <= 1; end_W(17, 181) <= 1; end_W(17, 182) <= 1; end_W(17, 183) <= 1; 
end_W(17, 184) <= 1; end_W(17, 185) <= 1; end_W(17, 186) <= 1; end_W(17, 187) <= 1; end_W(17, 188) <= 0; end_W(17, 189) <= 0; end_W(17, 190) <= 0; end_W(17, 191) <= 0; 
end_W(17, 192) <= 0; end_W(17, 193) <= 0; end_W(17, 194) <= 0; end_W(17, 195) <= 0; end_W(17, 196) <= 0; end_W(17, 197) <= 0; end_W(17, 198) <= 0; end_W(17, 199) <= 0; 
end_W(17, 200) <= 1; end_W(17, 201) <= 1; end_W(17, 202) <= 1; end_W(17, 203) <= 1; end_W(17, 204) <= 1; end_W(17, 205) <= 1; end_W(17, 206) <= 1; end_W(17, 207) <= 1; 
end_W(17, 208) <= 0; end_W(17, 209) <= 0; end_W(17, 210) <= 0; end_W(17, 211) <= 0; end_W(17, 212) <= 0; end_W(17, 213) <= 0; end_W(17, 214) <= 0; end_W(17, 215) <= 0; 
end_W(17, 216) <= 1; end_W(17, 217) <= 1; end_W(17, 218) <= 1; end_W(17, 219) <= 1; end_W(17, 220) <= 1; end_W(17, 221) <= 1; end_W(17, 222) <= 1; end_W(17, 223) <= 1; 
end_W(17, 224) <= 0; end_W(17, 225) <= 0; end_W(17, 226) <= 0; end_W(17, 227) <= 0; end_W(17, 228) <= 0; end_W(17, 229) <= 0; end_W(17, 230) <= 0; end_W(17, 231) <= 0; 
end_W(17, 232) <= 0; end_W(17, 233) <= 0; end_W(17, 234) <= 0; end_W(17, 235) <= 0; end_W(17, 236) <= 0; end_W(17, 237) <= 0; end_W(17, 238) <= 0; end_W(17, 239) <= 0; 
end_W(17, 240) <= 1; end_W(17, 241) <= 1; end_W(17, 242) <= 1; end_W(17, 243) <= 1; end_W(17, 244) <= 1; end_W(17, 245) <= 1; end_W(17, 246) <= 1; end_W(17, 247) <= 1; 
end_W(17, 248) <= 0; end_W(17, 249) <= 0; end_W(17, 250) <= 0; end_W(17, 251) <= 0; end_W(17, 252) <= 0; end_W(17, 253) <= 0; end_W(17, 254) <= 0; end_W(17, 255) <= 0; 
end_W(17, 256) <= 1; end_W(17, 257) <= 1; end_W(17, 258) <= 1; end_W(17, 259) <= 1; end_W(17, 260) <= 1; end_W(17, 261) <= 1; end_W(17, 262) <= 1; end_W(17, 263) <= 1; 
end_W(17, 264) <= 1; end_W(17, 265) <= 1; end_W(17, 266) <= 1; end_W(17, 267) <= 1; end_W(17, 268) <= 1; end_W(17, 269) <= 1; end_W(17, 270) <= 1; end_W(17, 271) <= 1; 
end_W(17, 272) <= 0; end_W(17, 273) <= 0; end_W(17, 274) <= 0; end_W(17, 275) <= 0; end_W(17, 276) <= 0; end_W(17, 277) <= 0; end_W(17, 278) <= 0; end_W(17, 279) <= 0; 
end_W(17, 280) <= 0; end_W(17, 281) <= 0; end_W(17, 282) <= 0; end_W(17, 283) <= 0; end_W(17, 284) <= 0; end_W(17, 285) <= 0; end_W(17, 286) <= 0; end_W(17, 287) <= 0; 
end_W(17, 288) <= 0; end_W(17, 289) <= 0; end_W(17, 290) <= 0; end_W(17, 291) <= 0; end_W(17, 292) <= 1; end_W(17, 293) <= 1; end_W(17, 294) <= 1; end_W(17, 295) <= 1; 
end_W(17, 296) <= 1; end_W(17, 297) <= 1; end_W(17, 298) <= 1; end_W(17, 299) <= 1; end_W(17, 300) <= 1; end_W(17, 301) <= 1; end_W(17, 302) <= 1; end_W(17, 303) <= 1; 
end_W(17, 304) <= 1; end_W(17, 305) <= 1; end_W(17, 306) <= 1; end_W(17, 307) <= 1; end_W(17, 308) <= 1; end_W(17, 309) <= 1; end_W(17, 310) <= 1; end_W(17, 311) <= 1; 
end_W(17, 312) <= 0; end_W(17, 313) <= 0; end_W(17, 314) <= 0; end_W(17, 315) <= 0; end_W(17, 316) <= 0; end_W(17, 317) <= 0; end_W(17, 318) <= 0; end_W(17, 319) <= 0; 
end_W(17, 320) <= 0; end_W(17, 321) <= 0; end_W(17, 322) <= 0; end_W(17, 323) <= 0; end_W(18, 0) <= 1; end_W(18, 1) <= 1; end_W(18, 2) <= 1; end_W(18, 3) <= 1; end_W(18, 4) <= 1; end_W(18, 5) <= 1; end_W(18, 6) <= 1; end_W(18, 7) <= 1; 
end_W(18, 8) <= 0; end_W(18, 9) <= 0; end_W(18, 10) <= 0; end_W(18, 11) <= 0; end_W(18, 12) <= 0; end_W(18, 13) <= 0; end_W(18, 14) <= 0; end_W(18, 15) <= 0; 
end_W(18, 16) <= 0; end_W(18, 17) <= 0; end_W(18, 18) <= 0; end_W(18, 19) <= 0; end_W(18, 20) <= 0; end_W(18, 21) <= 0; end_W(18, 22) <= 0; end_W(18, 23) <= 0; 
end_W(18, 24) <= 0; end_W(18, 25) <= 0; end_W(18, 26) <= 0; end_W(18, 27) <= 0; end_W(18, 28) <= 0; end_W(18, 29) <= 0; end_W(18, 30) <= 0; end_W(18, 31) <= 0; 
end_W(18, 32) <= 0; end_W(18, 33) <= 0; end_W(18, 34) <= 0; end_W(18, 35) <= 0; end_W(18, 36) <= 1; end_W(18, 37) <= 1; end_W(18, 38) <= 1; end_W(18, 39) <= 1; 
end_W(18, 40) <= 1; end_W(18, 41) <= 1; end_W(18, 42) <= 1; end_W(18, 43) <= 1; end_W(18, 44) <= 0; end_W(18, 45) <= 0; end_W(18, 46) <= 0; end_W(18, 47) <= 0; 
end_W(18, 48) <= 0; end_W(18, 49) <= 0; end_W(18, 50) <= 0; end_W(18, 51) <= 0; end_W(18, 52) <= 0; end_W(18, 53) <= 0; end_W(18, 54) <= 0; end_W(18, 55) <= 0; 
end_W(18, 56) <= 1; end_W(18, 57) <= 1; end_W(18, 58) <= 1; end_W(18, 59) <= 1; end_W(18, 60) <= 1; end_W(18, 61) <= 1; end_W(18, 62) <= 1; end_W(18, 63) <= 1; 
end_W(18, 64) <= 0; end_W(18, 65) <= 0; end_W(18, 66) <= 0; end_W(18, 67) <= 0; end_W(18, 68) <= 0; end_W(18, 69) <= 0; end_W(18, 70) <= 0; end_W(18, 71) <= 0; 
end_W(18, 72) <= 1; end_W(18, 73) <= 1; end_W(18, 74) <= 1; end_W(18, 75) <= 1; end_W(18, 76) <= 1; end_W(18, 77) <= 1; end_W(18, 78) <= 1; end_W(18, 79) <= 1; 
end_W(18, 80) <= 0; end_W(18, 81) <= 0; end_W(18, 82) <= 0; end_W(18, 83) <= 0; end_W(18, 84) <= 1; end_W(18, 85) <= 1; end_W(18, 86) <= 1; end_W(18, 87) <= 1; 
end_W(18, 88) <= 1; end_W(18, 89) <= 1; end_W(18, 90) <= 1; end_W(18, 91) <= 1; end_W(18, 92) <= 0; end_W(18, 93) <= 0; end_W(18, 94) <= 0; end_W(18, 95) <= 0; 
end_W(18, 96) <= 1; end_W(18, 97) <= 1; end_W(18, 98) <= 1; end_W(18, 99) <= 1; end_W(18, 100) <= 1; end_W(18, 101) <= 1; end_W(18, 102) <= 1; end_W(18, 103) <= 1; 
end_W(18, 104) <= 0; end_W(18, 105) <= 0; end_W(18, 106) <= 0; end_W(18, 107) <= 0; end_W(18, 108) <= 0; end_W(18, 109) <= 0; end_W(18, 110) <= 0; end_W(18, 111) <= 0; 
end_W(18, 112) <= 1; end_W(18, 113) <= 1; end_W(18, 114) <= 1; end_W(18, 115) <= 1; end_W(18, 116) <= 1; end_W(18, 117) <= 1; end_W(18, 118) <= 1; end_W(18, 119) <= 1; 
end_W(18, 120) <= 1; end_W(18, 121) <= 1; end_W(18, 122) <= 1; end_W(18, 123) <= 1; end_W(18, 124) <= 1; end_W(18, 125) <= 1; end_W(18, 126) <= 1; end_W(18, 127) <= 1; 
end_W(18, 128) <= 0; end_W(18, 129) <= 0; end_W(18, 130) <= 0; end_W(18, 131) <= 0; end_W(18, 132) <= 0; end_W(18, 133) <= 0; end_W(18, 134) <= 0; end_W(18, 135) <= 0; 
end_W(18, 136) <= 0; end_W(18, 137) <= 0; end_W(18, 138) <= 0; end_W(18, 139) <= 0; end_W(18, 140) <= 0; end_W(18, 141) <= 0; end_W(18, 142) <= 0; end_W(18, 143) <= 0; 
end_W(18, 144) <= 0; end_W(18, 145) <= 0; end_W(18, 146) <= 0; end_W(18, 147) <= 0; end_W(18, 148) <= 0; end_W(18, 149) <= 0; end_W(18, 150) <= 0; end_W(18, 151) <= 0; 
end_W(18, 152) <= 0; end_W(18, 153) <= 0; end_W(18, 154) <= 0; end_W(18, 155) <= 0; end_W(18, 156) <= 0; end_W(18, 157) <= 0; end_W(18, 158) <= 0; end_W(18, 159) <= 0; 
end_W(18, 160) <= 0; end_W(18, 161) <= 0; end_W(18, 162) <= 0; end_W(18, 163) <= 0; end_W(18, 164) <= 0; end_W(18, 165) <= 0; end_W(18, 166) <= 0; end_W(18, 167) <= 0; 
end_W(18, 168) <= 0; end_W(18, 169) <= 0; end_W(18, 170) <= 0; end_W(18, 171) <= 0; end_W(18, 172) <= 0; end_W(18, 173) <= 0; end_W(18, 174) <= 0; end_W(18, 175) <= 0; 
end_W(18, 176) <= 0; end_W(18, 177) <= 0; end_W(18, 178) <= 0; end_W(18, 179) <= 0; end_W(18, 180) <= 1; end_W(18, 181) <= 1; end_W(18, 182) <= 1; end_W(18, 183) <= 1; 
end_W(18, 184) <= 1; end_W(18, 185) <= 1; end_W(18, 186) <= 1; end_W(18, 187) <= 1; end_W(18, 188) <= 0; end_W(18, 189) <= 0; end_W(18, 190) <= 0; end_W(18, 191) <= 0; 
end_W(18, 192) <= 0; end_W(18, 193) <= 0; end_W(18, 194) <= 0; end_W(18, 195) <= 0; end_W(18, 196) <= 0; end_W(18, 197) <= 0; end_W(18, 198) <= 0; end_W(18, 199) <= 0; 
end_W(18, 200) <= 1; end_W(18, 201) <= 1; end_W(18, 202) <= 1; end_W(18, 203) <= 1; end_W(18, 204) <= 1; end_W(18, 205) <= 1; end_W(18, 206) <= 1; end_W(18, 207) <= 1; 
end_W(18, 208) <= 0; end_W(18, 209) <= 0; end_W(18, 210) <= 0; end_W(18, 211) <= 0; end_W(18, 212) <= 0; end_W(18, 213) <= 0; end_W(18, 214) <= 0; end_W(18, 215) <= 0; 
end_W(18, 216) <= 1; end_W(18, 217) <= 1; end_W(18, 218) <= 1; end_W(18, 219) <= 1; end_W(18, 220) <= 1; end_W(18, 221) <= 1; end_W(18, 222) <= 1; end_W(18, 223) <= 1; 
end_W(18, 224) <= 0; end_W(18, 225) <= 0; end_W(18, 226) <= 0; end_W(18, 227) <= 0; end_W(18, 228) <= 0; end_W(18, 229) <= 0; end_W(18, 230) <= 0; end_W(18, 231) <= 0; 
end_W(18, 232) <= 0; end_W(18, 233) <= 0; end_W(18, 234) <= 0; end_W(18, 235) <= 0; end_W(18, 236) <= 0; end_W(18, 237) <= 0; end_W(18, 238) <= 0; end_W(18, 239) <= 0; 
end_W(18, 240) <= 1; end_W(18, 241) <= 1; end_W(18, 242) <= 1; end_W(18, 243) <= 1; end_W(18, 244) <= 1; end_W(18, 245) <= 1; end_W(18, 246) <= 1; end_W(18, 247) <= 1; 
end_W(18, 248) <= 0; end_W(18, 249) <= 0; end_W(18, 250) <= 0; end_W(18, 251) <= 0; end_W(18, 252) <= 0; end_W(18, 253) <= 0; end_W(18, 254) <= 0; end_W(18, 255) <= 0; 
end_W(18, 256) <= 1; end_W(18, 257) <= 1; end_W(18, 258) <= 1; end_W(18, 259) <= 1; end_W(18, 260) <= 1; end_W(18, 261) <= 1; end_W(18, 262) <= 1; end_W(18, 263) <= 1; 
end_W(18, 264) <= 1; end_W(18, 265) <= 1; end_W(18, 266) <= 1; end_W(18, 267) <= 1; end_W(18, 268) <= 1; end_W(18, 269) <= 1; end_W(18, 270) <= 1; end_W(18, 271) <= 1; 
end_W(18, 272) <= 0; end_W(18, 273) <= 0; end_W(18, 274) <= 0; end_W(18, 275) <= 0; end_W(18, 276) <= 0; end_W(18, 277) <= 0; end_W(18, 278) <= 0; end_W(18, 279) <= 0; 
end_W(18, 280) <= 0; end_W(18, 281) <= 0; end_W(18, 282) <= 0; end_W(18, 283) <= 0; end_W(18, 284) <= 0; end_W(18, 285) <= 0; end_W(18, 286) <= 0; end_W(18, 287) <= 0; 
end_W(18, 288) <= 0; end_W(18, 289) <= 0; end_W(18, 290) <= 0; end_W(18, 291) <= 0; end_W(18, 292) <= 1; end_W(18, 293) <= 1; end_W(18, 294) <= 1; end_W(18, 295) <= 1; 
end_W(18, 296) <= 1; end_W(18, 297) <= 1; end_W(18, 298) <= 1; end_W(18, 299) <= 1; end_W(18, 300) <= 1; end_W(18, 301) <= 1; end_W(18, 302) <= 1; end_W(18, 303) <= 1; 
end_W(18, 304) <= 1; end_W(18, 305) <= 1; end_W(18, 306) <= 1; end_W(18, 307) <= 1; end_W(18, 308) <= 1; end_W(18, 309) <= 1; end_W(18, 310) <= 1; end_W(18, 311) <= 1; 
end_W(18, 312) <= 0; end_W(18, 313) <= 0; end_W(18, 314) <= 0; end_W(18, 315) <= 0; end_W(18, 316) <= 0; end_W(18, 317) <= 0; end_W(18, 318) <= 0; end_W(18, 319) <= 0; 
end_W(18, 320) <= 0; end_W(18, 321) <= 0; end_W(18, 322) <= 0; end_W(18, 323) <= 0; end_W(19, 0) <= 1; end_W(19, 1) <= 1; end_W(19, 2) <= 1; end_W(19, 3) <= 1; end_W(19, 4) <= 1; end_W(19, 5) <= 1; end_W(19, 6) <= 1; end_W(19, 7) <= 1; 
end_W(19, 8) <= 0; end_W(19, 9) <= 0; end_W(19, 10) <= 0; end_W(19, 11) <= 0; end_W(19, 12) <= 0; end_W(19, 13) <= 0; end_W(19, 14) <= 0; end_W(19, 15) <= 0; 
end_W(19, 16) <= 0; end_W(19, 17) <= 0; end_W(19, 18) <= 0; end_W(19, 19) <= 0; end_W(19, 20) <= 0; end_W(19, 21) <= 0; end_W(19, 22) <= 0; end_W(19, 23) <= 0; 
end_W(19, 24) <= 0; end_W(19, 25) <= 0; end_W(19, 26) <= 0; end_W(19, 27) <= 0; end_W(19, 28) <= 0; end_W(19, 29) <= 0; end_W(19, 30) <= 0; end_W(19, 31) <= 0; 
end_W(19, 32) <= 0; end_W(19, 33) <= 0; end_W(19, 34) <= 0; end_W(19, 35) <= 0; end_W(19, 36) <= 1; end_W(19, 37) <= 1; end_W(19, 38) <= 1; end_W(19, 39) <= 1; 
end_W(19, 40) <= 1; end_W(19, 41) <= 1; end_W(19, 42) <= 1; end_W(19, 43) <= 1; end_W(19, 44) <= 0; end_W(19, 45) <= 0; end_W(19, 46) <= 0; end_W(19, 47) <= 0; 
end_W(19, 48) <= 0; end_W(19, 49) <= 0; end_W(19, 50) <= 0; end_W(19, 51) <= 0; end_W(19, 52) <= 0; end_W(19, 53) <= 0; end_W(19, 54) <= 0; end_W(19, 55) <= 0; 
end_W(19, 56) <= 1; end_W(19, 57) <= 1; end_W(19, 58) <= 1; end_W(19, 59) <= 1; end_W(19, 60) <= 1; end_W(19, 61) <= 1; end_W(19, 62) <= 1; end_W(19, 63) <= 1; 
end_W(19, 64) <= 0; end_W(19, 65) <= 0; end_W(19, 66) <= 0; end_W(19, 67) <= 0; end_W(19, 68) <= 0; end_W(19, 69) <= 0; end_W(19, 70) <= 0; end_W(19, 71) <= 0; 
end_W(19, 72) <= 1; end_W(19, 73) <= 1; end_W(19, 74) <= 1; end_W(19, 75) <= 1; end_W(19, 76) <= 1; end_W(19, 77) <= 1; end_W(19, 78) <= 1; end_W(19, 79) <= 1; 
end_W(19, 80) <= 0; end_W(19, 81) <= 0; end_W(19, 82) <= 0; end_W(19, 83) <= 0; end_W(19, 84) <= 1; end_W(19, 85) <= 1; end_W(19, 86) <= 1; end_W(19, 87) <= 1; 
end_W(19, 88) <= 1; end_W(19, 89) <= 1; end_W(19, 90) <= 1; end_W(19, 91) <= 1; end_W(19, 92) <= 0; end_W(19, 93) <= 0; end_W(19, 94) <= 0; end_W(19, 95) <= 0; 
end_W(19, 96) <= 1; end_W(19, 97) <= 1; end_W(19, 98) <= 1; end_W(19, 99) <= 1; end_W(19, 100) <= 1; end_W(19, 101) <= 1; end_W(19, 102) <= 1; end_W(19, 103) <= 1; 
end_W(19, 104) <= 0; end_W(19, 105) <= 0; end_W(19, 106) <= 0; end_W(19, 107) <= 0; end_W(19, 108) <= 0; end_W(19, 109) <= 0; end_W(19, 110) <= 0; end_W(19, 111) <= 0; 
end_W(19, 112) <= 1; end_W(19, 113) <= 1; end_W(19, 114) <= 1; end_W(19, 115) <= 1; end_W(19, 116) <= 1; end_W(19, 117) <= 1; end_W(19, 118) <= 1; end_W(19, 119) <= 1; 
end_W(19, 120) <= 1; end_W(19, 121) <= 1; end_W(19, 122) <= 1; end_W(19, 123) <= 1; end_W(19, 124) <= 1; end_W(19, 125) <= 1; end_W(19, 126) <= 1; end_W(19, 127) <= 1; 
end_W(19, 128) <= 0; end_W(19, 129) <= 0; end_W(19, 130) <= 0; end_W(19, 131) <= 0; end_W(19, 132) <= 0; end_W(19, 133) <= 0; end_W(19, 134) <= 0; end_W(19, 135) <= 0; 
end_W(19, 136) <= 0; end_W(19, 137) <= 0; end_W(19, 138) <= 0; end_W(19, 139) <= 0; end_W(19, 140) <= 0; end_W(19, 141) <= 0; end_W(19, 142) <= 0; end_W(19, 143) <= 0; 
end_W(19, 144) <= 0; end_W(19, 145) <= 0; end_W(19, 146) <= 0; end_W(19, 147) <= 0; end_W(19, 148) <= 0; end_W(19, 149) <= 0; end_W(19, 150) <= 0; end_W(19, 151) <= 0; 
end_W(19, 152) <= 0; end_W(19, 153) <= 0; end_W(19, 154) <= 0; end_W(19, 155) <= 0; end_W(19, 156) <= 0; end_W(19, 157) <= 0; end_W(19, 158) <= 0; end_W(19, 159) <= 0; 
end_W(19, 160) <= 0; end_W(19, 161) <= 0; end_W(19, 162) <= 0; end_W(19, 163) <= 0; end_W(19, 164) <= 0; end_W(19, 165) <= 0; end_W(19, 166) <= 0; end_W(19, 167) <= 0; 
end_W(19, 168) <= 0; end_W(19, 169) <= 0; end_W(19, 170) <= 0; end_W(19, 171) <= 0; end_W(19, 172) <= 0; end_W(19, 173) <= 0; end_W(19, 174) <= 0; end_W(19, 175) <= 0; 
end_W(19, 176) <= 0; end_W(19, 177) <= 0; end_W(19, 178) <= 0; end_W(19, 179) <= 0; end_W(19, 180) <= 1; end_W(19, 181) <= 1; end_W(19, 182) <= 1; end_W(19, 183) <= 1; 
end_W(19, 184) <= 1; end_W(19, 185) <= 1; end_W(19, 186) <= 1; end_W(19, 187) <= 1; end_W(19, 188) <= 0; end_W(19, 189) <= 0; end_W(19, 190) <= 0; end_W(19, 191) <= 0; 
end_W(19, 192) <= 0; end_W(19, 193) <= 0; end_W(19, 194) <= 0; end_W(19, 195) <= 0; end_W(19, 196) <= 0; end_W(19, 197) <= 0; end_W(19, 198) <= 0; end_W(19, 199) <= 0; 
end_W(19, 200) <= 1; end_W(19, 201) <= 1; end_W(19, 202) <= 1; end_W(19, 203) <= 1; end_W(19, 204) <= 1; end_W(19, 205) <= 1; end_W(19, 206) <= 1; end_W(19, 207) <= 1; 
end_W(19, 208) <= 0; end_W(19, 209) <= 0; end_W(19, 210) <= 0; end_W(19, 211) <= 0; end_W(19, 212) <= 0; end_W(19, 213) <= 0; end_W(19, 214) <= 0; end_W(19, 215) <= 0; 
end_W(19, 216) <= 1; end_W(19, 217) <= 1; end_W(19, 218) <= 1; end_W(19, 219) <= 1; end_W(19, 220) <= 1; end_W(19, 221) <= 1; end_W(19, 222) <= 1; end_W(19, 223) <= 1; 
end_W(19, 224) <= 0; end_W(19, 225) <= 0; end_W(19, 226) <= 0; end_W(19, 227) <= 0; end_W(19, 228) <= 0; end_W(19, 229) <= 0; end_W(19, 230) <= 0; end_W(19, 231) <= 0; 
end_W(19, 232) <= 0; end_W(19, 233) <= 0; end_W(19, 234) <= 0; end_W(19, 235) <= 0; end_W(19, 236) <= 0; end_W(19, 237) <= 0; end_W(19, 238) <= 0; end_W(19, 239) <= 0; 
end_W(19, 240) <= 1; end_W(19, 241) <= 1; end_W(19, 242) <= 1; end_W(19, 243) <= 1; end_W(19, 244) <= 1; end_W(19, 245) <= 1; end_W(19, 246) <= 1; end_W(19, 247) <= 1; 
end_W(19, 248) <= 0; end_W(19, 249) <= 0; end_W(19, 250) <= 0; end_W(19, 251) <= 0; end_W(19, 252) <= 0; end_W(19, 253) <= 0; end_W(19, 254) <= 0; end_W(19, 255) <= 0; 
end_W(19, 256) <= 1; end_W(19, 257) <= 1; end_W(19, 258) <= 1; end_W(19, 259) <= 1; end_W(19, 260) <= 1; end_W(19, 261) <= 1; end_W(19, 262) <= 1; end_W(19, 263) <= 1; 
end_W(19, 264) <= 1; end_W(19, 265) <= 1; end_W(19, 266) <= 1; end_W(19, 267) <= 1; end_W(19, 268) <= 1; end_W(19, 269) <= 1; end_W(19, 270) <= 1; end_W(19, 271) <= 1; 
end_W(19, 272) <= 0; end_W(19, 273) <= 0; end_W(19, 274) <= 0; end_W(19, 275) <= 0; end_W(19, 276) <= 0; end_W(19, 277) <= 0; end_W(19, 278) <= 0; end_W(19, 279) <= 0; 
end_W(19, 280) <= 0; end_W(19, 281) <= 0; end_W(19, 282) <= 0; end_W(19, 283) <= 0; end_W(19, 284) <= 0; end_W(19, 285) <= 0; end_W(19, 286) <= 0; end_W(19, 287) <= 0; 
end_W(19, 288) <= 0; end_W(19, 289) <= 0; end_W(19, 290) <= 0; end_W(19, 291) <= 0; end_W(19, 292) <= 1; end_W(19, 293) <= 1; end_W(19, 294) <= 1; end_W(19, 295) <= 1; 
end_W(19, 296) <= 1; end_W(19, 297) <= 1; end_W(19, 298) <= 1; end_W(19, 299) <= 1; end_W(19, 300) <= 1; end_W(19, 301) <= 1; end_W(19, 302) <= 1; end_W(19, 303) <= 1; 
end_W(19, 304) <= 1; end_W(19, 305) <= 1; end_W(19, 306) <= 1; end_W(19, 307) <= 1; end_W(19, 308) <= 1; end_W(19, 309) <= 1; end_W(19, 310) <= 1; end_W(19, 311) <= 1; 
end_W(19, 312) <= 0; end_W(19, 313) <= 0; end_W(19, 314) <= 0; end_W(19, 315) <= 0; end_W(19, 316) <= 0; end_W(19, 317) <= 0; end_W(19, 318) <= 0; end_W(19, 319) <= 0; 
end_W(19, 320) <= 0; end_W(19, 321) <= 0; end_W(19, 322) <= 0; end_W(19, 323) <= 0; end_W(20, 0) <= 1; end_W(20, 1) <= 1; end_W(20, 2) <= 1; end_W(20, 3) <= 1; end_W(20, 4) <= 1; end_W(20, 5) <= 1; end_W(20, 6) <= 1; end_W(20, 7) <= 1; 
end_W(20, 8) <= 0; end_W(20, 9) <= 0; end_W(20, 10) <= 0; end_W(20, 11) <= 0; end_W(20, 12) <= 1; end_W(20, 13) <= 1; end_W(20, 14) <= 1; end_W(20, 15) <= 1; 
end_W(20, 16) <= 1; end_W(20, 17) <= 1; end_W(20, 18) <= 1; end_W(20, 19) <= 1; end_W(20, 20) <= 1; end_W(20, 21) <= 1; end_W(20, 22) <= 1; end_W(20, 23) <= 1; 
end_W(20, 24) <= 1; end_W(20, 25) <= 1; end_W(20, 26) <= 1; end_W(20, 27) <= 1; end_W(20, 28) <= 0; end_W(20, 29) <= 0; end_W(20, 30) <= 0; end_W(20, 31) <= 0; 
end_W(20, 32) <= 0; end_W(20, 33) <= 0; end_W(20, 34) <= 0; end_W(20, 35) <= 0; end_W(20, 36) <= 1; end_W(20, 37) <= 1; end_W(20, 38) <= 1; end_W(20, 39) <= 1; 
end_W(20, 40) <= 1; end_W(20, 41) <= 1; end_W(20, 42) <= 1; end_W(20, 43) <= 1; end_W(20, 44) <= 1; end_W(20, 45) <= 1; end_W(20, 46) <= 1; end_W(20, 47) <= 1; 
end_W(20, 48) <= 1; end_W(20, 49) <= 1; end_W(20, 50) <= 1; end_W(20, 51) <= 1; end_W(20, 52) <= 1; end_W(20, 53) <= 1; end_W(20, 54) <= 1; end_W(20, 55) <= 1; 
end_W(20, 56) <= 1; end_W(20, 57) <= 1; end_W(20, 58) <= 1; end_W(20, 59) <= 1; end_W(20, 60) <= 1; end_W(20, 61) <= 1; end_W(20, 62) <= 1; end_W(20, 63) <= 1; 
end_W(20, 64) <= 0; end_W(20, 65) <= 0; end_W(20, 66) <= 0; end_W(20, 67) <= 0; end_W(20, 68) <= 0; end_W(20, 69) <= 0; end_W(20, 70) <= 0; end_W(20, 71) <= 0; 
end_W(20, 72) <= 1; end_W(20, 73) <= 1; end_W(20, 74) <= 1; end_W(20, 75) <= 1; end_W(20, 76) <= 1; end_W(20, 77) <= 1; end_W(20, 78) <= 1; end_W(20, 79) <= 1; 
end_W(20, 80) <= 0; end_W(20, 81) <= 0; end_W(20, 82) <= 0; end_W(20, 83) <= 0; end_W(20, 84) <= 0; end_W(20, 85) <= 0; end_W(20, 86) <= 0; end_W(20, 87) <= 0; 
end_W(20, 88) <= 0; end_W(20, 89) <= 0; end_W(20, 90) <= 0; end_W(20, 91) <= 0; end_W(20, 92) <= 0; end_W(20, 93) <= 0; end_W(20, 94) <= 0; end_W(20, 95) <= 0; 
end_W(20, 96) <= 1; end_W(20, 97) <= 1; end_W(20, 98) <= 1; end_W(20, 99) <= 1; end_W(20, 100) <= 1; end_W(20, 101) <= 1; end_W(20, 102) <= 1; end_W(20, 103) <= 1; 
end_W(20, 104) <= 0; end_W(20, 105) <= 0; end_W(20, 106) <= 0; end_W(20, 107) <= 0; end_W(20, 108) <= 0; end_W(20, 109) <= 0; end_W(20, 110) <= 0; end_W(20, 111) <= 0; 
end_W(20, 112) <= 1; end_W(20, 113) <= 1; end_W(20, 114) <= 1; end_W(20, 115) <= 1; end_W(20, 116) <= 1; end_W(20, 117) <= 1; end_W(20, 118) <= 1; end_W(20, 119) <= 1; 
end_W(20, 120) <= 0; end_W(20, 121) <= 0; end_W(20, 122) <= 0; end_W(20, 123) <= 0; end_W(20, 124) <= 1; end_W(20, 125) <= 1; end_W(20, 126) <= 1; end_W(20, 127) <= 1; 
end_W(20, 128) <= 0; end_W(20, 129) <= 0; end_W(20, 130) <= 0; end_W(20, 131) <= 0; end_W(20, 132) <= 0; end_W(20, 133) <= 0; end_W(20, 134) <= 0; end_W(20, 135) <= 0; 
end_W(20, 136) <= 0; end_W(20, 137) <= 0; end_W(20, 138) <= 0; end_W(20, 139) <= 0; end_W(20, 140) <= 0; end_W(20, 141) <= 0; end_W(20, 142) <= 0; end_W(20, 143) <= 0; 
end_W(20, 144) <= 0; end_W(20, 145) <= 0; end_W(20, 146) <= 0; end_W(20, 147) <= 0; end_W(20, 148) <= 0; end_W(20, 149) <= 0; end_W(20, 150) <= 0; end_W(20, 151) <= 0; 
end_W(20, 152) <= 0; end_W(20, 153) <= 0; end_W(20, 154) <= 0; end_W(20, 155) <= 0; end_W(20, 156) <= 0; end_W(20, 157) <= 0; end_W(20, 158) <= 0; end_W(20, 159) <= 0; 
end_W(20, 160) <= 0; end_W(20, 161) <= 0; end_W(20, 162) <= 0; end_W(20, 163) <= 0; end_W(20, 164) <= 0; end_W(20, 165) <= 0; end_W(20, 166) <= 0; end_W(20, 167) <= 0; 
end_W(20, 168) <= 0; end_W(20, 169) <= 0; end_W(20, 170) <= 0; end_W(20, 171) <= 0; end_W(20, 172) <= 0; end_W(20, 173) <= 0; end_W(20, 174) <= 0; end_W(20, 175) <= 0; 
end_W(20, 176) <= 0; end_W(20, 177) <= 0; end_W(20, 178) <= 0; end_W(20, 179) <= 0; end_W(20, 180) <= 1; end_W(20, 181) <= 1; end_W(20, 182) <= 1; end_W(20, 183) <= 1; 
end_W(20, 184) <= 1; end_W(20, 185) <= 1; end_W(20, 186) <= 1; end_W(20, 187) <= 1; end_W(20, 188) <= 0; end_W(20, 189) <= 0; end_W(20, 190) <= 0; end_W(20, 191) <= 0; 
end_W(20, 192) <= 0; end_W(20, 193) <= 0; end_W(20, 194) <= 0; end_W(20, 195) <= 0; end_W(20, 196) <= 0; end_W(20, 197) <= 0; end_W(20, 198) <= 0; end_W(20, 199) <= 0; 
end_W(20, 200) <= 1; end_W(20, 201) <= 1; end_W(20, 202) <= 1; end_W(20, 203) <= 1; end_W(20, 204) <= 1; end_W(20, 205) <= 1; end_W(20, 206) <= 1; end_W(20, 207) <= 1; 
end_W(20, 208) <= 0; end_W(20, 209) <= 0; end_W(20, 210) <= 0; end_W(20, 211) <= 0; end_W(20, 212) <= 0; end_W(20, 213) <= 0; end_W(20, 214) <= 0; end_W(20, 215) <= 0; 
end_W(20, 216) <= 1; end_W(20, 217) <= 1; end_W(20, 218) <= 1; end_W(20, 219) <= 1; end_W(20, 220) <= 1; end_W(20, 221) <= 1; end_W(20, 222) <= 1; end_W(20, 223) <= 1; 
end_W(20, 224) <= 0; end_W(20, 225) <= 0; end_W(20, 226) <= 0; end_W(20, 227) <= 0; end_W(20, 228) <= 0; end_W(20, 229) <= 0; end_W(20, 230) <= 0; end_W(20, 231) <= 0; 
end_W(20, 232) <= 0; end_W(20, 233) <= 0; end_W(20, 234) <= 0; end_W(20, 235) <= 0; end_W(20, 236) <= 0; end_W(20, 237) <= 0; end_W(20, 238) <= 0; end_W(20, 239) <= 0; 
end_W(20, 240) <= 1; end_W(20, 241) <= 1; end_W(20, 242) <= 1; end_W(20, 243) <= 1; end_W(20, 244) <= 1; end_W(20, 245) <= 1; end_W(20, 246) <= 1; end_W(20, 247) <= 1; 
end_W(20, 248) <= 0; end_W(20, 249) <= 0; end_W(20, 250) <= 0; end_W(20, 251) <= 0; end_W(20, 252) <= 0; end_W(20, 253) <= 0; end_W(20, 254) <= 0; end_W(20, 255) <= 0; 
end_W(20, 256) <= 1; end_W(20, 257) <= 1; end_W(20, 258) <= 1; end_W(20, 259) <= 1; end_W(20, 260) <= 1; end_W(20, 261) <= 1; end_W(20, 262) <= 1; end_W(20, 263) <= 1; 
end_W(20, 264) <= 0; end_W(20, 265) <= 0; end_W(20, 266) <= 0; end_W(20, 267) <= 0; end_W(20, 268) <= 1; end_W(20, 269) <= 1; end_W(20, 270) <= 1; end_W(20, 271) <= 1; 
end_W(20, 272) <= 0; end_W(20, 273) <= 0; end_W(20, 274) <= 0; end_W(20, 275) <= 0; end_W(20, 276) <= 0; end_W(20, 277) <= 0; end_W(20, 278) <= 0; end_W(20, 279) <= 0; 
end_W(20, 280) <= 0; end_W(20, 281) <= 0; end_W(20, 282) <= 0; end_W(20, 283) <= 0; end_W(20, 284) <= 0; end_W(20, 285) <= 0; end_W(20, 286) <= 0; end_W(20, 287) <= 0; 
end_W(20, 288) <= 0; end_W(20, 289) <= 0; end_W(20, 290) <= 0; end_W(20, 291) <= 0; end_W(20, 292) <= 1; end_W(20, 293) <= 1; end_W(20, 294) <= 1; end_W(20, 295) <= 1; 
end_W(20, 296) <= 1; end_W(20, 297) <= 1; end_W(20, 298) <= 1; end_W(20, 299) <= 1; end_W(20, 300) <= 0; end_W(20, 301) <= 0; end_W(20, 302) <= 0; end_W(20, 303) <= 0; 
end_W(20, 304) <= 1; end_W(20, 305) <= 1; end_W(20, 306) <= 1; end_W(20, 307) <= 1; end_W(20, 308) <= 1; end_W(20, 309) <= 1; end_W(20, 310) <= 1; end_W(20, 311) <= 1; 
end_W(20, 312) <= 0; end_W(20, 313) <= 0; end_W(20, 314) <= 0; end_W(20, 315) <= 0; end_W(20, 316) <= 0; end_W(20, 317) <= 0; end_W(20, 318) <= 0; end_W(20, 319) <= 0; 
end_W(20, 320) <= 0; end_W(20, 321) <= 0; end_W(20, 322) <= 0; end_W(20, 323) <= 0; end_W(21, 0) <= 1; end_W(21, 1) <= 1; end_W(21, 2) <= 1; end_W(21, 3) <= 1; end_W(21, 4) <= 1; end_W(21, 5) <= 1; end_W(21, 6) <= 1; end_W(21, 7) <= 1; 
end_W(21, 8) <= 0; end_W(21, 9) <= 0; end_W(21, 10) <= 0; end_W(21, 11) <= 0; end_W(21, 12) <= 1; end_W(21, 13) <= 1; end_W(21, 14) <= 1; end_W(21, 15) <= 1; 
end_W(21, 16) <= 1; end_W(21, 17) <= 1; end_W(21, 18) <= 1; end_W(21, 19) <= 1; end_W(21, 20) <= 1; end_W(21, 21) <= 1; end_W(21, 22) <= 1; end_W(21, 23) <= 1; 
end_W(21, 24) <= 1; end_W(21, 25) <= 1; end_W(21, 26) <= 1; end_W(21, 27) <= 1; end_W(21, 28) <= 0; end_W(21, 29) <= 0; end_W(21, 30) <= 0; end_W(21, 31) <= 0; 
end_W(21, 32) <= 0; end_W(21, 33) <= 0; end_W(21, 34) <= 0; end_W(21, 35) <= 0; end_W(21, 36) <= 1; end_W(21, 37) <= 1; end_W(21, 38) <= 1; end_W(21, 39) <= 1; 
end_W(21, 40) <= 1; end_W(21, 41) <= 1; end_W(21, 42) <= 1; end_W(21, 43) <= 1; end_W(21, 44) <= 1; end_W(21, 45) <= 1; end_W(21, 46) <= 1; end_W(21, 47) <= 1; 
end_W(21, 48) <= 1; end_W(21, 49) <= 1; end_W(21, 50) <= 1; end_W(21, 51) <= 1; end_W(21, 52) <= 1; end_W(21, 53) <= 1; end_W(21, 54) <= 1; end_W(21, 55) <= 1; 
end_W(21, 56) <= 1; end_W(21, 57) <= 1; end_W(21, 58) <= 1; end_W(21, 59) <= 1; end_W(21, 60) <= 1; end_W(21, 61) <= 1; end_W(21, 62) <= 1; end_W(21, 63) <= 1; 
end_W(21, 64) <= 0; end_W(21, 65) <= 0; end_W(21, 66) <= 0; end_W(21, 67) <= 0; end_W(21, 68) <= 0; end_W(21, 69) <= 0; end_W(21, 70) <= 0; end_W(21, 71) <= 0; 
end_W(21, 72) <= 1; end_W(21, 73) <= 1; end_W(21, 74) <= 1; end_W(21, 75) <= 1; end_W(21, 76) <= 1; end_W(21, 77) <= 1; end_W(21, 78) <= 1; end_W(21, 79) <= 1; 
end_W(21, 80) <= 0; end_W(21, 81) <= 0; end_W(21, 82) <= 0; end_W(21, 83) <= 0; end_W(21, 84) <= 0; end_W(21, 85) <= 0; end_W(21, 86) <= 0; end_W(21, 87) <= 0; 
end_W(21, 88) <= 0; end_W(21, 89) <= 0; end_W(21, 90) <= 0; end_W(21, 91) <= 0; end_W(21, 92) <= 0; end_W(21, 93) <= 0; end_W(21, 94) <= 0; end_W(21, 95) <= 0; 
end_W(21, 96) <= 1; end_W(21, 97) <= 1; end_W(21, 98) <= 1; end_W(21, 99) <= 1; end_W(21, 100) <= 1; end_W(21, 101) <= 1; end_W(21, 102) <= 1; end_W(21, 103) <= 1; 
end_W(21, 104) <= 0; end_W(21, 105) <= 0; end_W(21, 106) <= 0; end_W(21, 107) <= 0; end_W(21, 108) <= 0; end_W(21, 109) <= 0; end_W(21, 110) <= 0; end_W(21, 111) <= 0; 
end_W(21, 112) <= 1; end_W(21, 113) <= 1; end_W(21, 114) <= 1; end_W(21, 115) <= 1; end_W(21, 116) <= 1; end_W(21, 117) <= 1; end_W(21, 118) <= 1; end_W(21, 119) <= 1; 
end_W(21, 120) <= 0; end_W(21, 121) <= 0; end_W(21, 122) <= 0; end_W(21, 123) <= 0; end_W(21, 124) <= 1; end_W(21, 125) <= 1; end_W(21, 126) <= 1; end_W(21, 127) <= 1; 
end_W(21, 128) <= 0; end_W(21, 129) <= 0; end_W(21, 130) <= 0; end_W(21, 131) <= 0; end_W(21, 132) <= 0; end_W(21, 133) <= 0; end_W(21, 134) <= 0; end_W(21, 135) <= 0; 
end_W(21, 136) <= 0; end_W(21, 137) <= 0; end_W(21, 138) <= 0; end_W(21, 139) <= 0; end_W(21, 140) <= 0; end_W(21, 141) <= 0; end_W(21, 142) <= 0; end_W(21, 143) <= 0; 
end_W(21, 144) <= 0; end_W(21, 145) <= 0; end_W(21, 146) <= 0; end_W(21, 147) <= 0; end_W(21, 148) <= 0; end_W(21, 149) <= 0; end_W(21, 150) <= 0; end_W(21, 151) <= 0; 
end_W(21, 152) <= 0; end_W(21, 153) <= 0; end_W(21, 154) <= 0; end_W(21, 155) <= 0; end_W(21, 156) <= 0; end_W(21, 157) <= 0; end_W(21, 158) <= 0; end_W(21, 159) <= 0; 
end_W(21, 160) <= 0; end_W(21, 161) <= 0; end_W(21, 162) <= 0; end_W(21, 163) <= 0; end_W(21, 164) <= 0; end_W(21, 165) <= 0; end_W(21, 166) <= 0; end_W(21, 167) <= 0; 
end_W(21, 168) <= 0; end_W(21, 169) <= 0; end_W(21, 170) <= 0; end_W(21, 171) <= 0; end_W(21, 172) <= 0; end_W(21, 173) <= 0; end_W(21, 174) <= 0; end_W(21, 175) <= 0; 
end_W(21, 176) <= 0; end_W(21, 177) <= 0; end_W(21, 178) <= 0; end_W(21, 179) <= 0; end_W(21, 180) <= 1; end_W(21, 181) <= 1; end_W(21, 182) <= 1; end_W(21, 183) <= 1; 
end_W(21, 184) <= 1; end_W(21, 185) <= 1; end_W(21, 186) <= 1; end_W(21, 187) <= 1; end_W(21, 188) <= 0; end_W(21, 189) <= 0; end_W(21, 190) <= 0; end_W(21, 191) <= 0; 
end_W(21, 192) <= 0; end_W(21, 193) <= 0; end_W(21, 194) <= 0; end_W(21, 195) <= 0; end_W(21, 196) <= 0; end_W(21, 197) <= 0; end_W(21, 198) <= 0; end_W(21, 199) <= 0; 
end_W(21, 200) <= 1; end_W(21, 201) <= 1; end_W(21, 202) <= 1; end_W(21, 203) <= 1; end_W(21, 204) <= 1; end_W(21, 205) <= 1; end_W(21, 206) <= 1; end_W(21, 207) <= 1; 
end_W(21, 208) <= 0; end_W(21, 209) <= 0; end_W(21, 210) <= 0; end_W(21, 211) <= 0; end_W(21, 212) <= 0; end_W(21, 213) <= 0; end_W(21, 214) <= 0; end_W(21, 215) <= 0; 
end_W(21, 216) <= 1; end_W(21, 217) <= 1; end_W(21, 218) <= 1; end_W(21, 219) <= 1; end_W(21, 220) <= 1; end_W(21, 221) <= 1; end_W(21, 222) <= 1; end_W(21, 223) <= 1; 
end_W(21, 224) <= 0; end_W(21, 225) <= 0; end_W(21, 226) <= 0; end_W(21, 227) <= 0; end_W(21, 228) <= 0; end_W(21, 229) <= 0; end_W(21, 230) <= 0; end_W(21, 231) <= 0; 
end_W(21, 232) <= 0; end_W(21, 233) <= 0; end_W(21, 234) <= 0; end_W(21, 235) <= 0; end_W(21, 236) <= 0; end_W(21, 237) <= 0; end_W(21, 238) <= 0; end_W(21, 239) <= 0; 
end_W(21, 240) <= 1; end_W(21, 241) <= 1; end_W(21, 242) <= 1; end_W(21, 243) <= 1; end_W(21, 244) <= 1; end_W(21, 245) <= 1; end_W(21, 246) <= 1; end_W(21, 247) <= 1; 
end_W(21, 248) <= 0; end_W(21, 249) <= 0; end_W(21, 250) <= 0; end_W(21, 251) <= 0; end_W(21, 252) <= 0; end_W(21, 253) <= 0; end_W(21, 254) <= 0; end_W(21, 255) <= 0; 
end_W(21, 256) <= 1; end_W(21, 257) <= 1; end_W(21, 258) <= 1; end_W(21, 259) <= 1; end_W(21, 260) <= 1; end_W(21, 261) <= 1; end_W(21, 262) <= 1; end_W(21, 263) <= 1; 
end_W(21, 264) <= 0; end_W(21, 265) <= 0; end_W(21, 266) <= 0; end_W(21, 267) <= 0; end_W(21, 268) <= 1; end_W(21, 269) <= 1; end_W(21, 270) <= 1; end_W(21, 271) <= 1; 
end_W(21, 272) <= 0; end_W(21, 273) <= 0; end_W(21, 274) <= 0; end_W(21, 275) <= 0; end_W(21, 276) <= 0; end_W(21, 277) <= 0; end_W(21, 278) <= 0; end_W(21, 279) <= 0; 
end_W(21, 280) <= 0; end_W(21, 281) <= 0; end_W(21, 282) <= 0; end_W(21, 283) <= 0; end_W(21, 284) <= 0; end_W(21, 285) <= 0; end_W(21, 286) <= 0; end_W(21, 287) <= 0; 
end_W(21, 288) <= 0; end_W(21, 289) <= 0; end_W(21, 290) <= 0; end_W(21, 291) <= 0; end_W(21, 292) <= 1; end_W(21, 293) <= 1; end_W(21, 294) <= 1; end_W(21, 295) <= 1; 
end_W(21, 296) <= 1; end_W(21, 297) <= 1; end_W(21, 298) <= 1; end_W(21, 299) <= 1; end_W(21, 300) <= 0; end_W(21, 301) <= 0; end_W(21, 302) <= 0; end_W(21, 303) <= 0; 
end_W(21, 304) <= 1; end_W(21, 305) <= 1; end_W(21, 306) <= 1; end_W(21, 307) <= 1; end_W(21, 308) <= 1; end_W(21, 309) <= 1; end_W(21, 310) <= 1; end_W(21, 311) <= 1; 
end_W(21, 312) <= 0; end_W(21, 313) <= 0; end_W(21, 314) <= 0; end_W(21, 315) <= 0; end_W(21, 316) <= 0; end_W(21, 317) <= 0; end_W(21, 318) <= 0; end_W(21, 319) <= 0; 
end_W(21, 320) <= 0; end_W(21, 321) <= 0; end_W(21, 322) <= 0; end_W(21, 323) <= 0; end_W(22, 0) <= 1; end_W(22, 1) <= 1; end_W(22, 2) <= 1; end_W(22, 3) <= 1; end_W(22, 4) <= 1; end_W(22, 5) <= 1; end_W(22, 6) <= 1; end_W(22, 7) <= 1; 
end_W(22, 8) <= 0; end_W(22, 9) <= 0; end_W(22, 10) <= 0; end_W(22, 11) <= 0; end_W(22, 12) <= 1; end_W(22, 13) <= 1; end_W(22, 14) <= 1; end_W(22, 15) <= 1; 
end_W(22, 16) <= 1; end_W(22, 17) <= 1; end_W(22, 18) <= 1; end_W(22, 19) <= 1; end_W(22, 20) <= 1; end_W(22, 21) <= 1; end_W(22, 22) <= 1; end_W(22, 23) <= 1; 
end_W(22, 24) <= 1; end_W(22, 25) <= 1; end_W(22, 26) <= 1; end_W(22, 27) <= 1; end_W(22, 28) <= 0; end_W(22, 29) <= 0; end_W(22, 30) <= 0; end_W(22, 31) <= 0; 
end_W(22, 32) <= 0; end_W(22, 33) <= 0; end_W(22, 34) <= 0; end_W(22, 35) <= 0; end_W(22, 36) <= 1; end_W(22, 37) <= 1; end_W(22, 38) <= 1; end_W(22, 39) <= 1; 
end_W(22, 40) <= 1; end_W(22, 41) <= 1; end_W(22, 42) <= 1; end_W(22, 43) <= 1; end_W(22, 44) <= 1; end_W(22, 45) <= 1; end_W(22, 46) <= 1; end_W(22, 47) <= 1; 
end_W(22, 48) <= 1; end_W(22, 49) <= 1; end_W(22, 50) <= 1; end_W(22, 51) <= 1; end_W(22, 52) <= 1; end_W(22, 53) <= 1; end_W(22, 54) <= 1; end_W(22, 55) <= 1; 
end_W(22, 56) <= 1; end_W(22, 57) <= 1; end_W(22, 58) <= 1; end_W(22, 59) <= 1; end_W(22, 60) <= 1; end_W(22, 61) <= 1; end_W(22, 62) <= 1; end_W(22, 63) <= 1; 
end_W(22, 64) <= 0; end_W(22, 65) <= 0; end_W(22, 66) <= 0; end_W(22, 67) <= 0; end_W(22, 68) <= 0; end_W(22, 69) <= 0; end_W(22, 70) <= 0; end_W(22, 71) <= 0; 
end_W(22, 72) <= 1; end_W(22, 73) <= 1; end_W(22, 74) <= 1; end_W(22, 75) <= 1; end_W(22, 76) <= 1; end_W(22, 77) <= 1; end_W(22, 78) <= 1; end_W(22, 79) <= 1; 
end_W(22, 80) <= 0; end_W(22, 81) <= 0; end_W(22, 82) <= 0; end_W(22, 83) <= 0; end_W(22, 84) <= 0; end_W(22, 85) <= 0; end_W(22, 86) <= 0; end_W(22, 87) <= 0; 
end_W(22, 88) <= 0; end_W(22, 89) <= 0; end_W(22, 90) <= 0; end_W(22, 91) <= 0; end_W(22, 92) <= 0; end_W(22, 93) <= 0; end_W(22, 94) <= 0; end_W(22, 95) <= 0; 
end_W(22, 96) <= 1; end_W(22, 97) <= 1; end_W(22, 98) <= 1; end_W(22, 99) <= 1; end_W(22, 100) <= 1; end_W(22, 101) <= 1; end_W(22, 102) <= 1; end_W(22, 103) <= 1; 
end_W(22, 104) <= 0; end_W(22, 105) <= 0; end_W(22, 106) <= 0; end_W(22, 107) <= 0; end_W(22, 108) <= 0; end_W(22, 109) <= 0; end_W(22, 110) <= 0; end_W(22, 111) <= 0; 
end_W(22, 112) <= 1; end_W(22, 113) <= 1; end_W(22, 114) <= 1; end_W(22, 115) <= 1; end_W(22, 116) <= 1; end_W(22, 117) <= 1; end_W(22, 118) <= 1; end_W(22, 119) <= 1; 
end_W(22, 120) <= 0; end_W(22, 121) <= 0; end_W(22, 122) <= 0; end_W(22, 123) <= 0; end_W(22, 124) <= 1; end_W(22, 125) <= 1; end_W(22, 126) <= 1; end_W(22, 127) <= 1; 
end_W(22, 128) <= 0; end_W(22, 129) <= 0; end_W(22, 130) <= 0; end_W(22, 131) <= 0; end_W(22, 132) <= 0; end_W(22, 133) <= 0; end_W(22, 134) <= 0; end_W(22, 135) <= 0; 
end_W(22, 136) <= 0; end_W(22, 137) <= 0; end_W(22, 138) <= 0; end_W(22, 139) <= 0; end_W(22, 140) <= 0; end_W(22, 141) <= 0; end_W(22, 142) <= 0; end_W(22, 143) <= 0; 
end_W(22, 144) <= 0; end_W(22, 145) <= 0; end_W(22, 146) <= 0; end_W(22, 147) <= 0; end_W(22, 148) <= 0; end_W(22, 149) <= 0; end_W(22, 150) <= 0; end_W(22, 151) <= 0; 
end_W(22, 152) <= 0; end_W(22, 153) <= 0; end_W(22, 154) <= 0; end_W(22, 155) <= 0; end_W(22, 156) <= 0; end_W(22, 157) <= 0; end_W(22, 158) <= 0; end_W(22, 159) <= 0; 
end_W(22, 160) <= 0; end_W(22, 161) <= 0; end_W(22, 162) <= 0; end_W(22, 163) <= 0; end_W(22, 164) <= 0; end_W(22, 165) <= 0; end_W(22, 166) <= 0; end_W(22, 167) <= 0; 
end_W(22, 168) <= 0; end_W(22, 169) <= 0; end_W(22, 170) <= 0; end_W(22, 171) <= 0; end_W(22, 172) <= 0; end_W(22, 173) <= 0; end_W(22, 174) <= 0; end_W(22, 175) <= 0; 
end_W(22, 176) <= 0; end_W(22, 177) <= 0; end_W(22, 178) <= 0; end_W(22, 179) <= 0; end_W(22, 180) <= 1; end_W(22, 181) <= 1; end_W(22, 182) <= 1; end_W(22, 183) <= 1; 
end_W(22, 184) <= 1; end_W(22, 185) <= 1; end_W(22, 186) <= 1; end_W(22, 187) <= 1; end_W(22, 188) <= 0; end_W(22, 189) <= 0; end_W(22, 190) <= 0; end_W(22, 191) <= 0; 
end_W(22, 192) <= 0; end_W(22, 193) <= 0; end_W(22, 194) <= 0; end_W(22, 195) <= 0; end_W(22, 196) <= 0; end_W(22, 197) <= 0; end_W(22, 198) <= 0; end_W(22, 199) <= 0; 
end_W(22, 200) <= 1; end_W(22, 201) <= 1; end_W(22, 202) <= 1; end_W(22, 203) <= 1; end_W(22, 204) <= 1; end_W(22, 205) <= 1; end_W(22, 206) <= 1; end_W(22, 207) <= 1; 
end_W(22, 208) <= 0; end_W(22, 209) <= 0; end_W(22, 210) <= 0; end_W(22, 211) <= 0; end_W(22, 212) <= 0; end_W(22, 213) <= 0; end_W(22, 214) <= 0; end_W(22, 215) <= 0; 
end_W(22, 216) <= 1; end_W(22, 217) <= 1; end_W(22, 218) <= 1; end_W(22, 219) <= 1; end_W(22, 220) <= 1; end_W(22, 221) <= 1; end_W(22, 222) <= 1; end_W(22, 223) <= 1; 
end_W(22, 224) <= 0; end_W(22, 225) <= 0; end_W(22, 226) <= 0; end_W(22, 227) <= 0; end_W(22, 228) <= 0; end_W(22, 229) <= 0; end_W(22, 230) <= 0; end_W(22, 231) <= 0; 
end_W(22, 232) <= 0; end_W(22, 233) <= 0; end_W(22, 234) <= 0; end_W(22, 235) <= 0; end_W(22, 236) <= 0; end_W(22, 237) <= 0; end_W(22, 238) <= 0; end_W(22, 239) <= 0; 
end_W(22, 240) <= 1; end_W(22, 241) <= 1; end_W(22, 242) <= 1; end_W(22, 243) <= 1; end_W(22, 244) <= 1; end_W(22, 245) <= 1; end_W(22, 246) <= 1; end_W(22, 247) <= 1; 
end_W(22, 248) <= 0; end_W(22, 249) <= 0; end_W(22, 250) <= 0; end_W(22, 251) <= 0; end_W(22, 252) <= 0; end_W(22, 253) <= 0; end_W(22, 254) <= 0; end_W(22, 255) <= 0; 
end_W(22, 256) <= 1; end_W(22, 257) <= 1; end_W(22, 258) <= 1; end_W(22, 259) <= 1; end_W(22, 260) <= 1; end_W(22, 261) <= 1; end_W(22, 262) <= 1; end_W(22, 263) <= 1; 
end_W(22, 264) <= 0; end_W(22, 265) <= 0; end_W(22, 266) <= 0; end_W(22, 267) <= 0; end_W(22, 268) <= 1; end_W(22, 269) <= 1; end_W(22, 270) <= 1; end_W(22, 271) <= 1; 
end_W(22, 272) <= 0; end_W(22, 273) <= 0; end_W(22, 274) <= 0; end_W(22, 275) <= 0; end_W(22, 276) <= 0; end_W(22, 277) <= 0; end_W(22, 278) <= 0; end_W(22, 279) <= 0; 
end_W(22, 280) <= 0; end_W(22, 281) <= 0; end_W(22, 282) <= 0; end_W(22, 283) <= 0; end_W(22, 284) <= 0; end_W(22, 285) <= 0; end_W(22, 286) <= 0; end_W(22, 287) <= 0; 
end_W(22, 288) <= 0; end_W(22, 289) <= 0; end_W(22, 290) <= 0; end_W(22, 291) <= 0; end_W(22, 292) <= 1; end_W(22, 293) <= 1; end_W(22, 294) <= 1; end_W(22, 295) <= 1; 
end_W(22, 296) <= 1; end_W(22, 297) <= 1; end_W(22, 298) <= 1; end_W(22, 299) <= 1; end_W(22, 300) <= 0; end_W(22, 301) <= 0; end_W(22, 302) <= 0; end_W(22, 303) <= 0; 
end_W(22, 304) <= 1; end_W(22, 305) <= 1; end_W(22, 306) <= 1; end_W(22, 307) <= 1; end_W(22, 308) <= 1; end_W(22, 309) <= 1; end_W(22, 310) <= 1; end_W(22, 311) <= 1; 
end_W(22, 312) <= 0; end_W(22, 313) <= 0; end_W(22, 314) <= 0; end_W(22, 315) <= 0; end_W(22, 316) <= 0; end_W(22, 317) <= 0; end_W(22, 318) <= 0; end_W(22, 319) <= 0; 
end_W(22, 320) <= 0; end_W(22, 321) <= 0; end_W(22, 322) <= 0; end_W(22, 323) <= 0; end_W(23, 0) <= 1; end_W(23, 1) <= 1; end_W(23, 2) <= 1; end_W(23, 3) <= 1; end_W(23, 4) <= 1; end_W(23, 5) <= 1; end_W(23, 6) <= 1; end_W(23, 7) <= 1; 
end_W(23, 8) <= 0; end_W(23, 9) <= 0; end_W(23, 10) <= 0; end_W(23, 11) <= 0; end_W(23, 12) <= 1; end_W(23, 13) <= 1; end_W(23, 14) <= 1; end_W(23, 15) <= 1; 
end_W(23, 16) <= 1; end_W(23, 17) <= 1; end_W(23, 18) <= 1; end_W(23, 19) <= 1; end_W(23, 20) <= 1; end_W(23, 21) <= 1; end_W(23, 22) <= 1; end_W(23, 23) <= 1; 
end_W(23, 24) <= 1; end_W(23, 25) <= 1; end_W(23, 26) <= 1; end_W(23, 27) <= 1; end_W(23, 28) <= 0; end_W(23, 29) <= 0; end_W(23, 30) <= 0; end_W(23, 31) <= 0; 
end_W(23, 32) <= 0; end_W(23, 33) <= 0; end_W(23, 34) <= 0; end_W(23, 35) <= 0; end_W(23, 36) <= 1; end_W(23, 37) <= 1; end_W(23, 38) <= 1; end_W(23, 39) <= 1; 
end_W(23, 40) <= 1; end_W(23, 41) <= 1; end_W(23, 42) <= 1; end_W(23, 43) <= 1; end_W(23, 44) <= 1; end_W(23, 45) <= 1; end_W(23, 46) <= 1; end_W(23, 47) <= 1; 
end_W(23, 48) <= 1; end_W(23, 49) <= 1; end_W(23, 50) <= 1; end_W(23, 51) <= 1; end_W(23, 52) <= 1; end_W(23, 53) <= 1; end_W(23, 54) <= 1; end_W(23, 55) <= 1; 
end_W(23, 56) <= 1; end_W(23, 57) <= 1; end_W(23, 58) <= 1; end_W(23, 59) <= 1; end_W(23, 60) <= 1; end_W(23, 61) <= 1; end_W(23, 62) <= 1; end_W(23, 63) <= 1; 
end_W(23, 64) <= 0; end_W(23, 65) <= 0; end_W(23, 66) <= 0; end_W(23, 67) <= 0; end_W(23, 68) <= 0; end_W(23, 69) <= 0; end_W(23, 70) <= 0; end_W(23, 71) <= 0; 
end_W(23, 72) <= 1; end_W(23, 73) <= 1; end_W(23, 74) <= 1; end_W(23, 75) <= 1; end_W(23, 76) <= 1; end_W(23, 77) <= 1; end_W(23, 78) <= 1; end_W(23, 79) <= 1; 
end_W(23, 80) <= 0; end_W(23, 81) <= 0; end_W(23, 82) <= 0; end_W(23, 83) <= 0; end_W(23, 84) <= 0; end_W(23, 85) <= 0; end_W(23, 86) <= 0; end_W(23, 87) <= 0; 
end_W(23, 88) <= 0; end_W(23, 89) <= 0; end_W(23, 90) <= 0; end_W(23, 91) <= 0; end_W(23, 92) <= 0; end_W(23, 93) <= 0; end_W(23, 94) <= 0; end_W(23, 95) <= 0; 
end_W(23, 96) <= 1; end_W(23, 97) <= 1; end_W(23, 98) <= 1; end_W(23, 99) <= 1; end_W(23, 100) <= 1; end_W(23, 101) <= 1; end_W(23, 102) <= 1; end_W(23, 103) <= 1; 
end_W(23, 104) <= 0; end_W(23, 105) <= 0; end_W(23, 106) <= 0; end_W(23, 107) <= 0; end_W(23, 108) <= 0; end_W(23, 109) <= 0; end_W(23, 110) <= 0; end_W(23, 111) <= 0; 
end_W(23, 112) <= 1; end_W(23, 113) <= 1; end_W(23, 114) <= 1; end_W(23, 115) <= 1; end_W(23, 116) <= 1; end_W(23, 117) <= 1; end_W(23, 118) <= 1; end_W(23, 119) <= 1; 
end_W(23, 120) <= 0; end_W(23, 121) <= 0; end_W(23, 122) <= 0; end_W(23, 123) <= 0; end_W(23, 124) <= 1; end_W(23, 125) <= 1; end_W(23, 126) <= 1; end_W(23, 127) <= 1; 
end_W(23, 128) <= 0; end_W(23, 129) <= 0; end_W(23, 130) <= 0; end_W(23, 131) <= 0; end_W(23, 132) <= 0; end_W(23, 133) <= 0; end_W(23, 134) <= 0; end_W(23, 135) <= 0; 
end_W(23, 136) <= 0; end_W(23, 137) <= 0; end_W(23, 138) <= 0; end_W(23, 139) <= 0; end_W(23, 140) <= 0; end_W(23, 141) <= 0; end_W(23, 142) <= 0; end_W(23, 143) <= 0; 
end_W(23, 144) <= 0; end_W(23, 145) <= 0; end_W(23, 146) <= 0; end_W(23, 147) <= 0; end_W(23, 148) <= 0; end_W(23, 149) <= 0; end_W(23, 150) <= 0; end_W(23, 151) <= 0; 
end_W(23, 152) <= 0; end_W(23, 153) <= 0; end_W(23, 154) <= 0; end_W(23, 155) <= 0; end_W(23, 156) <= 0; end_W(23, 157) <= 0; end_W(23, 158) <= 0; end_W(23, 159) <= 0; 
end_W(23, 160) <= 0; end_W(23, 161) <= 0; end_W(23, 162) <= 0; end_W(23, 163) <= 0; end_W(23, 164) <= 0; end_W(23, 165) <= 0; end_W(23, 166) <= 0; end_W(23, 167) <= 0; 
end_W(23, 168) <= 0; end_W(23, 169) <= 0; end_W(23, 170) <= 0; end_W(23, 171) <= 0; end_W(23, 172) <= 0; end_W(23, 173) <= 0; end_W(23, 174) <= 0; end_W(23, 175) <= 0; 
end_W(23, 176) <= 0; end_W(23, 177) <= 0; end_W(23, 178) <= 0; end_W(23, 179) <= 0; end_W(23, 180) <= 1; end_W(23, 181) <= 1; end_W(23, 182) <= 1; end_W(23, 183) <= 1; 
end_W(23, 184) <= 1; end_W(23, 185) <= 1; end_W(23, 186) <= 1; end_W(23, 187) <= 1; end_W(23, 188) <= 0; end_W(23, 189) <= 0; end_W(23, 190) <= 0; end_W(23, 191) <= 0; 
end_W(23, 192) <= 0; end_W(23, 193) <= 0; end_W(23, 194) <= 0; end_W(23, 195) <= 0; end_W(23, 196) <= 0; end_W(23, 197) <= 0; end_W(23, 198) <= 0; end_W(23, 199) <= 0; 
end_W(23, 200) <= 1; end_W(23, 201) <= 1; end_W(23, 202) <= 1; end_W(23, 203) <= 1; end_W(23, 204) <= 1; end_W(23, 205) <= 1; end_W(23, 206) <= 1; end_W(23, 207) <= 1; 
end_W(23, 208) <= 0; end_W(23, 209) <= 0; end_W(23, 210) <= 0; end_W(23, 211) <= 0; end_W(23, 212) <= 0; end_W(23, 213) <= 0; end_W(23, 214) <= 0; end_W(23, 215) <= 0; 
end_W(23, 216) <= 1; end_W(23, 217) <= 1; end_W(23, 218) <= 1; end_W(23, 219) <= 1; end_W(23, 220) <= 1; end_W(23, 221) <= 1; end_W(23, 222) <= 1; end_W(23, 223) <= 1; 
end_W(23, 224) <= 0; end_W(23, 225) <= 0; end_W(23, 226) <= 0; end_W(23, 227) <= 0; end_W(23, 228) <= 0; end_W(23, 229) <= 0; end_W(23, 230) <= 0; end_W(23, 231) <= 0; 
end_W(23, 232) <= 0; end_W(23, 233) <= 0; end_W(23, 234) <= 0; end_W(23, 235) <= 0; end_W(23, 236) <= 0; end_W(23, 237) <= 0; end_W(23, 238) <= 0; end_W(23, 239) <= 0; 
end_W(23, 240) <= 1; end_W(23, 241) <= 1; end_W(23, 242) <= 1; end_W(23, 243) <= 1; end_W(23, 244) <= 1; end_W(23, 245) <= 1; end_W(23, 246) <= 1; end_W(23, 247) <= 1; 
end_W(23, 248) <= 0; end_W(23, 249) <= 0; end_W(23, 250) <= 0; end_W(23, 251) <= 0; end_W(23, 252) <= 0; end_W(23, 253) <= 0; end_W(23, 254) <= 0; end_W(23, 255) <= 0; 
end_W(23, 256) <= 1; end_W(23, 257) <= 1; end_W(23, 258) <= 1; end_W(23, 259) <= 1; end_W(23, 260) <= 1; end_W(23, 261) <= 1; end_W(23, 262) <= 1; end_W(23, 263) <= 1; 
end_W(23, 264) <= 0; end_W(23, 265) <= 0; end_W(23, 266) <= 0; end_W(23, 267) <= 0; end_W(23, 268) <= 1; end_W(23, 269) <= 1; end_W(23, 270) <= 1; end_W(23, 271) <= 1; 
end_W(23, 272) <= 0; end_W(23, 273) <= 0; end_W(23, 274) <= 0; end_W(23, 275) <= 0; end_W(23, 276) <= 0; end_W(23, 277) <= 0; end_W(23, 278) <= 0; end_W(23, 279) <= 0; 
end_W(23, 280) <= 0; end_W(23, 281) <= 0; end_W(23, 282) <= 0; end_W(23, 283) <= 0; end_W(23, 284) <= 0; end_W(23, 285) <= 0; end_W(23, 286) <= 0; end_W(23, 287) <= 0; 
end_W(23, 288) <= 0; end_W(23, 289) <= 0; end_W(23, 290) <= 0; end_W(23, 291) <= 0; end_W(23, 292) <= 1; end_W(23, 293) <= 1; end_W(23, 294) <= 1; end_W(23, 295) <= 1; 
end_W(23, 296) <= 1; end_W(23, 297) <= 1; end_W(23, 298) <= 1; end_W(23, 299) <= 1; end_W(23, 300) <= 0; end_W(23, 301) <= 0; end_W(23, 302) <= 0; end_W(23, 303) <= 0; 
end_W(23, 304) <= 1; end_W(23, 305) <= 1; end_W(23, 306) <= 1; end_W(23, 307) <= 1; end_W(23, 308) <= 1; end_W(23, 309) <= 1; end_W(23, 310) <= 1; end_W(23, 311) <= 1; 
end_W(23, 312) <= 0; end_W(23, 313) <= 0; end_W(23, 314) <= 0; end_W(23, 315) <= 0; end_W(23, 316) <= 0; end_W(23, 317) <= 0; end_W(23, 318) <= 0; end_W(23, 319) <= 0; 
end_W(23, 320) <= 0; end_W(23, 321) <= 0; end_W(23, 322) <= 0; end_W(23, 323) <= 0; end_W(24, 0) <= 1; end_W(24, 1) <= 1; end_W(24, 2) <= 1; end_W(24, 3) <= 1; end_W(24, 4) <= 1; end_W(24, 5) <= 1; end_W(24, 6) <= 1; end_W(24, 7) <= 1; 
end_W(24, 8) <= 0; end_W(24, 9) <= 0; end_W(24, 10) <= 0; end_W(24, 11) <= 0; end_W(24, 12) <= 0; end_W(24, 13) <= 0; end_W(24, 14) <= 0; end_W(24, 15) <= 0; 
end_W(24, 16) <= 0; end_W(24, 17) <= 0; end_W(24, 18) <= 0; end_W(24, 19) <= 0; end_W(24, 20) <= 1; end_W(24, 21) <= 1; end_W(24, 22) <= 1; end_W(24, 23) <= 1; 
end_W(24, 24) <= 1; end_W(24, 25) <= 1; end_W(24, 26) <= 1; end_W(24, 27) <= 1; end_W(24, 28) <= 0; end_W(24, 29) <= 0; end_W(24, 30) <= 0; end_W(24, 31) <= 0; 
end_W(24, 32) <= 0; end_W(24, 33) <= 0; end_W(24, 34) <= 0; end_W(24, 35) <= 0; end_W(24, 36) <= 1; end_W(24, 37) <= 1; end_W(24, 38) <= 1; end_W(24, 39) <= 1; 
end_W(24, 40) <= 1; end_W(24, 41) <= 1; end_W(24, 42) <= 1; end_W(24, 43) <= 1; end_W(24, 44) <= 0; end_W(24, 45) <= 0; end_W(24, 46) <= 0; end_W(24, 47) <= 0; 
end_W(24, 48) <= 0; end_W(24, 49) <= 0; end_W(24, 50) <= 0; end_W(24, 51) <= 0; end_W(24, 52) <= 0; end_W(24, 53) <= 0; end_W(24, 54) <= 0; end_W(24, 55) <= 0; 
end_W(24, 56) <= 1; end_W(24, 57) <= 1; end_W(24, 58) <= 1; end_W(24, 59) <= 1; end_W(24, 60) <= 1; end_W(24, 61) <= 1; end_W(24, 62) <= 1; end_W(24, 63) <= 1; 
end_W(24, 64) <= 0; end_W(24, 65) <= 0; end_W(24, 66) <= 0; end_W(24, 67) <= 0; end_W(24, 68) <= 0; end_W(24, 69) <= 0; end_W(24, 70) <= 0; end_W(24, 71) <= 0; 
end_W(24, 72) <= 1; end_W(24, 73) <= 1; end_W(24, 74) <= 1; end_W(24, 75) <= 1; end_W(24, 76) <= 1; end_W(24, 77) <= 1; end_W(24, 78) <= 1; end_W(24, 79) <= 1; 
end_W(24, 80) <= 0; end_W(24, 81) <= 0; end_W(24, 82) <= 0; end_W(24, 83) <= 0; end_W(24, 84) <= 0; end_W(24, 85) <= 0; end_W(24, 86) <= 0; end_W(24, 87) <= 0; 
end_W(24, 88) <= 0; end_W(24, 89) <= 0; end_W(24, 90) <= 0; end_W(24, 91) <= 0; end_W(24, 92) <= 0; end_W(24, 93) <= 0; end_W(24, 94) <= 0; end_W(24, 95) <= 0; 
end_W(24, 96) <= 1; end_W(24, 97) <= 1; end_W(24, 98) <= 1; end_W(24, 99) <= 1; end_W(24, 100) <= 1; end_W(24, 101) <= 1; end_W(24, 102) <= 1; end_W(24, 103) <= 1; 
end_W(24, 104) <= 0; end_W(24, 105) <= 0; end_W(24, 106) <= 0; end_W(24, 107) <= 0; end_W(24, 108) <= 0; end_W(24, 109) <= 0; end_W(24, 110) <= 0; end_W(24, 111) <= 0; 
end_W(24, 112) <= 1; end_W(24, 113) <= 1; end_W(24, 114) <= 1; end_W(24, 115) <= 1; end_W(24, 116) <= 1; end_W(24, 117) <= 1; end_W(24, 118) <= 1; end_W(24, 119) <= 1; 
end_W(24, 120) <= 0; end_W(24, 121) <= 0; end_W(24, 122) <= 0; end_W(24, 123) <= 0; end_W(24, 124) <= 0; end_W(24, 125) <= 0; end_W(24, 126) <= 0; end_W(24, 127) <= 0; 
end_W(24, 128) <= 0; end_W(24, 129) <= 0; end_W(24, 130) <= 0; end_W(24, 131) <= 0; end_W(24, 132) <= 0; end_W(24, 133) <= 0; end_W(24, 134) <= 0; end_W(24, 135) <= 0; 
end_W(24, 136) <= 0; end_W(24, 137) <= 0; end_W(24, 138) <= 0; end_W(24, 139) <= 0; end_W(24, 140) <= 0; end_W(24, 141) <= 0; end_W(24, 142) <= 0; end_W(24, 143) <= 0; 
end_W(24, 144) <= 0; end_W(24, 145) <= 0; end_W(24, 146) <= 0; end_W(24, 147) <= 0; end_W(24, 148) <= 0; end_W(24, 149) <= 0; end_W(24, 150) <= 0; end_W(24, 151) <= 0; 
end_W(24, 152) <= 0; end_W(24, 153) <= 0; end_W(24, 154) <= 0; end_W(24, 155) <= 0; end_W(24, 156) <= 0; end_W(24, 157) <= 0; end_W(24, 158) <= 0; end_W(24, 159) <= 0; 
end_W(24, 160) <= 0; end_W(24, 161) <= 0; end_W(24, 162) <= 0; end_W(24, 163) <= 0; end_W(24, 164) <= 0; end_W(24, 165) <= 0; end_W(24, 166) <= 0; end_W(24, 167) <= 0; 
end_W(24, 168) <= 0; end_W(24, 169) <= 0; end_W(24, 170) <= 0; end_W(24, 171) <= 0; end_W(24, 172) <= 0; end_W(24, 173) <= 0; end_W(24, 174) <= 0; end_W(24, 175) <= 0; 
end_W(24, 176) <= 0; end_W(24, 177) <= 0; end_W(24, 178) <= 0; end_W(24, 179) <= 0; end_W(24, 180) <= 1; end_W(24, 181) <= 1; end_W(24, 182) <= 1; end_W(24, 183) <= 1; 
end_W(24, 184) <= 1; end_W(24, 185) <= 1; end_W(24, 186) <= 1; end_W(24, 187) <= 1; end_W(24, 188) <= 0; end_W(24, 189) <= 0; end_W(24, 190) <= 0; end_W(24, 191) <= 0; 
end_W(24, 192) <= 0; end_W(24, 193) <= 0; end_W(24, 194) <= 0; end_W(24, 195) <= 0; end_W(24, 196) <= 0; end_W(24, 197) <= 0; end_W(24, 198) <= 0; end_W(24, 199) <= 0; 
end_W(24, 200) <= 1; end_W(24, 201) <= 1; end_W(24, 202) <= 1; end_W(24, 203) <= 1; end_W(24, 204) <= 1; end_W(24, 205) <= 1; end_W(24, 206) <= 1; end_W(24, 207) <= 1; 
end_W(24, 208) <= 0; end_W(24, 209) <= 0; end_W(24, 210) <= 0; end_W(24, 211) <= 0; end_W(24, 212) <= 0; end_W(24, 213) <= 0; end_W(24, 214) <= 0; end_W(24, 215) <= 0; 
end_W(24, 216) <= 1; end_W(24, 217) <= 1; end_W(24, 218) <= 1; end_W(24, 219) <= 1; end_W(24, 220) <= 1; end_W(24, 221) <= 1; end_W(24, 222) <= 1; end_W(24, 223) <= 1; 
end_W(24, 224) <= 0; end_W(24, 225) <= 0; end_W(24, 226) <= 0; end_W(24, 227) <= 0; end_W(24, 228) <= 0; end_W(24, 229) <= 0; end_W(24, 230) <= 0; end_W(24, 231) <= 0; 
end_W(24, 232) <= 0; end_W(24, 233) <= 0; end_W(24, 234) <= 0; end_W(24, 235) <= 0; end_W(24, 236) <= 0; end_W(24, 237) <= 0; end_W(24, 238) <= 0; end_W(24, 239) <= 0; 
end_W(24, 240) <= 1; end_W(24, 241) <= 1; end_W(24, 242) <= 1; end_W(24, 243) <= 1; end_W(24, 244) <= 1; end_W(24, 245) <= 1; end_W(24, 246) <= 1; end_W(24, 247) <= 1; 
end_W(24, 248) <= 0; end_W(24, 249) <= 0; end_W(24, 250) <= 0; end_W(24, 251) <= 0; end_W(24, 252) <= 0; end_W(24, 253) <= 0; end_W(24, 254) <= 0; end_W(24, 255) <= 0; 
end_W(24, 256) <= 1; end_W(24, 257) <= 1; end_W(24, 258) <= 1; end_W(24, 259) <= 1; end_W(24, 260) <= 1; end_W(24, 261) <= 1; end_W(24, 262) <= 1; end_W(24, 263) <= 1; 
end_W(24, 264) <= 0; end_W(24, 265) <= 0; end_W(24, 266) <= 0; end_W(24, 267) <= 0; end_W(24, 268) <= 0; end_W(24, 269) <= 0; end_W(24, 270) <= 0; end_W(24, 271) <= 0; 
end_W(24, 272) <= 0; end_W(24, 273) <= 0; end_W(24, 274) <= 0; end_W(24, 275) <= 0; end_W(24, 276) <= 0; end_W(24, 277) <= 0; end_W(24, 278) <= 0; end_W(24, 279) <= 0; 
end_W(24, 280) <= 0; end_W(24, 281) <= 0; end_W(24, 282) <= 0; end_W(24, 283) <= 0; end_W(24, 284) <= 0; end_W(24, 285) <= 0; end_W(24, 286) <= 0; end_W(24, 287) <= 0; 
end_W(24, 288) <= 0; end_W(24, 289) <= 0; end_W(24, 290) <= 0; end_W(24, 291) <= 0; end_W(24, 292) <= 1; end_W(24, 293) <= 1; end_W(24, 294) <= 1; end_W(24, 295) <= 1; 
end_W(24, 296) <= 1; end_W(24, 297) <= 1; end_W(24, 298) <= 1; end_W(24, 299) <= 1; end_W(24, 300) <= 0; end_W(24, 301) <= 0; end_W(24, 302) <= 0; end_W(24, 303) <= 0; 
end_W(24, 304) <= 0; end_W(24, 305) <= 0; end_W(24, 306) <= 0; end_W(24, 307) <= 0; end_W(24, 308) <= 1; end_W(24, 309) <= 1; end_W(24, 310) <= 1; end_W(24, 311) <= 1; 
end_W(24, 312) <= 1; end_W(24, 313) <= 1; end_W(24, 314) <= 1; end_W(24, 315) <= 1; end_W(24, 316) <= 0; end_W(24, 317) <= 0; end_W(24, 318) <= 0; end_W(24, 319) <= 0; 
end_W(24, 320) <= 0; end_W(24, 321) <= 0; end_W(24, 322) <= 0; end_W(24, 323) <= 0; end_W(25, 0) <= 1; end_W(25, 1) <= 1; end_W(25, 2) <= 1; end_W(25, 3) <= 1; end_W(25, 4) <= 1; end_W(25, 5) <= 1; end_W(25, 6) <= 1; end_W(25, 7) <= 1; 
end_W(25, 8) <= 0; end_W(25, 9) <= 0; end_W(25, 10) <= 0; end_W(25, 11) <= 0; end_W(25, 12) <= 0; end_W(25, 13) <= 0; end_W(25, 14) <= 0; end_W(25, 15) <= 0; 
end_W(25, 16) <= 0; end_W(25, 17) <= 0; end_W(25, 18) <= 0; end_W(25, 19) <= 0; end_W(25, 20) <= 1; end_W(25, 21) <= 1; end_W(25, 22) <= 1; end_W(25, 23) <= 1; 
end_W(25, 24) <= 1; end_W(25, 25) <= 1; end_W(25, 26) <= 1; end_W(25, 27) <= 1; end_W(25, 28) <= 0; end_W(25, 29) <= 0; end_W(25, 30) <= 0; end_W(25, 31) <= 0; 
end_W(25, 32) <= 0; end_W(25, 33) <= 0; end_W(25, 34) <= 0; end_W(25, 35) <= 0; end_W(25, 36) <= 1; end_W(25, 37) <= 1; end_W(25, 38) <= 1; end_W(25, 39) <= 1; 
end_W(25, 40) <= 1; end_W(25, 41) <= 1; end_W(25, 42) <= 1; end_W(25, 43) <= 1; end_W(25, 44) <= 0; end_W(25, 45) <= 0; end_W(25, 46) <= 0; end_W(25, 47) <= 0; 
end_W(25, 48) <= 0; end_W(25, 49) <= 0; end_W(25, 50) <= 0; end_W(25, 51) <= 0; end_W(25, 52) <= 0; end_W(25, 53) <= 0; end_W(25, 54) <= 0; end_W(25, 55) <= 0; 
end_W(25, 56) <= 1; end_W(25, 57) <= 1; end_W(25, 58) <= 1; end_W(25, 59) <= 1; end_W(25, 60) <= 1; end_W(25, 61) <= 1; end_W(25, 62) <= 1; end_W(25, 63) <= 1; 
end_W(25, 64) <= 0; end_W(25, 65) <= 0; end_W(25, 66) <= 0; end_W(25, 67) <= 0; end_W(25, 68) <= 0; end_W(25, 69) <= 0; end_W(25, 70) <= 0; end_W(25, 71) <= 0; 
end_W(25, 72) <= 1; end_W(25, 73) <= 1; end_W(25, 74) <= 1; end_W(25, 75) <= 1; end_W(25, 76) <= 1; end_W(25, 77) <= 1; end_W(25, 78) <= 1; end_W(25, 79) <= 1; 
end_W(25, 80) <= 0; end_W(25, 81) <= 0; end_W(25, 82) <= 0; end_W(25, 83) <= 0; end_W(25, 84) <= 0; end_W(25, 85) <= 0; end_W(25, 86) <= 0; end_W(25, 87) <= 0; 
end_W(25, 88) <= 0; end_W(25, 89) <= 0; end_W(25, 90) <= 0; end_W(25, 91) <= 0; end_W(25, 92) <= 0; end_W(25, 93) <= 0; end_W(25, 94) <= 0; end_W(25, 95) <= 0; 
end_W(25, 96) <= 1; end_W(25, 97) <= 1; end_W(25, 98) <= 1; end_W(25, 99) <= 1; end_W(25, 100) <= 1; end_W(25, 101) <= 1; end_W(25, 102) <= 1; end_W(25, 103) <= 1; 
end_W(25, 104) <= 0; end_W(25, 105) <= 0; end_W(25, 106) <= 0; end_W(25, 107) <= 0; end_W(25, 108) <= 0; end_W(25, 109) <= 0; end_W(25, 110) <= 0; end_W(25, 111) <= 0; 
end_W(25, 112) <= 1; end_W(25, 113) <= 1; end_W(25, 114) <= 1; end_W(25, 115) <= 1; end_W(25, 116) <= 1; end_W(25, 117) <= 1; end_W(25, 118) <= 1; end_W(25, 119) <= 1; 
end_W(25, 120) <= 0; end_W(25, 121) <= 0; end_W(25, 122) <= 0; end_W(25, 123) <= 0; end_W(25, 124) <= 0; end_W(25, 125) <= 0; end_W(25, 126) <= 0; end_W(25, 127) <= 0; 
end_W(25, 128) <= 0; end_W(25, 129) <= 0; end_W(25, 130) <= 0; end_W(25, 131) <= 0; end_W(25, 132) <= 0; end_W(25, 133) <= 0; end_W(25, 134) <= 0; end_W(25, 135) <= 0; 
end_W(25, 136) <= 0; end_W(25, 137) <= 0; end_W(25, 138) <= 0; end_W(25, 139) <= 0; end_W(25, 140) <= 0; end_W(25, 141) <= 0; end_W(25, 142) <= 0; end_W(25, 143) <= 0; 
end_W(25, 144) <= 0; end_W(25, 145) <= 0; end_W(25, 146) <= 0; end_W(25, 147) <= 0; end_W(25, 148) <= 0; end_W(25, 149) <= 0; end_W(25, 150) <= 0; end_W(25, 151) <= 0; 
end_W(25, 152) <= 0; end_W(25, 153) <= 0; end_W(25, 154) <= 0; end_W(25, 155) <= 0; end_W(25, 156) <= 0; end_W(25, 157) <= 0; end_W(25, 158) <= 0; end_W(25, 159) <= 0; 
end_W(25, 160) <= 0; end_W(25, 161) <= 0; end_W(25, 162) <= 0; end_W(25, 163) <= 0; end_W(25, 164) <= 0; end_W(25, 165) <= 0; end_W(25, 166) <= 0; end_W(25, 167) <= 0; 
end_W(25, 168) <= 0; end_W(25, 169) <= 0; end_W(25, 170) <= 0; end_W(25, 171) <= 0; end_W(25, 172) <= 0; end_W(25, 173) <= 0; end_W(25, 174) <= 0; end_W(25, 175) <= 0; 
end_W(25, 176) <= 0; end_W(25, 177) <= 0; end_W(25, 178) <= 0; end_W(25, 179) <= 0; end_W(25, 180) <= 1; end_W(25, 181) <= 1; end_W(25, 182) <= 1; end_W(25, 183) <= 1; 
end_W(25, 184) <= 1; end_W(25, 185) <= 1; end_W(25, 186) <= 1; end_W(25, 187) <= 1; end_W(25, 188) <= 0; end_W(25, 189) <= 0; end_W(25, 190) <= 0; end_W(25, 191) <= 0; 
end_W(25, 192) <= 0; end_W(25, 193) <= 0; end_W(25, 194) <= 0; end_W(25, 195) <= 0; end_W(25, 196) <= 0; end_W(25, 197) <= 0; end_W(25, 198) <= 0; end_W(25, 199) <= 0; 
end_W(25, 200) <= 1; end_W(25, 201) <= 1; end_W(25, 202) <= 1; end_W(25, 203) <= 1; end_W(25, 204) <= 1; end_W(25, 205) <= 1; end_W(25, 206) <= 1; end_W(25, 207) <= 1; 
end_W(25, 208) <= 0; end_W(25, 209) <= 0; end_W(25, 210) <= 0; end_W(25, 211) <= 0; end_W(25, 212) <= 0; end_W(25, 213) <= 0; end_W(25, 214) <= 0; end_W(25, 215) <= 0; 
end_W(25, 216) <= 1; end_W(25, 217) <= 1; end_W(25, 218) <= 1; end_W(25, 219) <= 1; end_W(25, 220) <= 1; end_W(25, 221) <= 1; end_W(25, 222) <= 1; end_W(25, 223) <= 1; 
end_W(25, 224) <= 0; end_W(25, 225) <= 0; end_W(25, 226) <= 0; end_W(25, 227) <= 0; end_W(25, 228) <= 0; end_W(25, 229) <= 0; end_W(25, 230) <= 0; end_W(25, 231) <= 0; 
end_W(25, 232) <= 0; end_W(25, 233) <= 0; end_W(25, 234) <= 0; end_W(25, 235) <= 0; end_W(25, 236) <= 0; end_W(25, 237) <= 0; end_W(25, 238) <= 0; end_W(25, 239) <= 0; 
end_W(25, 240) <= 1; end_W(25, 241) <= 1; end_W(25, 242) <= 1; end_W(25, 243) <= 1; end_W(25, 244) <= 1; end_W(25, 245) <= 1; end_W(25, 246) <= 1; end_W(25, 247) <= 1; 
end_W(25, 248) <= 0; end_W(25, 249) <= 0; end_W(25, 250) <= 0; end_W(25, 251) <= 0; end_W(25, 252) <= 0; end_W(25, 253) <= 0; end_W(25, 254) <= 0; end_W(25, 255) <= 0; 
end_W(25, 256) <= 1; end_W(25, 257) <= 1; end_W(25, 258) <= 1; end_W(25, 259) <= 1; end_W(25, 260) <= 1; end_W(25, 261) <= 1; end_W(25, 262) <= 1; end_W(25, 263) <= 1; 
end_W(25, 264) <= 0; end_W(25, 265) <= 0; end_W(25, 266) <= 0; end_W(25, 267) <= 0; end_W(25, 268) <= 0; end_W(25, 269) <= 0; end_W(25, 270) <= 0; end_W(25, 271) <= 0; 
end_W(25, 272) <= 0; end_W(25, 273) <= 0; end_W(25, 274) <= 0; end_W(25, 275) <= 0; end_W(25, 276) <= 0; end_W(25, 277) <= 0; end_W(25, 278) <= 0; end_W(25, 279) <= 0; 
end_W(25, 280) <= 0; end_W(25, 281) <= 0; end_W(25, 282) <= 0; end_W(25, 283) <= 0; end_W(25, 284) <= 0; end_W(25, 285) <= 0; end_W(25, 286) <= 0; end_W(25, 287) <= 0; 
end_W(25, 288) <= 0; end_W(25, 289) <= 0; end_W(25, 290) <= 0; end_W(25, 291) <= 0; end_W(25, 292) <= 1; end_W(25, 293) <= 1; end_W(25, 294) <= 1; end_W(25, 295) <= 1; 
end_W(25, 296) <= 1; end_W(25, 297) <= 1; end_W(25, 298) <= 1; end_W(25, 299) <= 1; end_W(25, 300) <= 0; end_W(25, 301) <= 0; end_W(25, 302) <= 0; end_W(25, 303) <= 0; 
end_W(25, 304) <= 0; end_W(25, 305) <= 0; end_W(25, 306) <= 0; end_W(25, 307) <= 0; end_W(25, 308) <= 1; end_W(25, 309) <= 1; end_W(25, 310) <= 1; end_W(25, 311) <= 1; 
end_W(25, 312) <= 1; end_W(25, 313) <= 1; end_W(25, 314) <= 1; end_W(25, 315) <= 1; end_W(25, 316) <= 0; end_W(25, 317) <= 0; end_W(25, 318) <= 0; end_W(25, 319) <= 0; 
end_W(25, 320) <= 0; end_W(25, 321) <= 0; end_W(25, 322) <= 0; end_W(25, 323) <= 0; end_W(26, 0) <= 1; end_W(26, 1) <= 1; end_W(26, 2) <= 1; end_W(26, 3) <= 1; end_W(26, 4) <= 1; end_W(26, 5) <= 1; end_W(26, 6) <= 1; end_W(26, 7) <= 1; 
end_W(26, 8) <= 0; end_W(26, 9) <= 0; end_W(26, 10) <= 0; end_W(26, 11) <= 0; end_W(26, 12) <= 0; end_W(26, 13) <= 0; end_W(26, 14) <= 0; end_W(26, 15) <= 0; 
end_W(26, 16) <= 0; end_W(26, 17) <= 0; end_W(26, 18) <= 0; end_W(26, 19) <= 0; end_W(26, 20) <= 1; end_W(26, 21) <= 1; end_W(26, 22) <= 1; end_W(26, 23) <= 1; 
end_W(26, 24) <= 1; end_W(26, 25) <= 1; end_W(26, 26) <= 1; end_W(26, 27) <= 1; end_W(26, 28) <= 0; end_W(26, 29) <= 0; end_W(26, 30) <= 0; end_W(26, 31) <= 0; 
end_W(26, 32) <= 0; end_W(26, 33) <= 0; end_W(26, 34) <= 0; end_W(26, 35) <= 0; end_W(26, 36) <= 1; end_W(26, 37) <= 1; end_W(26, 38) <= 1; end_W(26, 39) <= 1; 
end_W(26, 40) <= 1; end_W(26, 41) <= 1; end_W(26, 42) <= 1; end_W(26, 43) <= 1; end_W(26, 44) <= 0; end_W(26, 45) <= 0; end_W(26, 46) <= 0; end_W(26, 47) <= 0; 
end_W(26, 48) <= 0; end_W(26, 49) <= 0; end_W(26, 50) <= 0; end_W(26, 51) <= 0; end_W(26, 52) <= 0; end_W(26, 53) <= 0; end_W(26, 54) <= 0; end_W(26, 55) <= 0; 
end_W(26, 56) <= 1; end_W(26, 57) <= 1; end_W(26, 58) <= 1; end_W(26, 59) <= 1; end_W(26, 60) <= 1; end_W(26, 61) <= 1; end_W(26, 62) <= 1; end_W(26, 63) <= 1; 
end_W(26, 64) <= 0; end_W(26, 65) <= 0; end_W(26, 66) <= 0; end_W(26, 67) <= 0; end_W(26, 68) <= 0; end_W(26, 69) <= 0; end_W(26, 70) <= 0; end_W(26, 71) <= 0; 
end_W(26, 72) <= 1; end_W(26, 73) <= 1; end_W(26, 74) <= 1; end_W(26, 75) <= 1; end_W(26, 76) <= 1; end_W(26, 77) <= 1; end_W(26, 78) <= 1; end_W(26, 79) <= 1; 
end_W(26, 80) <= 0; end_W(26, 81) <= 0; end_W(26, 82) <= 0; end_W(26, 83) <= 0; end_W(26, 84) <= 0; end_W(26, 85) <= 0; end_W(26, 86) <= 0; end_W(26, 87) <= 0; 
end_W(26, 88) <= 0; end_W(26, 89) <= 0; end_W(26, 90) <= 0; end_W(26, 91) <= 0; end_W(26, 92) <= 0; end_W(26, 93) <= 0; end_W(26, 94) <= 0; end_W(26, 95) <= 0; 
end_W(26, 96) <= 1; end_W(26, 97) <= 1; end_W(26, 98) <= 1; end_W(26, 99) <= 1; end_W(26, 100) <= 1; end_W(26, 101) <= 1; end_W(26, 102) <= 1; end_W(26, 103) <= 1; 
end_W(26, 104) <= 0; end_W(26, 105) <= 0; end_W(26, 106) <= 0; end_W(26, 107) <= 0; end_W(26, 108) <= 0; end_W(26, 109) <= 0; end_W(26, 110) <= 0; end_W(26, 111) <= 0; 
end_W(26, 112) <= 1; end_W(26, 113) <= 1; end_W(26, 114) <= 1; end_W(26, 115) <= 1; end_W(26, 116) <= 1; end_W(26, 117) <= 1; end_W(26, 118) <= 1; end_W(26, 119) <= 1; 
end_W(26, 120) <= 0; end_W(26, 121) <= 0; end_W(26, 122) <= 0; end_W(26, 123) <= 0; end_W(26, 124) <= 0; end_W(26, 125) <= 0; end_W(26, 126) <= 0; end_W(26, 127) <= 0; 
end_W(26, 128) <= 0; end_W(26, 129) <= 0; end_W(26, 130) <= 0; end_W(26, 131) <= 0; end_W(26, 132) <= 0; end_W(26, 133) <= 0; end_W(26, 134) <= 0; end_W(26, 135) <= 0; 
end_W(26, 136) <= 0; end_W(26, 137) <= 0; end_W(26, 138) <= 0; end_W(26, 139) <= 0; end_W(26, 140) <= 0; end_W(26, 141) <= 0; end_W(26, 142) <= 0; end_W(26, 143) <= 0; 
end_W(26, 144) <= 0; end_W(26, 145) <= 0; end_W(26, 146) <= 0; end_W(26, 147) <= 0; end_W(26, 148) <= 0; end_W(26, 149) <= 0; end_W(26, 150) <= 0; end_W(26, 151) <= 0; 
end_W(26, 152) <= 0; end_W(26, 153) <= 0; end_W(26, 154) <= 0; end_W(26, 155) <= 0; end_W(26, 156) <= 0; end_W(26, 157) <= 0; end_W(26, 158) <= 0; end_W(26, 159) <= 0; 
end_W(26, 160) <= 0; end_W(26, 161) <= 0; end_W(26, 162) <= 0; end_W(26, 163) <= 0; end_W(26, 164) <= 0; end_W(26, 165) <= 0; end_W(26, 166) <= 0; end_W(26, 167) <= 0; 
end_W(26, 168) <= 0; end_W(26, 169) <= 0; end_W(26, 170) <= 0; end_W(26, 171) <= 0; end_W(26, 172) <= 0; end_W(26, 173) <= 0; end_W(26, 174) <= 0; end_W(26, 175) <= 0; 
end_W(26, 176) <= 0; end_W(26, 177) <= 0; end_W(26, 178) <= 0; end_W(26, 179) <= 0; end_W(26, 180) <= 1; end_W(26, 181) <= 1; end_W(26, 182) <= 1; end_W(26, 183) <= 1; 
end_W(26, 184) <= 1; end_W(26, 185) <= 1; end_W(26, 186) <= 1; end_W(26, 187) <= 1; end_W(26, 188) <= 0; end_W(26, 189) <= 0; end_W(26, 190) <= 0; end_W(26, 191) <= 0; 
end_W(26, 192) <= 0; end_W(26, 193) <= 0; end_W(26, 194) <= 0; end_W(26, 195) <= 0; end_W(26, 196) <= 0; end_W(26, 197) <= 0; end_W(26, 198) <= 0; end_W(26, 199) <= 0; 
end_W(26, 200) <= 1; end_W(26, 201) <= 1; end_W(26, 202) <= 1; end_W(26, 203) <= 1; end_W(26, 204) <= 1; end_W(26, 205) <= 1; end_W(26, 206) <= 1; end_W(26, 207) <= 1; 
end_W(26, 208) <= 0; end_W(26, 209) <= 0; end_W(26, 210) <= 0; end_W(26, 211) <= 0; end_W(26, 212) <= 0; end_W(26, 213) <= 0; end_W(26, 214) <= 0; end_W(26, 215) <= 0; 
end_W(26, 216) <= 1; end_W(26, 217) <= 1; end_W(26, 218) <= 1; end_W(26, 219) <= 1; end_W(26, 220) <= 1; end_W(26, 221) <= 1; end_W(26, 222) <= 1; end_W(26, 223) <= 1; 
end_W(26, 224) <= 0; end_W(26, 225) <= 0; end_W(26, 226) <= 0; end_W(26, 227) <= 0; end_W(26, 228) <= 0; end_W(26, 229) <= 0; end_W(26, 230) <= 0; end_W(26, 231) <= 0; 
end_W(26, 232) <= 0; end_W(26, 233) <= 0; end_W(26, 234) <= 0; end_W(26, 235) <= 0; end_W(26, 236) <= 0; end_W(26, 237) <= 0; end_W(26, 238) <= 0; end_W(26, 239) <= 0; 
end_W(26, 240) <= 1; end_W(26, 241) <= 1; end_W(26, 242) <= 1; end_W(26, 243) <= 1; end_W(26, 244) <= 1; end_W(26, 245) <= 1; end_W(26, 246) <= 1; end_W(26, 247) <= 1; 
end_W(26, 248) <= 0; end_W(26, 249) <= 0; end_W(26, 250) <= 0; end_W(26, 251) <= 0; end_W(26, 252) <= 0; end_W(26, 253) <= 0; end_W(26, 254) <= 0; end_W(26, 255) <= 0; 
end_W(26, 256) <= 1; end_W(26, 257) <= 1; end_W(26, 258) <= 1; end_W(26, 259) <= 1; end_W(26, 260) <= 1; end_W(26, 261) <= 1; end_W(26, 262) <= 1; end_W(26, 263) <= 1; 
end_W(26, 264) <= 0; end_W(26, 265) <= 0; end_W(26, 266) <= 0; end_W(26, 267) <= 0; end_W(26, 268) <= 0; end_W(26, 269) <= 0; end_W(26, 270) <= 0; end_W(26, 271) <= 0; 
end_W(26, 272) <= 0; end_W(26, 273) <= 0; end_W(26, 274) <= 0; end_W(26, 275) <= 0; end_W(26, 276) <= 0; end_W(26, 277) <= 0; end_W(26, 278) <= 0; end_W(26, 279) <= 0; 
end_W(26, 280) <= 0; end_W(26, 281) <= 0; end_W(26, 282) <= 0; end_W(26, 283) <= 0; end_W(26, 284) <= 0; end_W(26, 285) <= 0; end_W(26, 286) <= 0; end_W(26, 287) <= 0; 
end_W(26, 288) <= 0; end_W(26, 289) <= 0; end_W(26, 290) <= 0; end_W(26, 291) <= 0; end_W(26, 292) <= 1; end_W(26, 293) <= 1; end_W(26, 294) <= 1; end_W(26, 295) <= 1; 
end_W(26, 296) <= 1; end_W(26, 297) <= 1; end_W(26, 298) <= 1; end_W(26, 299) <= 1; end_W(26, 300) <= 0; end_W(26, 301) <= 0; end_W(26, 302) <= 0; end_W(26, 303) <= 0; 
end_W(26, 304) <= 0; end_W(26, 305) <= 0; end_W(26, 306) <= 0; end_W(26, 307) <= 0; end_W(26, 308) <= 1; end_W(26, 309) <= 1; end_W(26, 310) <= 1; end_W(26, 311) <= 1; 
end_W(26, 312) <= 1; end_W(26, 313) <= 1; end_W(26, 314) <= 1; end_W(26, 315) <= 1; end_W(26, 316) <= 0; end_W(26, 317) <= 0; end_W(26, 318) <= 0; end_W(26, 319) <= 0; 
end_W(26, 320) <= 0; end_W(26, 321) <= 0; end_W(26, 322) <= 0; end_W(26, 323) <= 0; end_W(27, 0) <= 1; end_W(27, 1) <= 1; end_W(27, 2) <= 1; end_W(27, 3) <= 1; end_W(27, 4) <= 1; end_W(27, 5) <= 1; end_W(27, 6) <= 1; end_W(27, 7) <= 1; 
end_W(27, 8) <= 0; end_W(27, 9) <= 0; end_W(27, 10) <= 0; end_W(27, 11) <= 0; end_W(27, 12) <= 0; end_W(27, 13) <= 0; end_W(27, 14) <= 0; end_W(27, 15) <= 0; 
end_W(27, 16) <= 0; end_W(27, 17) <= 0; end_W(27, 18) <= 0; end_W(27, 19) <= 0; end_W(27, 20) <= 1; end_W(27, 21) <= 1; end_W(27, 22) <= 1; end_W(27, 23) <= 1; 
end_W(27, 24) <= 1; end_W(27, 25) <= 1; end_W(27, 26) <= 1; end_W(27, 27) <= 1; end_W(27, 28) <= 0; end_W(27, 29) <= 0; end_W(27, 30) <= 0; end_W(27, 31) <= 0; 
end_W(27, 32) <= 0; end_W(27, 33) <= 0; end_W(27, 34) <= 0; end_W(27, 35) <= 0; end_W(27, 36) <= 1; end_W(27, 37) <= 1; end_W(27, 38) <= 1; end_W(27, 39) <= 1; 
end_W(27, 40) <= 1; end_W(27, 41) <= 1; end_W(27, 42) <= 1; end_W(27, 43) <= 1; end_W(27, 44) <= 0; end_W(27, 45) <= 0; end_W(27, 46) <= 0; end_W(27, 47) <= 0; 
end_W(27, 48) <= 0; end_W(27, 49) <= 0; end_W(27, 50) <= 0; end_W(27, 51) <= 0; end_W(27, 52) <= 0; end_W(27, 53) <= 0; end_W(27, 54) <= 0; end_W(27, 55) <= 0; 
end_W(27, 56) <= 1; end_W(27, 57) <= 1; end_W(27, 58) <= 1; end_W(27, 59) <= 1; end_W(27, 60) <= 1; end_W(27, 61) <= 1; end_W(27, 62) <= 1; end_W(27, 63) <= 1; 
end_W(27, 64) <= 0; end_W(27, 65) <= 0; end_W(27, 66) <= 0; end_W(27, 67) <= 0; end_W(27, 68) <= 0; end_W(27, 69) <= 0; end_W(27, 70) <= 0; end_W(27, 71) <= 0; 
end_W(27, 72) <= 1; end_W(27, 73) <= 1; end_W(27, 74) <= 1; end_W(27, 75) <= 1; end_W(27, 76) <= 1; end_W(27, 77) <= 1; end_W(27, 78) <= 1; end_W(27, 79) <= 1; 
end_W(27, 80) <= 0; end_W(27, 81) <= 0; end_W(27, 82) <= 0; end_W(27, 83) <= 0; end_W(27, 84) <= 0; end_W(27, 85) <= 0; end_W(27, 86) <= 0; end_W(27, 87) <= 0; 
end_W(27, 88) <= 0; end_W(27, 89) <= 0; end_W(27, 90) <= 0; end_W(27, 91) <= 0; end_W(27, 92) <= 0; end_W(27, 93) <= 0; end_W(27, 94) <= 0; end_W(27, 95) <= 0; 
end_W(27, 96) <= 1; end_W(27, 97) <= 1; end_W(27, 98) <= 1; end_W(27, 99) <= 1; end_W(27, 100) <= 1; end_W(27, 101) <= 1; end_W(27, 102) <= 1; end_W(27, 103) <= 1; 
end_W(27, 104) <= 0; end_W(27, 105) <= 0; end_W(27, 106) <= 0; end_W(27, 107) <= 0; end_W(27, 108) <= 0; end_W(27, 109) <= 0; end_W(27, 110) <= 0; end_W(27, 111) <= 0; 
end_W(27, 112) <= 1; end_W(27, 113) <= 1; end_W(27, 114) <= 1; end_W(27, 115) <= 1; end_W(27, 116) <= 1; end_W(27, 117) <= 1; end_W(27, 118) <= 1; end_W(27, 119) <= 1; 
end_W(27, 120) <= 0; end_W(27, 121) <= 0; end_W(27, 122) <= 0; end_W(27, 123) <= 0; end_W(27, 124) <= 0; end_W(27, 125) <= 0; end_W(27, 126) <= 0; end_W(27, 127) <= 0; 
end_W(27, 128) <= 0; end_W(27, 129) <= 0; end_W(27, 130) <= 0; end_W(27, 131) <= 0; end_W(27, 132) <= 0; end_W(27, 133) <= 0; end_W(27, 134) <= 0; end_W(27, 135) <= 0; 
end_W(27, 136) <= 0; end_W(27, 137) <= 0; end_W(27, 138) <= 0; end_W(27, 139) <= 0; end_W(27, 140) <= 0; end_W(27, 141) <= 0; end_W(27, 142) <= 0; end_W(27, 143) <= 0; 
end_W(27, 144) <= 0; end_W(27, 145) <= 0; end_W(27, 146) <= 0; end_W(27, 147) <= 0; end_W(27, 148) <= 0; end_W(27, 149) <= 0; end_W(27, 150) <= 0; end_W(27, 151) <= 0; 
end_W(27, 152) <= 0; end_W(27, 153) <= 0; end_W(27, 154) <= 0; end_W(27, 155) <= 0; end_W(27, 156) <= 0; end_W(27, 157) <= 0; end_W(27, 158) <= 0; end_W(27, 159) <= 0; 
end_W(27, 160) <= 0; end_W(27, 161) <= 0; end_W(27, 162) <= 0; end_W(27, 163) <= 0; end_W(27, 164) <= 0; end_W(27, 165) <= 0; end_W(27, 166) <= 0; end_W(27, 167) <= 0; 
end_W(27, 168) <= 0; end_W(27, 169) <= 0; end_W(27, 170) <= 0; end_W(27, 171) <= 0; end_W(27, 172) <= 0; end_W(27, 173) <= 0; end_W(27, 174) <= 0; end_W(27, 175) <= 0; 
end_W(27, 176) <= 0; end_W(27, 177) <= 0; end_W(27, 178) <= 0; end_W(27, 179) <= 0; end_W(27, 180) <= 1; end_W(27, 181) <= 1; end_W(27, 182) <= 1; end_W(27, 183) <= 1; 
end_W(27, 184) <= 1; end_W(27, 185) <= 1; end_W(27, 186) <= 1; end_W(27, 187) <= 1; end_W(27, 188) <= 0; end_W(27, 189) <= 0; end_W(27, 190) <= 0; end_W(27, 191) <= 0; 
end_W(27, 192) <= 0; end_W(27, 193) <= 0; end_W(27, 194) <= 0; end_W(27, 195) <= 0; end_W(27, 196) <= 0; end_W(27, 197) <= 0; end_W(27, 198) <= 0; end_W(27, 199) <= 0; 
end_W(27, 200) <= 1; end_W(27, 201) <= 1; end_W(27, 202) <= 1; end_W(27, 203) <= 1; end_W(27, 204) <= 1; end_W(27, 205) <= 1; end_W(27, 206) <= 1; end_W(27, 207) <= 1; 
end_W(27, 208) <= 0; end_W(27, 209) <= 0; end_W(27, 210) <= 0; end_W(27, 211) <= 0; end_W(27, 212) <= 0; end_W(27, 213) <= 0; end_W(27, 214) <= 0; end_W(27, 215) <= 0; 
end_W(27, 216) <= 1; end_W(27, 217) <= 1; end_W(27, 218) <= 1; end_W(27, 219) <= 1; end_W(27, 220) <= 1; end_W(27, 221) <= 1; end_W(27, 222) <= 1; end_W(27, 223) <= 1; 
end_W(27, 224) <= 0; end_W(27, 225) <= 0; end_W(27, 226) <= 0; end_W(27, 227) <= 0; end_W(27, 228) <= 0; end_W(27, 229) <= 0; end_W(27, 230) <= 0; end_W(27, 231) <= 0; 
end_W(27, 232) <= 0; end_W(27, 233) <= 0; end_W(27, 234) <= 0; end_W(27, 235) <= 0; end_W(27, 236) <= 0; end_W(27, 237) <= 0; end_W(27, 238) <= 0; end_W(27, 239) <= 0; 
end_W(27, 240) <= 1; end_W(27, 241) <= 1; end_W(27, 242) <= 1; end_W(27, 243) <= 1; end_W(27, 244) <= 1; end_W(27, 245) <= 1; end_W(27, 246) <= 1; end_W(27, 247) <= 1; 
end_W(27, 248) <= 0; end_W(27, 249) <= 0; end_W(27, 250) <= 0; end_W(27, 251) <= 0; end_W(27, 252) <= 0; end_W(27, 253) <= 0; end_W(27, 254) <= 0; end_W(27, 255) <= 0; 
end_W(27, 256) <= 1; end_W(27, 257) <= 1; end_W(27, 258) <= 1; end_W(27, 259) <= 1; end_W(27, 260) <= 1; end_W(27, 261) <= 1; end_W(27, 262) <= 1; end_W(27, 263) <= 1; 
end_W(27, 264) <= 0; end_W(27, 265) <= 0; end_W(27, 266) <= 0; end_W(27, 267) <= 0; end_W(27, 268) <= 0; end_W(27, 269) <= 0; end_W(27, 270) <= 0; end_W(27, 271) <= 0; 
end_W(27, 272) <= 0; end_W(27, 273) <= 0; end_W(27, 274) <= 0; end_W(27, 275) <= 0; end_W(27, 276) <= 0; end_W(27, 277) <= 0; end_W(27, 278) <= 0; end_W(27, 279) <= 0; 
end_W(27, 280) <= 0; end_W(27, 281) <= 0; end_W(27, 282) <= 0; end_W(27, 283) <= 0; end_W(27, 284) <= 0; end_W(27, 285) <= 0; end_W(27, 286) <= 0; end_W(27, 287) <= 0; 
end_W(27, 288) <= 0; end_W(27, 289) <= 0; end_W(27, 290) <= 0; end_W(27, 291) <= 0; end_W(27, 292) <= 1; end_W(27, 293) <= 1; end_W(27, 294) <= 1; end_W(27, 295) <= 1; 
end_W(27, 296) <= 1; end_W(27, 297) <= 1; end_W(27, 298) <= 1; end_W(27, 299) <= 1; end_W(27, 300) <= 0; end_W(27, 301) <= 0; end_W(27, 302) <= 0; end_W(27, 303) <= 0; 
end_W(27, 304) <= 0; end_W(27, 305) <= 0; end_W(27, 306) <= 0; end_W(27, 307) <= 0; end_W(27, 308) <= 1; end_W(27, 309) <= 1; end_W(27, 310) <= 1; end_W(27, 311) <= 1; 
end_W(27, 312) <= 1; end_W(27, 313) <= 1; end_W(27, 314) <= 1; end_W(27, 315) <= 1; end_W(27, 316) <= 0; end_W(27, 317) <= 0; end_W(27, 318) <= 0; end_W(27, 319) <= 0; 
end_W(27, 320) <= 0; end_W(27, 321) <= 0; end_W(27, 322) <= 0; end_W(27, 323) <= 0; end_W(28, 0) <= 1; end_W(28, 1) <= 1; end_W(28, 2) <= 1; end_W(28, 3) <= 1; end_W(28, 4) <= 1; end_W(28, 5) <= 1; end_W(28, 6) <= 1; end_W(28, 7) <= 1; 
end_W(28, 8) <= 0; end_W(28, 9) <= 0; end_W(28, 10) <= 0; end_W(28, 11) <= 0; end_W(28, 12) <= 0; end_W(28, 13) <= 0; end_W(28, 14) <= 0; end_W(28, 15) <= 0; 
end_W(28, 16) <= 0; end_W(28, 17) <= 0; end_W(28, 18) <= 0; end_W(28, 19) <= 0; end_W(28, 20) <= 1; end_W(28, 21) <= 1; end_W(28, 22) <= 1; end_W(28, 23) <= 1; 
end_W(28, 24) <= 1; end_W(28, 25) <= 1; end_W(28, 26) <= 1; end_W(28, 27) <= 1; end_W(28, 28) <= 0; end_W(28, 29) <= 0; end_W(28, 30) <= 0; end_W(28, 31) <= 0; 
end_W(28, 32) <= 0; end_W(28, 33) <= 0; end_W(28, 34) <= 0; end_W(28, 35) <= 0; end_W(28, 36) <= 1; end_W(28, 37) <= 1; end_W(28, 38) <= 1; end_W(28, 39) <= 1; 
end_W(28, 40) <= 1; end_W(28, 41) <= 1; end_W(28, 42) <= 1; end_W(28, 43) <= 1; end_W(28, 44) <= 0; end_W(28, 45) <= 0; end_W(28, 46) <= 0; end_W(28, 47) <= 0; 
end_W(28, 48) <= 0; end_W(28, 49) <= 0; end_W(28, 50) <= 0; end_W(28, 51) <= 0; end_W(28, 52) <= 0; end_W(28, 53) <= 0; end_W(28, 54) <= 0; end_W(28, 55) <= 0; 
end_W(28, 56) <= 1; end_W(28, 57) <= 1; end_W(28, 58) <= 1; end_W(28, 59) <= 1; end_W(28, 60) <= 1; end_W(28, 61) <= 1; end_W(28, 62) <= 1; end_W(28, 63) <= 1; 
end_W(28, 64) <= 0; end_W(28, 65) <= 0; end_W(28, 66) <= 0; end_W(28, 67) <= 0; end_W(28, 68) <= 0; end_W(28, 69) <= 0; end_W(28, 70) <= 0; end_W(28, 71) <= 0; 
end_W(28, 72) <= 1; end_W(28, 73) <= 1; end_W(28, 74) <= 1; end_W(28, 75) <= 1; end_W(28, 76) <= 1; end_W(28, 77) <= 1; end_W(28, 78) <= 1; end_W(28, 79) <= 1; 
end_W(28, 80) <= 0; end_W(28, 81) <= 0; end_W(28, 82) <= 0; end_W(28, 83) <= 0; end_W(28, 84) <= 0; end_W(28, 85) <= 0; end_W(28, 86) <= 0; end_W(28, 87) <= 0; 
end_W(28, 88) <= 0; end_W(28, 89) <= 0; end_W(28, 90) <= 0; end_W(28, 91) <= 0; end_W(28, 92) <= 0; end_W(28, 93) <= 0; end_W(28, 94) <= 0; end_W(28, 95) <= 0; 
end_W(28, 96) <= 1; end_W(28, 97) <= 1; end_W(28, 98) <= 1; end_W(28, 99) <= 1; end_W(28, 100) <= 1; end_W(28, 101) <= 1; end_W(28, 102) <= 1; end_W(28, 103) <= 1; 
end_W(28, 104) <= 0; end_W(28, 105) <= 0; end_W(28, 106) <= 0; end_W(28, 107) <= 0; end_W(28, 108) <= 0; end_W(28, 109) <= 0; end_W(28, 110) <= 0; end_W(28, 111) <= 0; 
end_W(28, 112) <= 1; end_W(28, 113) <= 1; end_W(28, 114) <= 1; end_W(28, 115) <= 1; end_W(28, 116) <= 1; end_W(28, 117) <= 1; end_W(28, 118) <= 1; end_W(28, 119) <= 1; 
end_W(28, 120) <= 0; end_W(28, 121) <= 0; end_W(28, 122) <= 0; end_W(28, 123) <= 0; end_W(28, 124) <= 0; end_W(28, 125) <= 0; end_W(28, 126) <= 0; end_W(28, 127) <= 0; 
end_W(28, 128) <= 0; end_W(28, 129) <= 0; end_W(28, 130) <= 0; end_W(28, 131) <= 0; end_W(28, 132) <= 1; end_W(28, 133) <= 1; end_W(28, 134) <= 1; end_W(28, 135) <= 1; 
end_W(28, 136) <= 0; end_W(28, 137) <= 0; end_W(28, 138) <= 0; end_W(28, 139) <= 0; end_W(28, 140) <= 0; end_W(28, 141) <= 0; end_W(28, 142) <= 0; end_W(28, 143) <= 0; 
end_W(28, 144) <= 0; end_W(28, 145) <= 0; end_W(28, 146) <= 0; end_W(28, 147) <= 0; end_W(28, 148) <= 0; end_W(28, 149) <= 0; end_W(28, 150) <= 0; end_W(28, 151) <= 0; 
end_W(28, 152) <= 0; end_W(28, 153) <= 0; end_W(28, 154) <= 0; end_W(28, 155) <= 0; end_W(28, 156) <= 0; end_W(28, 157) <= 0; end_W(28, 158) <= 0; end_W(28, 159) <= 0; 
end_W(28, 160) <= 0; end_W(28, 161) <= 0; end_W(28, 162) <= 0; end_W(28, 163) <= 0; end_W(28, 164) <= 0; end_W(28, 165) <= 0; end_W(28, 166) <= 0; end_W(28, 167) <= 0; 
end_W(28, 168) <= 0; end_W(28, 169) <= 0; end_W(28, 170) <= 0; end_W(28, 171) <= 0; end_W(28, 172) <= 0; end_W(28, 173) <= 0; end_W(28, 174) <= 0; end_W(28, 175) <= 0; 
end_W(28, 176) <= 0; end_W(28, 177) <= 0; end_W(28, 178) <= 0; end_W(28, 179) <= 0; end_W(28, 180) <= 1; end_W(28, 181) <= 1; end_W(28, 182) <= 1; end_W(28, 183) <= 1; 
end_W(28, 184) <= 1; end_W(28, 185) <= 1; end_W(28, 186) <= 1; end_W(28, 187) <= 1; end_W(28, 188) <= 0; end_W(28, 189) <= 0; end_W(28, 190) <= 0; end_W(28, 191) <= 0; 
end_W(28, 192) <= 0; end_W(28, 193) <= 0; end_W(28, 194) <= 0; end_W(28, 195) <= 0; end_W(28, 196) <= 0; end_W(28, 197) <= 0; end_W(28, 198) <= 0; end_W(28, 199) <= 0; 
end_W(28, 200) <= 1; end_W(28, 201) <= 1; end_W(28, 202) <= 1; end_W(28, 203) <= 1; end_W(28, 204) <= 1; end_W(28, 205) <= 1; end_W(28, 206) <= 1; end_W(28, 207) <= 1; 
end_W(28, 208) <= 0; end_W(28, 209) <= 0; end_W(28, 210) <= 0; end_W(28, 211) <= 0; end_W(28, 212) <= 0; end_W(28, 213) <= 0; end_W(28, 214) <= 0; end_W(28, 215) <= 0; 
end_W(28, 216) <= 0; end_W(28, 217) <= 0; end_W(28, 218) <= 0; end_W(28, 219) <= 0; end_W(28, 220) <= 1; end_W(28, 221) <= 1; end_W(28, 222) <= 1; end_W(28, 223) <= 1; 
end_W(28, 224) <= 1; end_W(28, 225) <= 1; end_W(28, 226) <= 1; end_W(28, 227) <= 1; end_W(28, 228) <= 0; end_W(28, 229) <= 0; end_W(28, 230) <= 0; end_W(28, 231) <= 0; 
end_W(28, 232) <= 0; end_W(28, 233) <= 0; end_W(28, 234) <= 0; end_W(28, 235) <= 0; end_W(28, 236) <= 1; end_W(28, 237) <= 1; end_W(28, 238) <= 1; end_W(28, 239) <= 1; 
end_W(28, 240) <= 1; end_W(28, 241) <= 1; end_W(28, 242) <= 1; end_W(28, 243) <= 1; end_W(28, 244) <= 0; end_W(28, 245) <= 0; end_W(28, 246) <= 0; end_W(28, 247) <= 0; 
end_W(28, 248) <= 0; end_W(28, 249) <= 0; end_W(28, 250) <= 0; end_W(28, 251) <= 0; end_W(28, 252) <= 0; end_W(28, 253) <= 0; end_W(28, 254) <= 0; end_W(28, 255) <= 0; 
end_W(28, 256) <= 1; end_W(28, 257) <= 1; end_W(28, 258) <= 1; end_W(28, 259) <= 1; end_W(28, 260) <= 1; end_W(28, 261) <= 1; end_W(28, 262) <= 1; end_W(28, 263) <= 1; 
end_W(28, 264) <= 0; end_W(28, 265) <= 0; end_W(28, 266) <= 0; end_W(28, 267) <= 0; end_W(28, 268) <= 0; end_W(28, 269) <= 0; end_W(28, 270) <= 0; end_W(28, 271) <= 0; 
end_W(28, 272) <= 0; end_W(28, 273) <= 0; end_W(28, 274) <= 0; end_W(28, 275) <= 0; end_W(28, 276) <= 1; end_W(28, 277) <= 1; end_W(28, 278) <= 1; end_W(28, 279) <= 1; 
end_W(28, 280) <= 0; end_W(28, 281) <= 0; end_W(28, 282) <= 0; end_W(28, 283) <= 0; end_W(28, 284) <= 0; end_W(28, 285) <= 0; end_W(28, 286) <= 0; end_W(28, 287) <= 0; 
end_W(28, 288) <= 0; end_W(28, 289) <= 0; end_W(28, 290) <= 0; end_W(28, 291) <= 0; end_W(28, 292) <= 1; end_W(28, 293) <= 1; end_W(28, 294) <= 1; end_W(28, 295) <= 1; 
end_W(28, 296) <= 1; end_W(28, 297) <= 1; end_W(28, 298) <= 1; end_W(28, 299) <= 1; end_W(28, 300) <= 0; end_W(28, 301) <= 0; end_W(28, 302) <= 0; end_W(28, 303) <= 0; 
end_W(28, 304) <= 0; end_W(28, 305) <= 0; end_W(28, 306) <= 0; end_W(28, 307) <= 0; end_W(28, 308) <= 1; end_W(28, 309) <= 1; end_W(28, 310) <= 1; end_W(28, 311) <= 1; 
end_W(28, 312) <= 1; end_W(28, 313) <= 1; end_W(28, 314) <= 1; end_W(28, 315) <= 1; end_W(28, 316) <= 0; end_W(28, 317) <= 0; end_W(28, 318) <= 0; end_W(28, 319) <= 0; 
end_W(28, 320) <= 0; end_W(28, 321) <= 0; end_W(28, 322) <= 0; end_W(28, 323) <= 0; end_W(29, 0) <= 1; end_W(29, 1) <= 1; end_W(29, 2) <= 1; end_W(29, 3) <= 1; end_W(29, 4) <= 1; end_W(29, 5) <= 1; end_W(29, 6) <= 1; end_W(29, 7) <= 1; 
end_W(29, 8) <= 0; end_W(29, 9) <= 0; end_W(29, 10) <= 0; end_W(29, 11) <= 0; end_W(29, 12) <= 0; end_W(29, 13) <= 0; end_W(29, 14) <= 0; end_W(29, 15) <= 0; 
end_W(29, 16) <= 0; end_W(29, 17) <= 0; end_W(29, 18) <= 0; end_W(29, 19) <= 0; end_W(29, 20) <= 1; end_W(29, 21) <= 1; end_W(29, 22) <= 1; end_W(29, 23) <= 1; 
end_W(29, 24) <= 1; end_W(29, 25) <= 1; end_W(29, 26) <= 1; end_W(29, 27) <= 1; end_W(29, 28) <= 0; end_W(29, 29) <= 0; end_W(29, 30) <= 0; end_W(29, 31) <= 0; 
end_W(29, 32) <= 0; end_W(29, 33) <= 0; end_W(29, 34) <= 0; end_W(29, 35) <= 0; end_W(29, 36) <= 1; end_W(29, 37) <= 1; end_W(29, 38) <= 1; end_W(29, 39) <= 1; 
end_W(29, 40) <= 1; end_W(29, 41) <= 1; end_W(29, 42) <= 1; end_W(29, 43) <= 1; end_W(29, 44) <= 0; end_W(29, 45) <= 0; end_W(29, 46) <= 0; end_W(29, 47) <= 0; 
end_W(29, 48) <= 0; end_W(29, 49) <= 0; end_W(29, 50) <= 0; end_W(29, 51) <= 0; end_W(29, 52) <= 0; end_W(29, 53) <= 0; end_W(29, 54) <= 0; end_W(29, 55) <= 0; 
end_W(29, 56) <= 1; end_W(29, 57) <= 1; end_W(29, 58) <= 1; end_W(29, 59) <= 1; end_W(29, 60) <= 1; end_W(29, 61) <= 1; end_W(29, 62) <= 1; end_W(29, 63) <= 1; 
end_W(29, 64) <= 0; end_W(29, 65) <= 0; end_W(29, 66) <= 0; end_W(29, 67) <= 0; end_W(29, 68) <= 0; end_W(29, 69) <= 0; end_W(29, 70) <= 0; end_W(29, 71) <= 0; 
end_W(29, 72) <= 1; end_W(29, 73) <= 1; end_W(29, 74) <= 1; end_W(29, 75) <= 1; end_W(29, 76) <= 1; end_W(29, 77) <= 1; end_W(29, 78) <= 1; end_W(29, 79) <= 1; 
end_W(29, 80) <= 0; end_W(29, 81) <= 0; end_W(29, 82) <= 0; end_W(29, 83) <= 0; end_W(29, 84) <= 0; end_W(29, 85) <= 0; end_W(29, 86) <= 0; end_W(29, 87) <= 0; 
end_W(29, 88) <= 0; end_W(29, 89) <= 0; end_W(29, 90) <= 0; end_W(29, 91) <= 0; end_W(29, 92) <= 0; end_W(29, 93) <= 0; end_W(29, 94) <= 0; end_W(29, 95) <= 0; 
end_W(29, 96) <= 1; end_W(29, 97) <= 1; end_W(29, 98) <= 1; end_W(29, 99) <= 1; end_W(29, 100) <= 1; end_W(29, 101) <= 1; end_W(29, 102) <= 1; end_W(29, 103) <= 1; 
end_W(29, 104) <= 0; end_W(29, 105) <= 0; end_W(29, 106) <= 0; end_W(29, 107) <= 0; end_W(29, 108) <= 0; end_W(29, 109) <= 0; end_W(29, 110) <= 0; end_W(29, 111) <= 0; 
end_W(29, 112) <= 1; end_W(29, 113) <= 1; end_W(29, 114) <= 1; end_W(29, 115) <= 1; end_W(29, 116) <= 1; end_W(29, 117) <= 1; end_W(29, 118) <= 1; end_W(29, 119) <= 1; 
end_W(29, 120) <= 0; end_W(29, 121) <= 0; end_W(29, 122) <= 0; end_W(29, 123) <= 0; end_W(29, 124) <= 0; end_W(29, 125) <= 0; end_W(29, 126) <= 0; end_W(29, 127) <= 0; 
end_W(29, 128) <= 0; end_W(29, 129) <= 0; end_W(29, 130) <= 0; end_W(29, 131) <= 0; end_W(29, 132) <= 1; end_W(29, 133) <= 1; end_W(29, 134) <= 1; end_W(29, 135) <= 1; 
end_W(29, 136) <= 0; end_W(29, 137) <= 0; end_W(29, 138) <= 0; end_W(29, 139) <= 0; end_W(29, 140) <= 0; end_W(29, 141) <= 0; end_W(29, 142) <= 0; end_W(29, 143) <= 0; 
end_W(29, 144) <= 0; end_W(29, 145) <= 0; end_W(29, 146) <= 0; end_W(29, 147) <= 0; end_W(29, 148) <= 0; end_W(29, 149) <= 0; end_W(29, 150) <= 0; end_W(29, 151) <= 0; 
end_W(29, 152) <= 0; end_W(29, 153) <= 0; end_W(29, 154) <= 0; end_W(29, 155) <= 0; end_W(29, 156) <= 0; end_W(29, 157) <= 0; end_W(29, 158) <= 0; end_W(29, 159) <= 0; 
end_W(29, 160) <= 0; end_W(29, 161) <= 0; end_W(29, 162) <= 0; end_W(29, 163) <= 0; end_W(29, 164) <= 0; end_W(29, 165) <= 0; end_W(29, 166) <= 0; end_W(29, 167) <= 0; 
end_W(29, 168) <= 0; end_W(29, 169) <= 0; end_W(29, 170) <= 0; end_W(29, 171) <= 0; end_W(29, 172) <= 0; end_W(29, 173) <= 0; end_W(29, 174) <= 0; end_W(29, 175) <= 0; 
end_W(29, 176) <= 0; end_W(29, 177) <= 0; end_W(29, 178) <= 0; end_W(29, 179) <= 0; end_W(29, 180) <= 1; end_W(29, 181) <= 1; end_W(29, 182) <= 1; end_W(29, 183) <= 1; 
end_W(29, 184) <= 1; end_W(29, 185) <= 1; end_W(29, 186) <= 1; end_W(29, 187) <= 1; end_W(29, 188) <= 0; end_W(29, 189) <= 0; end_W(29, 190) <= 0; end_W(29, 191) <= 0; 
end_W(29, 192) <= 0; end_W(29, 193) <= 0; end_W(29, 194) <= 0; end_W(29, 195) <= 0; end_W(29, 196) <= 0; end_W(29, 197) <= 0; end_W(29, 198) <= 0; end_W(29, 199) <= 0; 
end_W(29, 200) <= 1; end_W(29, 201) <= 1; end_W(29, 202) <= 1; end_W(29, 203) <= 1; end_W(29, 204) <= 1; end_W(29, 205) <= 1; end_W(29, 206) <= 1; end_W(29, 207) <= 1; 
end_W(29, 208) <= 0; end_W(29, 209) <= 0; end_W(29, 210) <= 0; end_W(29, 211) <= 0; end_W(29, 212) <= 0; end_W(29, 213) <= 0; end_W(29, 214) <= 0; end_W(29, 215) <= 0; 
end_W(29, 216) <= 0; end_W(29, 217) <= 0; end_W(29, 218) <= 0; end_W(29, 219) <= 0; end_W(29, 220) <= 1; end_W(29, 221) <= 1; end_W(29, 222) <= 1; end_W(29, 223) <= 1; 
end_W(29, 224) <= 1; end_W(29, 225) <= 1; end_W(29, 226) <= 1; end_W(29, 227) <= 1; end_W(29, 228) <= 0; end_W(29, 229) <= 0; end_W(29, 230) <= 0; end_W(29, 231) <= 0; 
end_W(29, 232) <= 0; end_W(29, 233) <= 0; end_W(29, 234) <= 0; end_W(29, 235) <= 0; end_W(29, 236) <= 1; end_W(29, 237) <= 1; end_W(29, 238) <= 1; end_W(29, 239) <= 1; 
end_W(29, 240) <= 1; end_W(29, 241) <= 1; end_W(29, 242) <= 1; end_W(29, 243) <= 1; end_W(29, 244) <= 0; end_W(29, 245) <= 0; end_W(29, 246) <= 0; end_W(29, 247) <= 0; 
end_W(29, 248) <= 0; end_W(29, 249) <= 0; end_W(29, 250) <= 0; end_W(29, 251) <= 0; end_W(29, 252) <= 0; end_W(29, 253) <= 0; end_W(29, 254) <= 0; end_W(29, 255) <= 0; 
end_W(29, 256) <= 1; end_W(29, 257) <= 1; end_W(29, 258) <= 1; end_W(29, 259) <= 1; end_W(29, 260) <= 1; end_W(29, 261) <= 1; end_W(29, 262) <= 1; end_W(29, 263) <= 1; 
end_W(29, 264) <= 0; end_W(29, 265) <= 0; end_W(29, 266) <= 0; end_W(29, 267) <= 0; end_W(29, 268) <= 0; end_W(29, 269) <= 0; end_W(29, 270) <= 0; end_W(29, 271) <= 0; 
end_W(29, 272) <= 0; end_W(29, 273) <= 0; end_W(29, 274) <= 0; end_W(29, 275) <= 0; end_W(29, 276) <= 1; end_W(29, 277) <= 1; end_W(29, 278) <= 1; end_W(29, 279) <= 1; 
end_W(29, 280) <= 0; end_W(29, 281) <= 0; end_W(29, 282) <= 0; end_W(29, 283) <= 0; end_W(29, 284) <= 0; end_W(29, 285) <= 0; end_W(29, 286) <= 0; end_W(29, 287) <= 0; 
end_W(29, 288) <= 0; end_W(29, 289) <= 0; end_W(29, 290) <= 0; end_W(29, 291) <= 0; end_W(29, 292) <= 1; end_W(29, 293) <= 1; end_W(29, 294) <= 1; end_W(29, 295) <= 1; 
end_W(29, 296) <= 1; end_W(29, 297) <= 1; end_W(29, 298) <= 1; end_W(29, 299) <= 1; end_W(29, 300) <= 0; end_W(29, 301) <= 0; end_W(29, 302) <= 0; end_W(29, 303) <= 0; 
end_W(29, 304) <= 0; end_W(29, 305) <= 0; end_W(29, 306) <= 0; end_W(29, 307) <= 0; end_W(29, 308) <= 1; end_W(29, 309) <= 1; end_W(29, 310) <= 1; end_W(29, 311) <= 1; 
end_W(29, 312) <= 1; end_W(29, 313) <= 1; end_W(29, 314) <= 1; end_W(29, 315) <= 1; end_W(29, 316) <= 0; end_W(29, 317) <= 0; end_W(29, 318) <= 0; end_W(29, 319) <= 0; 
end_W(29, 320) <= 0; end_W(29, 321) <= 0; end_W(29, 322) <= 0; end_W(29, 323) <= 0; end_W(30, 0) <= 1; end_W(30, 1) <= 1; end_W(30, 2) <= 1; end_W(30, 3) <= 1; end_W(30, 4) <= 1; end_W(30, 5) <= 1; end_W(30, 6) <= 1; end_W(30, 7) <= 1; 
end_W(30, 8) <= 0; end_W(30, 9) <= 0; end_W(30, 10) <= 0; end_W(30, 11) <= 0; end_W(30, 12) <= 0; end_W(30, 13) <= 0; end_W(30, 14) <= 0; end_W(30, 15) <= 0; 
end_W(30, 16) <= 0; end_W(30, 17) <= 0; end_W(30, 18) <= 0; end_W(30, 19) <= 0; end_W(30, 20) <= 1; end_W(30, 21) <= 1; end_W(30, 22) <= 1; end_W(30, 23) <= 1; 
end_W(30, 24) <= 1; end_W(30, 25) <= 1; end_W(30, 26) <= 1; end_W(30, 27) <= 1; end_W(30, 28) <= 0; end_W(30, 29) <= 0; end_W(30, 30) <= 0; end_W(30, 31) <= 0; 
end_W(30, 32) <= 0; end_W(30, 33) <= 0; end_W(30, 34) <= 0; end_W(30, 35) <= 0; end_W(30, 36) <= 1; end_W(30, 37) <= 1; end_W(30, 38) <= 1; end_W(30, 39) <= 1; 
end_W(30, 40) <= 1; end_W(30, 41) <= 1; end_W(30, 42) <= 1; end_W(30, 43) <= 1; end_W(30, 44) <= 0; end_W(30, 45) <= 0; end_W(30, 46) <= 0; end_W(30, 47) <= 0; 
end_W(30, 48) <= 0; end_W(30, 49) <= 0; end_W(30, 50) <= 0; end_W(30, 51) <= 0; end_W(30, 52) <= 0; end_W(30, 53) <= 0; end_W(30, 54) <= 0; end_W(30, 55) <= 0; 
end_W(30, 56) <= 1; end_W(30, 57) <= 1; end_W(30, 58) <= 1; end_W(30, 59) <= 1; end_W(30, 60) <= 1; end_W(30, 61) <= 1; end_W(30, 62) <= 1; end_W(30, 63) <= 1; 
end_W(30, 64) <= 0; end_W(30, 65) <= 0; end_W(30, 66) <= 0; end_W(30, 67) <= 0; end_W(30, 68) <= 0; end_W(30, 69) <= 0; end_W(30, 70) <= 0; end_W(30, 71) <= 0; 
end_W(30, 72) <= 1; end_W(30, 73) <= 1; end_W(30, 74) <= 1; end_W(30, 75) <= 1; end_W(30, 76) <= 1; end_W(30, 77) <= 1; end_W(30, 78) <= 1; end_W(30, 79) <= 1; 
end_W(30, 80) <= 0; end_W(30, 81) <= 0; end_W(30, 82) <= 0; end_W(30, 83) <= 0; end_W(30, 84) <= 0; end_W(30, 85) <= 0; end_W(30, 86) <= 0; end_W(30, 87) <= 0; 
end_W(30, 88) <= 0; end_W(30, 89) <= 0; end_W(30, 90) <= 0; end_W(30, 91) <= 0; end_W(30, 92) <= 0; end_W(30, 93) <= 0; end_W(30, 94) <= 0; end_W(30, 95) <= 0; 
end_W(30, 96) <= 1; end_W(30, 97) <= 1; end_W(30, 98) <= 1; end_W(30, 99) <= 1; end_W(30, 100) <= 1; end_W(30, 101) <= 1; end_W(30, 102) <= 1; end_W(30, 103) <= 1; 
end_W(30, 104) <= 0; end_W(30, 105) <= 0; end_W(30, 106) <= 0; end_W(30, 107) <= 0; end_W(30, 108) <= 0; end_W(30, 109) <= 0; end_W(30, 110) <= 0; end_W(30, 111) <= 0; 
end_W(30, 112) <= 1; end_W(30, 113) <= 1; end_W(30, 114) <= 1; end_W(30, 115) <= 1; end_W(30, 116) <= 1; end_W(30, 117) <= 1; end_W(30, 118) <= 1; end_W(30, 119) <= 1; 
end_W(30, 120) <= 0; end_W(30, 121) <= 0; end_W(30, 122) <= 0; end_W(30, 123) <= 0; end_W(30, 124) <= 0; end_W(30, 125) <= 0; end_W(30, 126) <= 0; end_W(30, 127) <= 0; 
end_W(30, 128) <= 0; end_W(30, 129) <= 0; end_W(30, 130) <= 0; end_W(30, 131) <= 0; end_W(30, 132) <= 1; end_W(30, 133) <= 1; end_W(30, 134) <= 1; end_W(30, 135) <= 1; 
end_W(30, 136) <= 0; end_W(30, 137) <= 0; end_W(30, 138) <= 0; end_W(30, 139) <= 0; end_W(30, 140) <= 0; end_W(30, 141) <= 0; end_W(30, 142) <= 0; end_W(30, 143) <= 0; 
end_W(30, 144) <= 0; end_W(30, 145) <= 0; end_W(30, 146) <= 0; end_W(30, 147) <= 0; end_W(30, 148) <= 0; end_W(30, 149) <= 0; end_W(30, 150) <= 0; end_W(30, 151) <= 0; 
end_W(30, 152) <= 0; end_W(30, 153) <= 0; end_W(30, 154) <= 0; end_W(30, 155) <= 0; end_W(30, 156) <= 0; end_W(30, 157) <= 0; end_W(30, 158) <= 0; end_W(30, 159) <= 0; 
end_W(30, 160) <= 0; end_W(30, 161) <= 0; end_W(30, 162) <= 0; end_W(30, 163) <= 0; end_W(30, 164) <= 0; end_W(30, 165) <= 0; end_W(30, 166) <= 0; end_W(30, 167) <= 0; 
end_W(30, 168) <= 0; end_W(30, 169) <= 0; end_W(30, 170) <= 0; end_W(30, 171) <= 0; end_W(30, 172) <= 0; end_W(30, 173) <= 0; end_W(30, 174) <= 0; end_W(30, 175) <= 0; 
end_W(30, 176) <= 0; end_W(30, 177) <= 0; end_W(30, 178) <= 0; end_W(30, 179) <= 0; end_W(30, 180) <= 1; end_W(30, 181) <= 1; end_W(30, 182) <= 1; end_W(30, 183) <= 1; 
end_W(30, 184) <= 1; end_W(30, 185) <= 1; end_W(30, 186) <= 1; end_W(30, 187) <= 1; end_W(30, 188) <= 0; end_W(30, 189) <= 0; end_W(30, 190) <= 0; end_W(30, 191) <= 0; 
end_W(30, 192) <= 0; end_W(30, 193) <= 0; end_W(30, 194) <= 0; end_W(30, 195) <= 0; end_W(30, 196) <= 0; end_W(30, 197) <= 0; end_W(30, 198) <= 0; end_W(30, 199) <= 0; 
end_W(30, 200) <= 1; end_W(30, 201) <= 1; end_W(30, 202) <= 1; end_W(30, 203) <= 1; end_W(30, 204) <= 1; end_W(30, 205) <= 1; end_W(30, 206) <= 1; end_W(30, 207) <= 1; 
end_W(30, 208) <= 0; end_W(30, 209) <= 0; end_W(30, 210) <= 0; end_W(30, 211) <= 0; end_W(30, 212) <= 0; end_W(30, 213) <= 0; end_W(30, 214) <= 0; end_W(30, 215) <= 0; 
end_W(30, 216) <= 0; end_W(30, 217) <= 0; end_W(30, 218) <= 0; end_W(30, 219) <= 0; end_W(30, 220) <= 1; end_W(30, 221) <= 1; end_W(30, 222) <= 1; end_W(30, 223) <= 1; 
end_W(30, 224) <= 1; end_W(30, 225) <= 1; end_W(30, 226) <= 1; end_W(30, 227) <= 1; end_W(30, 228) <= 0; end_W(30, 229) <= 0; end_W(30, 230) <= 0; end_W(30, 231) <= 0; 
end_W(30, 232) <= 0; end_W(30, 233) <= 0; end_W(30, 234) <= 0; end_W(30, 235) <= 0; end_W(30, 236) <= 1; end_W(30, 237) <= 1; end_W(30, 238) <= 1; end_W(30, 239) <= 1; 
end_W(30, 240) <= 1; end_W(30, 241) <= 1; end_W(30, 242) <= 1; end_W(30, 243) <= 1; end_W(30, 244) <= 0; end_W(30, 245) <= 0; end_W(30, 246) <= 0; end_W(30, 247) <= 0; 
end_W(30, 248) <= 0; end_W(30, 249) <= 0; end_W(30, 250) <= 0; end_W(30, 251) <= 0; end_W(30, 252) <= 0; end_W(30, 253) <= 0; end_W(30, 254) <= 0; end_W(30, 255) <= 0; 
end_W(30, 256) <= 1; end_W(30, 257) <= 1; end_W(30, 258) <= 1; end_W(30, 259) <= 1; end_W(30, 260) <= 1; end_W(30, 261) <= 1; end_W(30, 262) <= 1; end_W(30, 263) <= 1; 
end_W(30, 264) <= 0; end_W(30, 265) <= 0; end_W(30, 266) <= 0; end_W(30, 267) <= 0; end_W(30, 268) <= 0; end_W(30, 269) <= 0; end_W(30, 270) <= 0; end_W(30, 271) <= 0; 
end_W(30, 272) <= 0; end_W(30, 273) <= 0; end_W(30, 274) <= 0; end_W(30, 275) <= 0; end_W(30, 276) <= 1; end_W(30, 277) <= 1; end_W(30, 278) <= 1; end_W(30, 279) <= 1; 
end_W(30, 280) <= 0; end_W(30, 281) <= 0; end_W(30, 282) <= 0; end_W(30, 283) <= 0; end_W(30, 284) <= 0; end_W(30, 285) <= 0; end_W(30, 286) <= 0; end_W(30, 287) <= 0; 
end_W(30, 288) <= 0; end_W(30, 289) <= 0; end_W(30, 290) <= 0; end_W(30, 291) <= 0; end_W(30, 292) <= 1; end_W(30, 293) <= 1; end_W(30, 294) <= 1; end_W(30, 295) <= 1; 
end_W(30, 296) <= 1; end_W(30, 297) <= 1; end_W(30, 298) <= 1; end_W(30, 299) <= 1; end_W(30, 300) <= 0; end_W(30, 301) <= 0; end_W(30, 302) <= 0; end_W(30, 303) <= 0; 
end_W(30, 304) <= 0; end_W(30, 305) <= 0; end_W(30, 306) <= 0; end_W(30, 307) <= 0; end_W(30, 308) <= 1; end_W(30, 309) <= 1; end_W(30, 310) <= 1; end_W(30, 311) <= 1; 
end_W(30, 312) <= 1; end_W(30, 313) <= 1; end_W(30, 314) <= 1; end_W(30, 315) <= 1; end_W(30, 316) <= 0; end_W(30, 317) <= 0; end_W(30, 318) <= 0; end_W(30, 319) <= 0; 
end_W(30, 320) <= 0; end_W(30, 321) <= 0; end_W(30, 322) <= 0; end_W(30, 323) <= 0; end_W(31, 0) <= 1; end_W(31, 1) <= 1; end_W(31, 2) <= 1; end_W(31, 3) <= 1; end_W(31, 4) <= 1; end_W(31, 5) <= 1; end_W(31, 6) <= 1; end_W(31, 7) <= 1; 
end_W(31, 8) <= 0; end_W(31, 9) <= 0; end_W(31, 10) <= 0; end_W(31, 11) <= 0; end_W(31, 12) <= 0; end_W(31, 13) <= 0; end_W(31, 14) <= 0; end_W(31, 15) <= 0; 
end_W(31, 16) <= 0; end_W(31, 17) <= 0; end_W(31, 18) <= 0; end_W(31, 19) <= 0; end_W(31, 20) <= 1; end_W(31, 21) <= 1; end_W(31, 22) <= 1; end_W(31, 23) <= 1; 
end_W(31, 24) <= 1; end_W(31, 25) <= 1; end_W(31, 26) <= 1; end_W(31, 27) <= 1; end_W(31, 28) <= 0; end_W(31, 29) <= 0; end_W(31, 30) <= 0; end_W(31, 31) <= 0; 
end_W(31, 32) <= 0; end_W(31, 33) <= 0; end_W(31, 34) <= 0; end_W(31, 35) <= 0; end_W(31, 36) <= 1; end_W(31, 37) <= 1; end_W(31, 38) <= 1; end_W(31, 39) <= 1; 
end_W(31, 40) <= 1; end_W(31, 41) <= 1; end_W(31, 42) <= 1; end_W(31, 43) <= 1; end_W(31, 44) <= 0; end_W(31, 45) <= 0; end_W(31, 46) <= 0; end_W(31, 47) <= 0; 
end_W(31, 48) <= 0; end_W(31, 49) <= 0; end_W(31, 50) <= 0; end_W(31, 51) <= 0; end_W(31, 52) <= 0; end_W(31, 53) <= 0; end_W(31, 54) <= 0; end_W(31, 55) <= 0; 
end_W(31, 56) <= 1; end_W(31, 57) <= 1; end_W(31, 58) <= 1; end_W(31, 59) <= 1; end_W(31, 60) <= 1; end_W(31, 61) <= 1; end_W(31, 62) <= 1; end_W(31, 63) <= 1; 
end_W(31, 64) <= 0; end_W(31, 65) <= 0; end_W(31, 66) <= 0; end_W(31, 67) <= 0; end_W(31, 68) <= 0; end_W(31, 69) <= 0; end_W(31, 70) <= 0; end_W(31, 71) <= 0; 
end_W(31, 72) <= 1; end_W(31, 73) <= 1; end_W(31, 74) <= 1; end_W(31, 75) <= 1; end_W(31, 76) <= 1; end_W(31, 77) <= 1; end_W(31, 78) <= 1; end_W(31, 79) <= 1; 
end_W(31, 80) <= 0; end_W(31, 81) <= 0; end_W(31, 82) <= 0; end_W(31, 83) <= 0; end_W(31, 84) <= 0; end_W(31, 85) <= 0; end_W(31, 86) <= 0; end_W(31, 87) <= 0; 
end_W(31, 88) <= 0; end_W(31, 89) <= 0; end_W(31, 90) <= 0; end_W(31, 91) <= 0; end_W(31, 92) <= 0; end_W(31, 93) <= 0; end_W(31, 94) <= 0; end_W(31, 95) <= 0; 
end_W(31, 96) <= 1; end_W(31, 97) <= 1; end_W(31, 98) <= 1; end_W(31, 99) <= 1; end_W(31, 100) <= 1; end_W(31, 101) <= 1; end_W(31, 102) <= 1; end_W(31, 103) <= 1; 
end_W(31, 104) <= 0; end_W(31, 105) <= 0; end_W(31, 106) <= 0; end_W(31, 107) <= 0; end_W(31, 108) <= 0; end_W(31, 109) <= 0; end_W(31, 110) <= 0; end_W(31, 111) <= 0; 
end_W(31, 112) <= 1; end_W(31, 113) <= 1; end_W(31, 114) <= 1; end_W(31, 115) <= 1; end_W(31, 116) <= 1; end_W(31, 117) <= 1; end_W(31, 118) <= 1; end_W(31, 119) <= 1; 
end_W(31, 120) <= 0; end_W(31, 121) <= 0; end_W(31, 122) <= 0; end_W(31, 123) <= 0; end_W(31, 124) <= 0; end_W(31, 125) <= 0; end_W(31, 126) <= 0; end_W(31, 127) <= 0; 
end_W(31, 128) <= 0; end_W(31, 129) <= 0; end_W(31, 130) <= 0; end_W(31, 131) <= 0; end_W(31, 132) <= 1; end_W(31, 133) <= 1; end_W(31, 134) <= 1; end_W(31, 135) <= 1; 
end_W(31, 136) <= 0; end_W(31, 137) <= 0; end_W(31, 138) <= 0; end_W(31, 139) <= 0; end_W(31, 140) <= 0; end_W(31, 141) <= 0; end_W(31, 142) <= 0; end_W(31, 143) <= 0; 
end_W(31, 144) <= 0; end_W(31, 145) <= 0; end_W(31, 146) <= 0; end_W(31, 147) <= 0; end_W(31, 148) <= 0; end_W(31, 149) <= 0; end_W(31, 150) <= 0; end_W(31, 151) <= 0; 
end_W(31, 152) <= 0; end_W(31, 153) <= 0; end_W(31, 154) <= 0; end_W(31, 155) <= 0; end_W(31, 156) <= 0; end_W(31, 157) <= 0; end_W(31, 158) <= 0; end_W(31, 159) <= 0; 
end_W(31, 160) <= 0; end_W(31, 161) <= 0; end_W(31, 162) <= 0; end_W(31, 163) <= 0; end_W(31, 164) <= 0; end_W(31, 165) <= 0; end_W(31, 166) <= 0; end_W(31, 167) <= 0; 
end_W(31, 168) <= 0; end_W(31, 169) <= 0; end_W(31, 170) <= 0; end_W(31, 171) <= 0; end_W(31, 172) <= 0; end_W(31, 173) <= 0; end_W(31, 174) <= 0; end_W(31, 175) <= 0; 
end_W(31, 176) <= 0; end_W(31, 177) <= 0; end_W(31, 178) <= 0; end_W(31, 179) <= 0; end_W(31, 180) <= 1; end_W(31, 181) <= 1; end_W(31, 182) <= 1; end_W(31, 183) <= 1; 
end_W(31, 184) <= 1; end_W(31, 185) <= 1; end_W(31, 186) <= 1; end_W(31, 187) <= 1; end_W(31, 188) <= 0; end_W(31, 189) <= 0; end_W(31, 190) <= 0; end_W(31, 191) <= 0; 
end_W(31, 192) <= 0; end_W(31, 193) <= 0; end_W(31, 194) <= 0; end_W(31, 195) <= 0; end_W(31, 196) <= 0; end_W(31, 197) <= 0; end_W(31, 198) <= 0; end_W(31, 199) <= 0; 
end_W(31, 200) <= 1; end_W(31, 201) <= 1; end_W(31, 202) <= 1; end_W(31, 203) <= 1; end_W(31, 204) <= 1; end_W(31, 205) <= 1; end_W(31, 206) <= 1; end_W(31, 207) <= 1; 
end_W(31, 208) <= 0; end_W(31, 209) <= 0; end_W(31, 210) <= 0; end_W(31, 211) <= 0; end_W(31, 212) <= 0; end_W(31, 213) <= 0; end_W(31, 214) <= 0; end_W(31, 215) <= 0; 
end_W(31, 216) <= 0; end_W(31, 217) <= 0; end_W(31, 218) <= 0; end_W(31, 219) <= 0; end_W(31, 220) <= 1; end_W(31, 221) <= 1; end_W(31, 222) <= 1; end_W(31, 223) <= 1; 
end_W(31, 224) <= 1; end_W(31, 225) <= 1; end_W(31, 226) <= 1; end_W(31, 227) <= 1; end_W(31, 228) <= 0; end_W(31, 229) <= 0; end_W(31, 230) <= 0; end_W(31, 231) <= 0; 
end_W(31, 232) <= 0; end_W(31, 233) <= 0; end_W(31, 234) <= 0; end_W(31, 235) <= 0; end_W(31, 236) <= 1; end_W(31, 237) <= 1; end_W(31, 238) <= 1; end_W(31, 239) <= 1; 
end_W(31, 240) <= 1; end_W(31, 241) <= 1; end_W(31, 242) <= 1; end_W(31, 243) <= 1; end_W(31, 244) <= 0; end_W(31, 245) <= 0; end_W(31, 246) <= 0; end_W(31, 247) <= 0; 
end_W(31, 248) <= 0; end_W(31, 249) <= 0; end_W(31, 250) <= 0; end_W(31, 251) <= 0; end_W(31, 252) <= 0; end_W(31, 253) <= 0; end_W(31, 254) <= 0; end_W(31, 255) <= 0; 
end_W(31, 256) <= 1; end_W(31, 257) <= 1; end_W(31, 258) <= 1; end_W(31, 259) <= 1; end_W(31, 260) <= 1; end_W(31, 261) <= 1; end_W(31, 262) <= 1; end_W(31, 263) <= 1; 
end_W(31, 264) <= 0; end_W(31, 265) <= 0; end_W(31, 266) <= 0; end_W(31, 267) <= 0; end_W(31, 268) <= 0; end_W(31, 269) <= 0; end_W(31, 270) <= 0; end_W(31, 271) <= 0; 
end_W(31, 272) <= 0; end_W(31, 273) <= 0; end_W(31, 274) <= 0; end_W(31, 275) <= 0; end_W(31, 276) <= 1; end_W(31, 277) <= 1; end_W(31, 278) <= 1; end_W(31, 279) <= 1; 
end_W(31, 280) <= 0; end_W(31, 281) <= 0; end_W(31, 282) <= 0; end_W(31, 283) <= 0; end_W(31, 284) <= 0; end_W(31, 285) <= 0; end_W(31, 286) <= 0; end_W(31, 287) <= 0; 
end_W(31, 288) <= 0; end_W(31, 289) <= 0; end_W(31, 290) <= 0; end_W(31, 291) <= 0; end_W(31, 292) <= 1; end_W(31, 293) <= 1; end_W(31, 294) <= 1; end_W(31, 295) <= 1; 
end_W(31, 296) <= 1; end_W(31, 297) <= 1; end_W(31, 298) <= 1; end_W(31, 299) <= 1; end_W(31, 300) <= 0; end_W(31, 301) <= 0; end_W(31, 302) <= 0; end_W(31, 303) <= 0; 
end_W(31, 304) <= 0; end_W(31, 305) <= 0; end_W(31, 306) <= 0; end_W(31, 307) <= 0; end_W(31, 308) <= 1; end_W(31, 309) <= 1; end_W(31, 310) <= 1; end_W(31, 311) <= 1; 
end_W(31, 312) <= 1; end_W(31, 313) <= 1; end_W(31, 314) <= 1; end_W(31, 315) <= 1; end_W(31, 316) <= 0; end_W(31, 317) <= 0; end_W(31, 318) <= 0; end_W(31, 319) <= 0; 
end_W(31, 320) <= 0; end_W(31, 321) <= 0; end_W(31, 322) <= 0; end_W(31, 323) <= 0; end_W(32, 0) <= 0; end_W(32, 1) <= 0; end_W(32, 2) <= 0; end_W(32, 3) <= 0; end_W(32, 4) <= 1; end_W(32, 5) <= 1; end_W(32, 6) <= 1; end_W(32, 7) <= 1; 
end_W(32, 8) <= 1; end_W(32, 9) <= 1; end_W(32, 10) <= 1; end_W(32, 11) <= 1; end_W(32, 12) <= 0; end_W(32, 13) <= 0; end_W(32, 14) <= 0; end_W(32, 15) <= 0; 
end_W(32, 16) <= 0; end_W(32, 17) <= 0; end_W(32, 18) <= 0; end_W(32, 19) <= 0; end_W(32, 20) <= 1; end_W(32, 21) <= 1; end_W(32, 22) <= 1; end_W(32, 23) <= 1; 
end_W(32, 24) <= 1; end_W(32, 25) <= 1; end_W(32, 26) <= 1; end_W(32, 27) <= 1; end_W(32, 28) <= 0; end_W(32, 29) <= 0; end_W(32, 30) <= 0; end_W(32, 31) <= 0; 
end_W(32, 32) <= 0; end_W(32, 33) <= 0; end_W(32, 34) <= 0; end_W(32, 35) <= 0; end_W(32, 36) <= 1; end_W(32, 37) <= 1; end_W(32, 38) <= 1; end_W(32, 39) <= 1; 
end_W(32, 40) <= 1; end_W(32, 41) <= 1; end_W(32, 42) <= 1; end_W(32, 43) <= 1; end_W(32, 44) <= 0; end_W(32, 45) <= 0; end_W(32, 46) <= 0; end_W(32, 47) <= 0; 
end_W(32, 48) <= 0; end_W(32, 49) <= 0; end_W(32, 50) <= 0; end_W(32, 51) <= 0; end_W(32, 52) <= 0; end_W(32, 53) <= 0; end_W(32, 54) <= 0; end_W(32, 55) <= 0; 
end_W(32, 56) <= 1; end_W(32, 57) <= 1; end_W(32, 58) <= 1; end_W(32, 59) <= 1; end_W(32, 60) <= 1; end_W(32, 61) <= 1; end_W(32, 62) <= 1; end_W(32, 63) <= 1; 
end_W(32, 64) <= 0; end_W(32, 65) <= 0; end_W(32, 66) <= 0; end_W(32, 67) <= 0; end_W(32, 68) <= 0; end_W(32, 69) <= 0; end_W(32, 70) <= 0; end_W(32, 71) <= 0; 
end_W(32, 72) <= 1; end_W(32, 73) <= 1; end_W(32, 74) <= 1; end_W(32, 75) <= 1; end_W(32, 76) <= 1; end_W(32, 77) <= 1; end_W(32, 78) <= 1; end_W(32, 79) <= 1; 
end_W(32, 80) <= 0; end_W(32, 81) <= 0; end_W(32, 82) <= 0; end_W(32, 83) <= 0; end_W(32, 84) <= 0; end_W(32, 85) <= 0; end_W(32, 86) <= 0; end_W(32, 87) <= 0; 
end_W(32, 88) <= 0; end_W(32, 89) <= 0; end_W(32, 90) <= 0; end_W(32, 91) <= 0; end_W(32, 92) <= 0; end_W(32, 93) <= 0; end_W(32, 94) <= 0; end_W(32, 95) <= 0; 
end_W(32, 96) <= 1; end_W(32, 97) <= 1; end_W(32, 98) <= 1; end_W(32, 99) <= 1; end_W(32, 100) <= 1; end_W(32, 101) <= 1; end_W(32, 102) <= 1; end_W(32, 103) <= 1; 
end_W(32, 104) <= 0; end_W(32, 105) <= 0; end_W(32, 106) <= 0; end_W(32, 107) <= 0; end_W(32, 108) <= 0; end_W(32, 109) <= 0; end_W(32, 110) <= 0; end_W(32, 111) <= 0; 
end_W(32, 112) <= 1; end_W(32, 113) <= 1; end_W(32, 114) <= 1; end_W(32, 115) <= 1; end_W(32, 116) <= 1; end_W(32, 117) <= 1; end_W(32, 118) <= 1; end_W(32, 119) <= 1; 
end_W(32, 120) <= 0; end_W(32, 121) <= 0; end_W(32, 122) <= 0; end_W(32, 123) <= 0; end_W(32, 124) <= 0; end_W(32, 125) <= 0; end_W(32, 126) <= 0; end_W(32, 127) <= 0; 
end_W(32, 128) <= 1; end_W(32, 129) <= 1; end_W(32, 130) <= 1; end_W(32, 131) <= 1; end_W(32, 132) <= 1; end_W(32, 133) <= 1; end_W(32, 134) <= 1; end_W(32, 135) <= 1; 
end_W(32, 136) <= 0; end_W(32, 137) <= 0; end_W(32, 138) <= 0; end_W(32, 139) <= 0; end_W(32, 140) <= 0; end_W(32, 141) <= 0; end_W(32, 142) <= 0; end_W(32, 143) <= 0; 
end_W(32, 144) <= 0; end_W(32, 145) <= 0; end_W(32, 146) <= 0; end_W(32, 147) <= 0; end_W(32, 148) <= 0; end_W(32, 149) <= 0; end_W(32, 150) <= 0; end_W(32, 151) <= 0; 
end_W(32, 152) <= 0; end_W(32, 153) <= 0; end_W(32, 154) <= 0; end_W(32, 155) <= 0; end_W(32, 156) <= 0; end_W(32, 157) <= 0; end_W(32, 158) <= 0; end_W(32, 159) <= 0; 
end_W(32, 160) <= 0; end_W(32, 161) <= 0; end_W(32, 162) <= 0; end_W(32, 163) <= 0; end_W(32, 164) <= 0; end_W(32, 165) <= 0; end_W(32, 166) <= 0; end_W(32, 167) <= 0; 
end_W(32, 168) <= 0; end_W(32, 169) <= 0; end_W(32, 170) <= 0; end_W(32, 171) <= 0; end_W(32, 172) <= 0; end_W(32, 173) <= 0; end_W(32, 174) <= 0; end_W(32, 175) <= 0; 
end_W(32, 176) <= 0; end_W(32, 177) <= 0; end_W(32, 178) <= 0; end_W(32, 179) <= 0; end_W(32, 180) <= 1; end_W(32, 181) <= 1; end_W(32, 182) <= 1; end_W(32, 183) <= 1; 
end_W(32, 184) <= 1; end_W(32, 185) <= 1; end_W(32, 186) <= 1; end_W(32, 187) <= 1; end_W(32, 188) <= 0; end_W(32, 189) <= 0; end_W(32, 190) <= 0; end_W(32, 191) <= 0; 
end_W(32, 192) <= 0; end_W(32, 193) <= 0; end_W(32, 194) <= 0; end_W(32, 195) <= 0; end_W(32, 196) <= 0; end_W(32, 197) <= 0; end_W(32, 198) <= 0; end_W(32, 199) <= 0; 
end_W(32, 200) <= 1; end_W(32, 201) <= 1; end_W(32, 202) <= 1; end_W(32, 203) <= 1; end_W(32, 204) <= 1; end_W(32, 205) <= 1; end_W(32, 206) <= 1; end_W(32, 207) <= 1; 
end_W(32, 208) <= 0; end_W(32, 209) <= 0; end_W(32, 210) <= 0; end_W(32, 211) <= 0; end_W(32, 212) <= 0; end_W(32, 213) <= 0; end_W(32, 214) <= 0; end_W(32, 215) <= 0; 
end_W(32, 216) <= 0; end_W(32, 217) <= 0; end_W(32, 218) <= 0; end_W(32, 219) <= 0; end_W(32, 220) <= 0; end_W(32, 221) <= 0; end_W(32, 222) <= 0; end_W(32, 223) <= 0; 
end_W(32, 224) <= 1; end_W(32, 225) <= 1; end_W(32, 226) <= 1; end_W(32, 227) <= 1; end_W(32, 228) <= 1; end_W(32, 229) <= 1; end_W(32, 230) <= 1; end_W(32, 231) <= 1; 
end_W(32, 232) <= 1; end_W(32, 233) <= 1; end_W(32, 234) <= 1; end_W(32, 235) <= 1; end_W(32, 236) <= 1; end_W(32, 237) <= 1; end_W(32, 238) <= 1; end_W(32, 239) <= 1; 
end_W(32, 240) <= 0; end_W(32, 241) <= 0; end_W(32, 242) <= 0; end_W(32, 243) <= 0; end_W(32, 244) <= 0; end_W(32, 245) <= 0; end_W(32, 246) <= 0; end_W(32, 247) <= 0; 
end_W(32, 248) <= 0; end_W(32, 249) <= 0; end_W(32, 250) <= 0; end_W(32, 251) <= 0; end_W(32, 252) <= 0; end_W(32, 253) <= 0; end_W(32, 254) <= 0; end_W(32, 255) <= 0; 
end_W(32, 256) <= 1; end_W(32, 257) <= 1; end_W(32, 258) <= 1; end_W(32, 259) <= 1; end_W(32, 260) <= 1; end_W(32, 261) <= 1; end_W(32, 262) <= 1; end_W(32, 263) <= 1; 
end_W(32, 264) <= 0; end_W(32, 265) <= 0; end_W(32, 266) <= 0; end_W(32, 267) <= 0; end_W(32, 268) <= 0; end_W(32, 269) <= 0; end_W(32, 270) <= 0; end_W(32, 271) <= 0; 
end_W(32, 272) <= 1; end_W(32, 273) <= 1; end_W(32, 274) <= 1; end_W(32, 275) <= 1; end_W(32, 276) <= 1; end_W(32, 277) <= 1; end_W(32, 278) <= 1; end_W(32, 279) <= 1; 
end_W(32, 280) <= 0; end_W(32, 281) <= 0; end_W(32, 282) <= 0; end_W(32, 283) <= 0; end_W(32, 284) <= 0; end_W(32, 285) <= 0; end_W(32, 286) <= 0; end_W(32, 287) <= 0; 
end_W(32, 288) <= 0; end_W(32, 289) <= 0; end_W(32, 290) <= 0; end_W(32, 291) <= 0; end_W(32, 292) <= 1; end_W(32, 293) <= 1; end_W(32, 294) <= 1; end_W(32, 295) <= 1; 
end_W(32, 296) <= 1; end_W(32, 297) <= 1; end_W(32, 298) <= 1; end_W(32, 299) <= 1; end_W(32, 300) <= 0; end_W(32, 301) <= 0; end_W(32, 302) <= 0; end_W(32, 303) <= 0; 
end_W(32, 304) <= 0; end_W(32, 305) <= 0; end_W(32, 306) <= 0; end_W(32, 307) <= 0; end_W(32, 308) <= 1; end_W(32, 309) <= 1; end_W(32, 310) <= 1; end_W(32, 311) <= 1; 
end_W(32, 312) <= 1; end_W(32, 313) <= 1; end_W(32, 314) <= 1; end_W(32, 315) <= 1; end_W(32, 316) <= 0; end_W(32, 317) <= 0; end_W(32, 318) <= 0; end_W(32, 319) <= 0; 
end_W(32, 320) <= 0; end_W(32, 321) <= 0; end_W(32, 322) <= 0; end_W(32, 323) <= 0; end_W(33, 0) <= 0; end_W(33, 1) <= 0; end_W(33, 2) <= 0; end_W(33, 3) <= 0; end_W(33, 4) <= 1; end_W(33, 5) <= 1; end_W(33, 6) <= 1; end_W(33, 7) <= 1; 
end_W(33, 8) <= 1; end_W(33, 9) <= 1; end_W(33, 10) <= 1; end_W(33, 11) <= 1; end_W(33, 12) <= 0; end_W(33, 13) <= 0; end_W(33, 14) <= 0; end_W(33, 15) <= 0; 
end_W(33, 16) <= 0; end_W(33, 17) <= 0; end_W(33, 18) <= 0; end_W(33, 19) <= 0; end_W(33, 20) <= 1; end_W(33, 21) <= 1; end_W(33, 22) <= 1; end_W(33, 23) <= 1; 
end_W(33, 24) <= 1; end_W(33, 25) <= 1; end_W(33, 26) <= 1; end_W(33, 27) <= 1; end_W(33, 28) <= 0; end_W(33, 29) <= 0; end_W(33, 30) <= 0; end_W(33, 31) <= 0; 
end_W(33, 32) <= 0; end_W(33, 33) <= 0; end_W(33, 34) <= 0; end_W(33, 35) <= 0; end_W(33, 36) <= 1; end_W(33, 37) <= 1; end_W(33, 38) <= 1; end_W(33, 39) <= 1; 
end_W(33, 40) <= 1; end_W(33, 41) <= 1; end_W(33, 42) <= 1; end_W(33, 43) <= 1; end_W(33, 44) <= 0; end_W(33, 45) <= 0; end_W(33, 46) <= 0; end_W(33, 47) <= 0; 
end_W(33, 48) <= 0; end_W(33, 49) <= 0; end_W(33, 50) <= 0; end_W(33, 51) <= 0; end_W(33, 52) <= 0; end_W(33, 53) <= 0; end_W(33, 54) <= 0; end_W(33, 55) <= 0; 
end_W(33, 56) <= 1; end_W(33, 57) <= 1; end_W(33, 58) <= 1; end_W(33, 59) <= 1; end_W(33, 60) <= 1; end_W(33, 61) <= 1; end_W(33, 62) <= 1; end_W(33, 63) <= 1; 
end_W(33, 64) <= 0; end_W(33, 65) <= 0; end_W(33, 66) <= 0; end_W(33, 67) <= 0; end_W(33, 68) <= 0; end_W(33, 69) <= 0; end_W(33, 70) <= 0; end_W(33, 71) <= 0; 
end_W(33, 72) <= 1; end_W(33, 73) <= 1; end_W(33, 74) <= 1; end_W(33, 75) <= 1; end_W(33, 76) <= 1; end_W(33, 77) <= 1; end_W(33, 78) <= 1; end_W(33, 79) <= 1; 
end_W(33, 80) <= 0; end_W(33, 81) <= 0; end_W(33, 82) <= 0; end_W(33, 83) <= 0; end_W(33, 84) <= 0; end_W(33, 85) <= 0; end_W(33, 86) <= 0; end_W(33, 87) <= 0; 
end_W(33, 88) <= 0; end_W(33, 89) <= 0; end_W(33, 90) <= 0; end_W(33, 91) <= 0; end_W(33, 92) <= 0; end_W(33, 93) <= 0; end_W(33, 94) <= 0; end_W(33, 95) <= 0; 
end_W(33, 96) <= 1; end_W(33, 97) <= 1; end_W(33, 98) <= 1; end_W(33, 99) <= 1; end_W(33, 100) <= 1; end_W(33, 101) <= 1; end_W(33, 102) <= 1; end_W(33, 103) <= 1; 
end_W(33, 104) <= 0; end_W(33, 105) <= 0; end_W(33, 106) <= 0; end_W(33, 107) <= 0; end_W(33, 108) <= 0; end_W(33, 109) <= 0; end_W(33, 110) <= 0; end_W(33, 111) <= 0; 
end_W(33, 112) <= 1; end_W(33, 113) <= 1; end_W(33, 114) <= 1; end_W(33, 115) <= 1; end_W(33, 116) <= 1; end_W(33, 117) <= 1; end_W(33, 118) <= 1; end_W(33, 119) <= 1; 
end_W(33, 120) <= 0; end_W(33, 121) <= 0; end_W(33, 122) <= 0; end_W(33, 123) <= 0; end_W(33, 124) <= 0; end_W(33, 125) <= 0; end_W(33, 126) <= 0; end_W(33, 127) <= 0; 
end_W(33, 128) <= 1; end_W(33, 129) <= 1; end_W(33, 130) <= 1; end_W(33, 131) <= 1; end_W(33, 132) <= 1; end_W(33, 133) <= 1; end_W(33, 134) <= 1; end_W(33, 135) <= 1; 
end_W(33, 136) <= 0; end_W(33, 137) <= 0; end_W(33, 138) <= 0; end_W(33, 139) <= 0; end_W(33, 140) <= 0; end_W(33, 141) <= 0; end_W(33, 142) <= 0; end_W(33, 143) <= 0; 
end_W(33, 144) <= 0; end_W(33, 145) <= 0; end_W(33, 146) <= 0; end_W(33, 147) <= 0; end_W(33, 148) <= 0; end_W(33, 149) <= 0; end_W(33, 150) <= 0; end_W(33, 151) <= 0; 
end_W(33, 152) <= 0; end_W(33, 153) <= 0; end_W(33, 154) <= 0; end_W(33, 155) <= 0; end_W(33, 156) <= 0; end_W(33, 157) <= 0; end_W(33, 158) <= 0; end_W(33, 159) <= 0; 
end_W(33, 160) <= 0; end_W(33, 161) <= 0; end_W(33, 162) <= 0; end_W(33, 163) <= 0; end_W(33, 164) <= 0; end_W(33, 165) <= 0; end_W(33, 166) <= 0; end_W(33, 167) <= 0; 
end_W(33, 168) <= 0; end_W(33, 169) <= 0; end_W(33, 170) <= 0; end_W(33, 171) <= 0; end_W(33, 172) <= 0; end_W(33, 173) <= 0; end_W(33, 174) <= 0; end_W(33, 175) <= 0; 
end_W(33, 176) <= 0; end_W(33, 177) <= 0; end_W(33, 178) <= 0; end_W(33, 179) <= 0; end_W(33, 180) <= 1; end_W(33, 181) <= 1; end_W(33, 182) <= 1; end_W(33, 183) <= 1; 
end_W(33, 184) <= 1; end_W(33, 185) <= 1; end_W(33, 186) <= 1; end_W(33, 187) <= 1; end_W(33, 188) <= 0; end_W(33, 189) <= 0; end_W(33, 190) <= 0; end_W(33, 191) <= 0; 
end_W(33, 192) <= 0; end_W(33, 193) <= 0; end_W(33, 194) <= 0; end_W(33, 195) <= 0; end_W(33, 196) <= 0; end_W(33, 197) <= 0; end_W(33, 198) <= 0; end_W(33, 199) <= 0; 
end_W(33, 200) <= 1; end_W(33, 201) <= 1; end_W(33, 202) <= 1; end_W(33, 203) <= 1; end_W(33, 204) <= 1; end_W(33, 205) <= 1; end_W(33, 206) <= 1; end_W(33, 207) <= 1; 
end_W(33, 208) <= 0; end_W(33, 209) <= 0; end_W(33, 210) <= 0; end_W(33, 211) <= 0; end_W(33, 212) <= 0; end_W(33, 213) <= 0; end_W(33, 214) <= 0; end_W(33, 215) <= 0; 
end_W(33, 216) <= 0; end_W(33, 217) <= 0; end_W(33, 218) <= 0; end_W(33, 219) <= 0; end_W(33, 220) <= 0; end_W(33, 221) <= 0; end_W(33, 222) <= 0; end_W(33, 223) <= 0; 
end_W(33, 224) <= 1; end_W(33, 225) <= 1; end_W(33, 226) <= 1; end_W(33, 227) <= 1; end_W(33, 228) <= 1; end_W(33, 229) <= 1; end_W(33, 230) <= 1; end_W(33, 231) <= 1; 
end_W(33, 232) <= 1; end_W(33, 233) <= 1; end_W(33, 234) <= 1; end_W(33, 235) <= 1; end_W(33, 236) <= 1; end_W(33, 237) <= 1; end_W(33, 238) <= 1; end_W(33, 239) <= 1; 
end_W(33, 240) <= 0; end_W(33, 241) <= 0; end_W(33, 242) <= 0; end_W(33, 243) <= 0; end_W(33, 244) <= 0; end_W(33, 245) <= 0; end_W(33, 246) <= 0; end_W(33, 247) <= 0; 
end_W(33, 248) <= 0; end_W(33, 249) <= 0; end_W(33, 250) <= 0; end_W(33, 251) <= 0; end_W(33, 252) <= 0; end_W(33, 253) <= 0; end_W(33, 254) <= 0; end_W(33, 255) <= 0; 
end_W(33, 256) <= 1; end_W(33, 257) <= 1; end_W(33, 258) <= 1; end_W(33, 259) <= 1; end_W(33, 260) <= 1; end_W(33, 261) <= 1; end_W(33, 262) <= 1; end_W(33, 263) <= 1; 
end_W(33, 264) <= 0; end_W(33, 265) <= 0; end_W(33, 266) <= 0; end_W(33, 267) <= 0; end_W(33, 268) <= 0; end_W(33, 269) <= 0; end_W(33, 270) <= 0; end_W(33, 271) <= 0; 
end_W(33, 272) <= 1; end_W(33, 273) <= 1; end_W(33, 274) <= 1; end_W(33, 275) <= 1; end_W(33, 276) <= 1; end_W(33, 277) <= 1; end_W(33, 278) <= 1; end_W(33, 279) <= 1; 
end_W(33, 280) <= 0; end_W(33, 281) <= 0; end_W(33, 282) <= 0; end_W(33, 283) <= 0; end_W(33, 284) <= 0; end_W(33, 285) <= 0; end_W(33, 286) <= 0; end_W(33, 287) <= 0; 
end_W(33, 288) <= 0; end_W(33, 289) <= 0; end_W(33, 290) <= 0; end_W(33, 291) <= 0; end_W(33, 292) <= 1; end_W(33, 293) <= 1; end_W(33, 294) <= 1; end_W(33, 295) <= 1; 
end_W(33, 296) <= 1; end_W(33, 297) <= 1; end_W(33, 298) <= 1; end_W(33, 299) <= 1; end_W(33, 300) <= 0; end_W(33, 301) <= 0; end_W(33, 302) <= 0; end_W(33, 303) <= 0; 
end_W(33, 304) <= 0; end_W(33, 305) <= 0; end_W(33, 306) <= 0; end_W(33, 307) <= 0; end_W(33, 308) <= 1; end_W(33, 309) <= 1; end_W(33, 310) <= 1; end_W(33, 311) <= 1; 
end_W(33, 312) <= 1; end_W(33, 313) <= 1; end_W(33, 314) <= 1; end_W(33, 315) <= 1; end_W(33, 316) <= 0; end_W(33, 317) <= 0; end_W(33, 318) <= 0; end_W(33, 319) <= 0; 
end_W(33, 320) <= 0; end_W(33, 321) <= 0; end_W(33, 322) <= 0; end_W(33, 323) <= 0; end_W(34, 0) <= 0; end_W(34, 1) <= 0; end_W(34, 2) <= 0; end_W(34, 3) <= 0; end_W(34, 4) <= 1; end_W(34, 5) <= 1; end_W(34, 6) <= 1; end_W(34, 7) <= 1; 
end_W(34, 8) <= 1; end_W(34, 9) <= 1; end_W(34, 10) <= 1; end_W(34, 11) <= 1; end_W(34, 12) <= 0; end_W(34, 13) <= 0; end_W(34, 14) <= 0; end_W(34, 15) <= 0; 
end_W(34, 16) <= 0; end_W(34, 17) <= 0; end_W(34, 18) <= 0; end_W(34, 19) <= 0; end_W(34, 20) <= 1; end_W(34, 21) <= 1; end_W(34, 22) <= 1; end_W(34, 23) <= 1; 
end_W(34, 24) <= 1; end_W(34, 25) <= 1; end_W(34, 26) <= 1; end_W(34, 27) <= 1; end_W(34, 28) <= 0; end_W(34, 29) <= 0; end_W(34, 30) <= 0; end_W(34, 31) <= 0; 
end_W(34, 32) <= 0; end_W(34, 33) <= 0; end_W(34, 34) <= 0; end_W(34, 35) <= 0; end_W(34, 36) <= 1; end_W(34, 37) <= 1; end_W(34, 38) <= 1; end_W(34, 39) <= 1; 
end_W(34, 40) <= 1; end_W(34, 41) <= 1; end_W(34, 42) <= 1; end_W(34, 43) <= 1; end_W(34, 44) <= 0; end_W(34, 45) <= 0; end_W(34, 46) <= 0; end_W(34, 47) <= 0; 
end_W(34, 48) <= 0; end_W(34, 49) <= 0; end_W(34, 50) <= 0; end_W(34, 51) <= 0; end_W(34, 52) <= 0; end_W(34, 53) <= 0; end_W(34, 54) <= 0; end_W(34, 55) <= 0; 
end_W(34, 56) <= 1; end_W(34, 57) <= 1; end_W(34, 58) <= 1; end_W(34, 59) <= 1; end_W(34, 60) <= 1; end_W(34, 61) <= 1; end_W(34, 62) <= 1; end_W(34, 63) <= 1; 
end_W(34, 64) <= 0; end_W(34, 65) <= 0; end_W(34, 66) <= 0; end_W(34, 67) <= 0; end_W(34, 68) <= 0; end_W(34, 69) <= 0; end_W(34, 70) <= 0; end_W(34, 71) <= 0; 
end_W(34, 72) <= 1; end_W(34, 73) <= 1; end_W(34, 74) <= 1; end_W(34, 75) <= 1; end_W(34, 76) <= 1; end_W(34, 77) <= 1; end_W(34, 78) <= 1; end_W(34, 79) <= 1; 
end_W(34, 80) <= 0; end_W(34, 81) <= 0; end_W(34, 82) <= 0; end_W(34, 83) <= 0; end_W(34, 84) <= 0; end_W(34, 85) <= 0; end_W(34, 86) <= 0; end_W(34, 87) <= 0; 
end_W(34, 88) <= 0; end_W(34, 89) <= 0; end_W(34, 90) <= 0; end_W(34, 91) <= 0; end_W(34, 92) <= 0; end_W(34, 93) <= 0; end_W(34, 94) <= 0; end_W(34, 95) <= 0; 
end_W(34, 96) <= 1; end_W(34, 97) <= 1; end_W(34, 98) <= 1; end_W(34, 99) <= 1; end_W(34, 100) <= 1; end_W(34, 101) <= 1; end_W(34, 102) <= 1; end_W(34, 103) <= 1; 
end_W(34, 104) <= 0; end_W(34, 105) <= 0; end_W(34, 106) <= 0; end_W(34, 107) <= 0; end_W(34, 108) <= 0; end_W(34, 109) <= 0; end_W(34, 110) <= 0; end_W(34, 111) <= 0; 
end_W(34, 112) <= 1; end_W(34, 113) <= 1; end_W(34, 114) <= 1; end_W(34, 115) <= 1; end_W(34, 116) <= 1; end_W(34, 117) <= 1; end_W(34, 118) <= 1; end_W(34, 119) <= 1; 
end_W(34, 120) <= 0; end_W(34, 121) <= 0; end_W(34, 122) <= 0; end_W(34, 123) <= 0; end_W(34, 124) <= 0; end_W(34, 125) <= 0; end_W(34, 126) <= 0; end_W(34, 127) <= 0; 
end_W(34, 128) <= 1; end_W(34, 129) <= 1; end_W(34, 130) <= 1; end_W(34, 131) <= 1; end_W(34, 132) <= 1; end_W(34, 133) <= 1; end_W(34, 134) <= 1; end_W(34, 135) <= 1; 
end_W(34, 136) <= 0; end_W(34, 137) <= 0; end_W(34, 138) <= 0; end_W(34, 139) <= 0; end_W(34, 140) <= 0; end_W(34, 141) <= 0; end_W(34, 142) <= 0; end_W(34, 143) <= 0; 
end_W(34, 144) <= 0; end_W(34, 145) <= 0; end_W(34, 146) <= 0; end_W(34, 147) <= 0; end_W(34, 148) <= 0; end_W(34, 149) <= 0; end_W(34, 150) <= 0; end_W(34, 151) <= 0; 
end_W(34, 152) <= 0; end_W(34, 153) <= 0; end_W(34, 154) <= 0; end_W(34, 155) <= 0; end_W(34, 156) <= 0; end_W(34, 157) <= 0; end_W(34, 158) <= 0; end_W(34, 159) <= 0; 
end_W(34, 160) <= 0; end_W(34, 161) <= 0; end_W(34, 162) <= 0; end_W(34, 163) <= 0; end_W(34, 164) <= 0; end_W(34, 165) <= 0; end_W(34, 166) <= 0; end_W(34, 167) <= 0; 
end_W(34, 168) <= 0; end_W(34, 169) <= 0; end_W(34, 170) <= 0; end_W(34, 171) <= 0; end_W(34, 172) <= 0; end_W(34, 173) <= 0; end_W(34, 174) <= 0; end_W(34, 175) <= 0; 
end_W(34, 176) <= 0; end_W(34, 177) <= 0; end_W(34, 178) <= 0; end_W(34, 179) <= 0; end_W(34, 180) <= 1; end_W(34, 181) <= 1; end_W(34, 182) <= 1; end_W(34, 183) <= 1; 
end_W(34, 184) <= 1; end_W(34, 185) <= 1; end_W(34, 186) <= 1; end_W(34, 187) <= 1; end_W(34, 188) <= 0; end_W(34, 189) <= 0; end_W(34, 190) <= 0; end_W(34, 191) <= 0; 
end_W(34, 192) <= 0; end_W(34, 193) <= 0; end_W(34, 194) <= 0; end_W(34, 195) <= 0; end_W(34, 196) <= 0; end_W(34, 197) <= 0; end_W(34, 198) <= 0; end_W(34, 199) <= 0; 
end_W(34, 200) <= 1; end_W(34, 201) <= 1; end_W(34, 202) <= 1; end_W(34, 203) <= 1; end_W(34, 204) <= 1; end_W(34, 205) <= 1; end_W(34, 206) <= 1; end_W(34, 207) <= 1; 
end_W(34, 208) <= 0; end_W(34, 209) <= 0; end_W(34, 210) <= 0; end_W(34, 211) <= 0; end_W(34, 212) <= 0; end_W(34, 213) <= 0; end_W(34, 214) <= 0; end_W(34, 215) <= 0; 
end_W(34, 216) <= 0; end_W(34, 217) <= 0; end_W(34, 218) <= 0; end_W(34, 219) <= 0; end_W(34, 220) <= 0; end_W(34, 221) <= 0; end_W(34, 222) <= 0; end_W(34, 223) <= 0; 
end_W(34, 224) <= 1; end_W(34, 225) <= 1; end_W(34, 226) <= 1; end_W(34, 227) <= 1; end_W(34, 228) <= 1; end_W(34, 229) <= 1; end_W(34, 230) <= 1; end_W(34, 231) <= 1; 
end_W(34, 232) <= 1; end_W(34, 233) <= 1; end_W(34, 234) <= 1; end_W(34, 235) <= 1; end_W(34, 236) <= 1; end_W(34, 237) <= 1; end_W(34, 238) <= 1; end_W(34, 239) <= 1; 
end_W(34, 240) <= 0; end_W(34, 241) <= 0; end_W(34, 242) <= 0; end_W(34, 243) <= 0; end_W(34, 244) <= 0; end_W(34, 245) <= 0; end_W(34, 246) <= 0; end_W(34, 247) <= 0; 
end_W(34, 248) <= 0; end_W(34, 249) <= 0; end_W(34, 250) <= 0; end_W(34, 251) <= 0; end_W(34, 252) <= 0; end_W(34, 253) <= 0; end_W(34, 254) <= 0; end_W(34, 255) <= 0; 
end_W(34, 256) <= 1; end_W(34, 257) <= 1; end_W(34, 258) <= 1; end_W(34, 259) <= 1; end_W(34, 260) <= 1; end_W(34, 261) <= 1; end_W(34, 262) <= 1; end_W(34, 263) <= 1; 
end_W(34, 264) <= 0; end_W(34, 265) <= 0; end_W(34, 266) <= 0; end_W(34, 267) <= 0; end_W(34, 268) <= 0; end_W(34, 269) <= 0; end_W(34, 270) <= 0; end_W(34, 271) <= 0; 
end_W(34, 272) <= 1; end_W(34, 273) <= 1; end_W(34, 274) <= 1; end_W(34, 275) <= 1; end_W(34, 276) <= 1; end_W(34, 277) <= 1; end_W(34, 278) <= 1; end_W(34, 279) <= 1; 
end_W(34, 280) <= 0; end_W(34, 281) <= 0; end_W(34, 282) <= 0; end_W(34, 283) <= 0; end_W(34, 284) <= 0; end_W(34, 285) <= 0; end_W(34, 286) <= 0; end_W(34, 287) <= 0; 
end_W(34, 288) <= 0; end_W(34, 289) <= 0; end_W(34, 290) <= 0; end_W(34, 291) <= 0; end_W(34, 292) <= 1; end_W(34, 293) <= 1; end_W(34, 294) <= 1; end_W(34, 295) <= 1; 
end_W(34, 296) <= 1; end_W(34, 297) <= 1; end_W(34, 298) <= 1; end_W(34, 299) <= 1; end_W(34, 300) <= 0; end_W(34, 301) <= 0; end_W(34, 302) <= 0; end_W(34, 303) <= 0; 
end_W(34, 304) <= 0; end_W(34, 305) <= 0; end_W(34, 306) <= 0; end_W(34, 307) <= 0; end_W(34, 308) <= 1; end_W(34, 309) <= 1; end_W(34, 310) <= 1; end_W(34, 311) <= 1; 
end_W(34, 312) <= 1; end_W(34, 313) <= 1; end_W(34, 314) <= 1; end_W(34, 315) <= 1; end_W(34, 316) <= 0; end_W(34, 317) <= 0; end_W(34, 318) <= 0; end_W(34, 319) <= 0; 
end_W(34, 320) <= 0; end_W(34, 321) <= 0; end_W(34, 322) <= 0; end_W(34, 323) <= 0; end_W(35, 0) <= 0; end_W(35, 1) <= 0; end_W(35, 2) <= 0; end_W(35, 3) <= 0; end_W(35, 4) <= 1; end_W(35, 5) <= 1; end_W(35, 6) <= 1; end_W(35, 7) <= 1; 
end_W(35, 8) <= 1; end_W(35, 9) <= 1; end_W(35, 10) <= 1; end_W(35, 11) <= 1; end_W(35, 12) <= 0; end_W(35, 13) <= 0; end_W(35, 14) <= 0; end_W(35, 15) <= 0; 
end_W(35, 16) <= 0; end_W(35, 17) <= 0; end_W(35, 18) <= 0; end_W(35, 19) <= 0; end_W(35, 20) <= 1; end_W(35, 21) <= 1; end_W(35, 22) <= 1; end_W(35, 23) <= 1; 
end_W(35, 24) <= 1; end_W(35, 25) <= 1; end_W(35, 26) <= 1; end_W(35, 27) <= 1; end_W(35, 28) <= 0; end_W(35, 29) <= 0; end_W(35, 30) <= 0; end_W(35, 31) <= 0; 
end_W(35, 32) <= 0; end_W(35, 33) <= 0; end_W(35, 34) <= 0; end_W(35, 35) <= 0; end_W(35, 36) <= 1; end_W(35, 37) <= 1; end_W(35, 38) <= 1; end_W(35, 39) <= 1; 
end_W(35, 40) <= 1; end_W(35, 41) <= 1; end_W(35, 42) <= 1; end_W(35, 43) <= 1; end_W(35, 44) <= 0; end_W(35, 45) <= 0; end_W(35, 46) <= 0; end_W(35, 47) <= 0; 
end_W(35, 48) <= 0; end_W(35, 49) <= 0; end_W(35, 50) <= 0; end_W(35, 51) <= 0; end_W(35, 52) <= 0; end_W(35, 53) <= 0; end_W(35, 54) <= 0; end_W(35, 55) <= 0; 
end_W(35, 56) <= 1; end_W(35, 57) <= 1; end_W(35, 58) <= 1; end_W(35, 59) <= 1; end_W(35, 60) <= 1; end_W(35, 61) <= 1; end_W(35, 62) <= 1; end_W(35, 63) <= 1; 
end_W(35, 64) <= 0; end_W(35, 65) <= 0; end_W(35, 66) <= 0; end_W(35, 67) <= 0; end_W(35, 68) <= 0; end_W(35, 69) <= 0; end_W(35, 70) <= 0; end_W(35, 71) <= 0; 
end_W(35, 72) <= 1; end_W(35, 73) <= 1; end_W(35, 74) <= 1; end_W(35, 75) <= 1; end_W(35, 76) <= 1; end_W(35, 77) <= 1; end_W(35, 78) <= 1; end_W(35, 79) <= 1; 
end_W(35, 80) <= 0; end_W(35, 81) <= 0; end_W(35, 82) <= 0; end_W(35, 83) <= 0; end_W(35, 84) <= 0; end_W(35, 85) <= 0; end_W(35, 86) <= 0; end_W(35, 87) <= 0; 
end_W(35, 88) <= 0; end_W(35, 89) <= 0; end_W(35, 90) <= 0; end_W(35, 91) <= 0; end_W(35, 92) <= 0; end_W(35, 93) <= 0; end_W(35, 94) <= 0; end_W(35, 95) <= 0; 
end_W(35, 96) <= 1; end_W(35, 97) <= 1; end_W(35, 98) <= 1; end_W(35, 99) <= 1; end_W(35, 100) <= 1; end_W(35, 101) <= 1; end_W(35, 102) <= 1; end_W(35, 103) <= 1; 
end_W(35, 104) <= 0; end_W(35, 105) <= 0; end_W(35, 106) <= 0; end_W(35, 107) <= 0; end_W(35, 108) <= 0; end_W(35, 109) <= 0; end_W(35, 110) <= 0; end_W(35, 111) <= 0; 
end_W(35, 112) <= 1; end_W(35, 113) <= 1; end_W(35, 114) <= 1; end_W(35, 115) <= 1; end_W(35, 116) <= 1; end_W(35, 117) <= 1; end_W(35, 118) <= 1; end_W(35, 119) <= 1; 
end_W(35, 120) <= 0; end_W(35, 121) <= 0; end_W(35, 122) <= 0; end_W(35, 123) <= 0; end_W(35, 124) <= 0; end_W(35, 125) <= 0; end_W(35, 126) <= 0; end_W(35, 127) <= 0; 
end_W(35, 128) <= 1; end_W(35, 129) <= 1; end_W(35, 130) <= 1; end_W(35, 131) <= 1; end_W(35, 132) <= 1; end_W(35, 133) <= 1; end_W(35, 134) <= 1; end_W(35, 135) <= 1; 
end_W(35, 136) <= 0; end_W(35, 137) <= 0; end_W(35, 138) <= 0; end_W(35, 139) <= 0; end_W(35, 140) <= 0; end_W(35, 141) <= 0; end_W(35, 142) <= 0; end_W(35, 143) <= 0; 
end_W(35, 144) <= 0; end_W(35, 145) <= 0; end_W(35, 146) <= 0; end_W(35, 147) <= 0; end_W(35, 148) <= 0; end_W(35, 149) <= 0; end_W(35, 150) <= 0; end_W(35, 151) <= 0; 
end_W(35, 152) <= 0; end_W(35, 153) <= 0; end_W(35, 154) <= 0; end_W(35, 155) <= 0; end_W(35, 156) <= 0; end_W(35, 157) <= 0; end_W(35, 158) <= 0; end_W(35, 159) <= 0; 
end_W(35, 160) <= 0; end_W(35, 161) <= 0; end_W(35, 162) <= 0; end_W(35, 163) <= 0; end_W(35, 164) <= 0; end_W(35, 165) <= 0; end_W(35, 166) <= 0; end_W(35, 167) <= 0; 
end_W(35, 168) <= 0; end_W(35, 169) <= 0; end_W(35, 170) <= 0; end_W(35, 171) <= 0; end_W(35, 172) <= 0; end_W(35, 173) <= 0; end_W(35, 174) <= 0; end_W(35, 175) <= 0; 
end_W(35, 176) <= 0; end_W(35, 177) <= 0; end_W(35, 178) <= 0; end_W(35, 179) <= 0; end_W(35, 180) <= 1; end_W(35, 181) <= 1; end_W(35, 182) <= 1; end_W(35, 183) <= 1; 
end_W(35, 184) <= 1; end_W(35, 185) <= 1; end_W(35, 186) <= 1; end_W(35, 187) <= 1; end_W(35, 188) <= 0; end_W(35, 189) <= 0; end_W(35, 190) <= 0; end_W(35, 191) <= 0; 
end_W(35, 192) <= 0; end_W(35, 193) <= 0; end_W(35, 194) <= 0; end_W(35, 195) <= 0; end_W(35, 196) <= 0; end_W(35, 197) <= 0; end_W(35, 198) <= 0; end_W(35, 199) <= 0; 
end_W(35, 200) <= 1; end_W(35, 201) <= 1; end_W(35, 202) <= 1; end_W(35, 203) <= 1; end_W(35, 204) <= 1; end_W(35, 205) <= 1; end_W(35, 206) <= 1; end_W(35, 207) <= 1; 
end_W(35, 208) <= 0; end_W(35, 209) <= 0; end_W(35, 210) <= 0; end_W(35, 211) <= 0; end_W(35, 212) <= 0; end_W(35, 213) <= 0; end_W(35, 214) <= 0; end_W(35, 215) <= 0; 
end_W(35, 216) <= 0; end_W(35, 217) <= 0; end_W(35, 218) <= 0; end_W(35, 219) <= 0; end_W(35, 220) <= 0; end_W(35, 221) <= 0; end_W(35, 222) <= 0; end_W(35, 223) <= 0; 
end_W(35, 224) <= 1; end_W(35, 225) <= 1; end_W(35, 226) <= 1; end_W(35, 227) <= 1; end_W(35, 228) <= 1; end_W(35, 229) <= 1; end_W(35, 230) <= 1; end_W(35, 231) <= 1; 
end_W(35, 232) <= 1; end_W(35, 233) <= 1; end_W(35, 234) <= 1; end_W(35, 235) <= 1; end_W(35, 236) <= 1; end_W(35, 237) <= 1; end_W(35, 238) <= 1; end_W(35, 239) <= 1; 
end_W(35, 240) <= 0; end_W(35, 241) <= 0; end_W(35, 242) <= 0; end_W(35, 243) <= 0; end_W(35, 244) <= 0; end_W(35, 245) <= 0; end_W(35, 246) <= 0; end_W(35, 247) <= 0; 
end_W(35, 248) <= 0; end_W(35, 249) <= 0; end_W(35, 250) <= 0; end_W(35, 251) <= 0; end_W(35, 252) <= 0; end_W(35, 253) <= 0; end_W(35, 254) <= 0; end_W(35, 255) <= 0; 
end_W(35, 256) <= 1; end_W(35, 257) <= 1; end_W(35, 258) <= 1; end_W(35, 259) <= 1; end_W(35, 260) <= 1; end_W(35, 261) <= 1; end_W(35, 262) <= 1; end_W(35, 263) <= 1; 
end_W(35, 264) <= 0; end_W(35, 265) <= 0; end_W(35, 266) <= 0; end_W(35, 267) <= 0; end_W(35, 268) <= 0; end_W(35, 269) <= 0; end_W(35, 270) <= 0; end_W(35, 271) <= 0; 
end_W(35, 272) <= 1; end_W(35, 273) <= 1; end_W(35, 274) <= 1; end_W(35, 275) <= 1; end_W(35, 276) <= 1; end_W(35, 277) <= 1; end_W(35, 278) <= 1; end_W(35, 279) <= 1; 
end_W(35, 280) <= 0; end_W(35, 281) <= 0; end_W(35, 282) <= 0; end_W(35, 283) <= 0; end_W(35, 284) <= 0; end_W(35, 285) <= 0; end_W(35, 286) <= 0; end_W(35, 287) <= 0; 
end_W(35, 288) <= 0; end_W(35, 289) <= 0; end_W(35, 290) <= 0; end_W(35, 291) <= 0; end_W(35, 292) <= 1; end_W(35, 293) <= 1; end_W(35, 294) <= 1; end_W(35, 295) <= 1; 
end_W(35, 296) <= 1; end_W(35, 297) <= 1; end_W(35, 298) <= 1; end_W(35, 299) <= 1; end_W(35, 300) <= 0; end_W(35, 301) <= 0; end_W(35, 302) <= 0; end_W(35, 303) <= 0; 
end_W(35, 304) <= 0; end_W(35, 305) <= 0; end_W(35, 306) <= 0; end_W(35, 307) <= 0; end_W(35, 308) <= 1; end_W(35, 309) <= 1; end_W(35, 310) <= 1; end_W(35, 311) <= 1; 
end_W(35, 312) <= 1; end_W(35, 313) <= 1; end_W(35, 314) <= 1; end_W(35, 315) <= 1; end_W(35, 316) <= 0; end_W(35, 317) <= 0; end_W(35, 318) <= 0; end_W(35, 319) <= 0; 
end_W(35, 320) <= 0; end_W(35, 321) <= 0; end_W(35, 322) <= 0; end_W(35, 323) <= 0; end_W(36, 0) <= 0; end_W(36, 1) <= 0; end_W(36, 2) <= 0; end_W(36, 3) <= 0; end_W(36, 4) <= 0; end_W(36, 5) <= 0; end_W(36, 6) <= 0; end_W(36, 7) <= 0; 
end_W(36, 8) <= 1; end_W(36, 9) <= 1; end_W(36, 10) <= 1; end_W(36, 11) <= 1; end_W(36, 12) <= 1; end_W(36, 13) <= 1; end_W(36, 14) <= 1; end_W(36, 15) <= 1; 
end_W(36, 16) <= 1; end_W(36, 17) <= 1; end_W(36, 18) <= 1; end_W(36, 19) <= 1; end_W(36, 20) <= 0; end_W(36, 21) <= 0; end_W(36, 22) <= 0; end_W(36, 23) <= 0; 
end_W(36, 24) <= 1; end_W(36, 25) <= 1; end_W(36, 26) <= 1; end_W(36, 27) <= 1; end_W(36, 28) <= 0; end_W(36, 29) <= 0; end_W(36, 30) <= 0; end_W(36, 31) <= 0; 
end_W(36, 32) <= 0; end_W(36, 33) <= 0; end_W(36, 34) <= 0; end_W(36, 35) <= 0; end_W(36, 36) <= 1; end_W(36, 37) <= 1; end_W(36, 38) <= 1; end_W(36, 39) <= 1; 
end_W(36, 40) <= 1; end_W(36, 41) <= 1; end_W(36, 42) <= 1; end_W(36, 43) <= 1; end_W(36, 44) <= 0; end_W(36, 45) <= 0; end_W(36, 46) <= 0; end_W(36, 47) <= 0; 
end_W(36, 48) <= 0; end_W(36, 49) <= 0; end_W(36, 50) <= 0; end_W(36, 51) <= 0; end_W(36, 52) <= 0; end_W(36, 53) <= 0; end_W(36, 54) <= 0; end_W(36, 55) <= 0; 
end_W(36, 56) <= 1; end_W(36, 57) <= 1; end_W(36, 58) <= 1; end_W(36, 59) <= 1; end_W(36, 60) <= 1; end_W(36, 61) <= 1; end_W(36, 62) <= 1; end_W(36, 63) <= 1; 
end_W(36, 64) <= 0; end_W(36, 65) <= 0; end_W(36, 66) <= 0; end_W(36, 67) <= 0; end_W(36, 68) <= 0; end_W(36, 69) <= 0; end_W(36, 70) <= 0; end_W(36, 71) <= 0; 
end_W(36, 72) <= 1; end_W(36, 73) <= 1; end_W(36, 74) <= 1; end_W(36, 75) <= 1; end_W(36, 76) <= 1; end_W(36, 77) <= 1; end_W(36, 78) <= 1; end_W(36, 79) <= 1; 
end_W(36, 80) <= 0; end_W(36, 81) <= 0; end_W(36, 82) <= 0; end_W(36, 83) <= 0; end_W(36, 84) <= 0; end_W(36, 85) <= 0; end_W(36, 86) <= 0; end_W(36, 87) <= 0; 
end_W(36, 88) <= 0; end_W(36, 89) <= 0; end_W(36, 90) <= 0; end_W(36, 91) <= 0; end_W(36, 92) <= 0; end_W(36, 93) <= 0; end_W(36, 94) <= 0; end_W(36, 95) <= 0; 
end_W(36, 96) <= 1; end_W(36, 97) <= 1; end_W(36, 98) <= 1; end_W(36, 99) <= 1; end_W(36, 100) <= 1; end_W(36, 101) <= 1; end_W(36, 102) <= 1; end_W(36, 103) <= 1; 
end_W(36, 104) <= 0; end_W(36, 105) <= 0; end_W(36, 106) <= 0; end_W(36, 107) <= 0; end_W(36, 108) <= 1; end_W(36, 109) <= 1; end_W(36, 110) <= 1; end_W(36, 111) <= 1; 
end_W(36, 112) <= 1; end_W(36, 113) <= 1; end_W(36, 114) <= 1; end_W(36, 115) <= 1; end_W(36, 116) <= 1; end_W(36, 117) <= 1; end_W(36, 118) <= 1; end_W(36, 119) <= 1; 
end_W(36, 120) <= 1; end_W(36, 121) <= 1; end_W(36, 122) <= 1; end_W(36, 123) <= 1; end_W(36, 124) <= 1; end_W(36, 125) <= 1; end_W(36, 126) <= 1; end_W(36, 127) <= 1; 
end_W(36, 128) <= 1; end_W(36, 129) <= 1; end_W(36, 130) <= 1; end_W(36, 131) <= 1; end_W(36, 132) <= 1; end_W(36, 133) <= 1; end_W(36, 134) <= 1; end_W(36, 135) <= 1; 
end_W(36, 136) <= 0; end_W(36, 137) <= 0; end_W(36, 138) <= 0; end_W(36, 139) <= 0; end_W(36, 140) <= 0; end_W(36, 141) <= 0; end_W(36, 142) <= 0; end_W(36, 143) <= 0; 
end_W(36, 144) <= 0; end_W(36, 145) <= 0; end_W(36, 146) <= 0; end_W(36, 147) <= 0; end_W(36, 148) <= 0; end_W(36, 149) <= 0; end_W(36, 150) <= 0; end_W(36, 151) <= 0; 
end_W(36, 152) <= 0; end_W(36, 153) <= 0; end_W(36, 154) <= 0; end_W(36, 155) <= 0; end_W(36, 156) <= 0; end_W(36, 157) <= 0; end_W(36, 158) <= 0; end_W(36, 159) <= 0; 
end_W(36, 160) <= 0; end_W(36, 161) <= 0; end_W(36, 162) <= 0; end_W(36, 163) <= 0; end_W(36, 164) <= 0; end_W(36, 165) <= 0; end_W(36, 166) <= 0; end_W(36, 167) <= 0; 
end_W(36, 168) <= 0; end_W(36, 169) <= 0; end_W(36, 170) <= 0; end_W(36, 171) <= 0; end_W(36, 172) <= 0; end_W(36, 173) <= 0; end_W(36, 174) <= 0; end_W(36, 175) <= 0; 
end_W(36, 176) <= 0; end_W(36, 177) <= 0; end_W(36, 178) <= 0; end_W(36, 179) <= 0; end_W(36, 180) <= 0; end_W(36, 181) <= 0; end_W(36, 182) <= 0; end_W(36, 183) <= 0; 
end_W(36, 184) <= 1; end_W(36, 185) <= 1; end_W(36, 186) <= 1; end_W(36, 187) <= 1; end_W(36, 188) <= 1; end_W(36, 189) <= 1; end_W(36, 190) <= 1; end_W(36, 191) <= 1; 
end_W(36, 192) <= 1; end_W(36, 193) <= 1; end_W(36, 194) <= 1; end_W(36, 195) <= 1; end_W(36, 196) <= 1; end_W(36, 197) <= 1; end_W(36, 198) <= 1; end_W(36, 199) <= 1; 
end_W(36, 200) <= 1; end_W(36, 201) <= 1; end_W(36, 202) <= 1; end_W(36, 203) <= 1; end_W(36, 204) <= 0; end_W(36, 205) <= 0; end_W(36, 206) <= 0; end_W(36, 207) <= 0; 
end_W(36, 208) <= 0; end_W(36, 209) <= 0; end_W(36, 210) <= 0; end_W(36, 211) <= 0; end_W(36, 212) <= 0; end_W(36, 213) <= 0; end_W(36, 214) <= 0; end_W(36, 215) <= 0; 
end_W(36, 216) <= 0; end_W(36, 217) <= 0; end_W(36, 218) <= 0; end_W(36, 219) <= 0; end_W(36, 220) <= 0; end_W(36, 221) <= 0; end_W(36, 222) <= 0; end_W(36, 223) <= 0; 
end_W(36, 224) <= 0; end_W(36, 225) <= 0; end_W(36, 226) <= 0; end_W(36, 227) <= 0; end_W(36, 228) <= 1; end_W(36, 229) <= 1; end_W(36, 230) <= 1; end_W(36, 231) <= 1; 
end_W(36, 232) <= 1; end_W(36, 233) <= 1; end_W(36, 234) <= 1; end_W(36, 235) <= 1; end_W(36, 236) <= 0; end_W(36, 237) <= 0; end_W(36, 238) <= 0; end_W(36, 239) <= 0; 
end_W(36, 240) <= 0; end_W(36, 241) <= 0; end_W(36, 242) <= 0; end_W(36, 243) <= 0; end_W(36, 244) <= 0; end_W(36, 245) <= 0; end_W(36, 246) <= 0; end_W(36, 247) <= 0; 
end_W(36, 248) <= 0; end_W(36, 249) <= 0; end_W(36, 250) <= 0; end_W(36, 251) <= 0; end_W(36, 252) <= 1; end_W(36, 253) <= 1; end_W(36, 254) <= 1; end_W(36, 255) <= 1; 
end_W(36, 256) <= 1; end_W(36, 257) <= 1; end_W(36, 258) <= 1; end_W(36, 259) <= 1; end_W(36, 260) <= 1; end_W(36, 261) <= 1; end_W(36, 262) <= 1; end_W(36, 263) <= 1; 
end_W(36, 264) <= 1; end_W(36, 265) <= 1; end_W(36, 266) <= 1; end_W(36, 267) <= 1; end_W(36, 268) <= 1; end_W(36, 269) <= 1; end_W(36, 270) <= 1; end_W(36, 271) <= 1; 
end_W(36, 272) <= 1; end_W(36, 273) <= 1; end_W(36, 274) <= 1; end_W(36, 275) <= 1; end_W(36, 276) <= 1; end_W(36, 277) <= 1; end_W(36, 278) <= 1; end_W(36, 279) <= 1; 
end_W(36, 280) <= 0; end_W(36, 281) <= 0; end_W(36, 282) <= 0; end_W(36, 283) <= 0; end_W(36, 284) <= 0; end_W(36, 285) <= 0; end_W(36, 286) <= 0; end_W(36, 287) <= 0; 
end_W(36, 288) <= 1; end_W(36, 289) <= 1; end_W(36, 290) <= 1; end_W(36, 291) <= 1; end_W(36, 292) <= 1; end_W(36, 293) <= 1; end_W(36, 294) <= 1; end_W(36, 295) <= 1; 
end_W(36, 296) <= 1; end_W(36, 297) <= 1; end_W(36, 298) <= 1; end_W(36, 299) <= 1; end_W(36, 300) <= 0; end_W(36, 301) <= 0; end_W(36, 302) <= 0; end_W(36, 303) <= 0; 
end_W(36, 304) <= 0; end_W(36, 305) <= 0; end_W(36, 306) <= 0; end_W(36, 307) <= 0; end_W(36, 308) <= 1; end_W(36, 309) <= 1; end_W(36, 310) <= 1; end_W(36, 311) <= 1; 
end_W(36, 312) <= 1; end_W(36, 313) <= 1; end_W(36, 314) <= 1; end_W(36, 315) <= 1; end_W(36, 316) <= 0; end_W(36, 317) <= 0; end_W(36, 318) <= 0; end_W(36, 319) <= 0; 
end_W(36, 320) <= 0; end_W(36, 321) <= 0; end_W(36, 322) <= 0; end_W(36, 323) <= 0; end_W(37, 0) <= 0; end_W(37, 1) <= 0; end_W(37, 2) <= 0; end_W(37, 3) <= 0; end_W(37, 4) <= 0; end_W(37, 5) <= 0; end_W(37, 6) <= 0; end_W(37, 7) <= 0; 
end_W(37, 8) <= 1; end_W(37, 9) <= 1; end_W(37, 10) <= 1; end_W(37, 11) <= 1; end_W(37, 12) <= 1; end_W(37, 13) <= 1; end_W(37, 14) <= 1; end_W(37, 15) <= 1; 
end_W(37, 16) <= 1; end_W(37, 17) <= 1; end_W(37, 18) <= 1; end_W(37, 19) <= 1; end_W(37, 20) <= 0; end_W(37, 21) <= 0; end_W(37, 22) <= 0; end_W(37, 23) <= 0; 
end_W(37, 24) <= 1; end_W(37, 25) <= 1; end_W(37, 26) <= 1; end_W(37, 27) <= 1; end_W(37, 28) <= 0; end_W(37, 29) <= 0; end_W(37, 30) <= 0; end_W(37, 31) <= 0; 
end_W(37, 32) <= 0; end_W(37, 33) <= 0; end_W(37, 34) <= 0; end_W(37, 35) <= 0; end_W(37, 36) <= 1; end_W(37, 37) <= 1; end_W(37, 38) <= 1; end_W(37, 39) <= 1; 
end_W(37, 40) <= 1; end_W(37, 41) <= 1; end_W(37, 42) <= 1; end_W(37, 43) <= 1; end_W(37, 44) <= 0; end_W(37, 45) <= 0; end_W(37, 46) <= 0; end_W(37, 47) <= 0; 
end_W(37, 48) <= 0; end_W(37, 49) <= 0; end_W(37, 50) <= 0; end_W(37, 51) <= 0; end_W(37, 52) <= 0; end_W(37, 53) <= 0; end_W(37, 54) <= 0; end_W(37, 55) <= 0; 
end_W(37, 56) <= 1; end_W(37, 57) <= 1; end_W(37, 58) <= 1; end_W(37, 59) <= 1; end_W(37, 60) <= 1; end_W(37, 61) <= 1; end_W(37, 62) <= 1; end_W(37, 63) <= 1; 
end_W(37, 64) <= 0; end_W(37, 65) <= 0; end_W(37, 66) <= 0; end_W(37, 67) <= 0; end_W(37, 68) <= 0; end_W(37, 69) <= 0; end_W(37, 70) <= 0; end_W(37, 71) <= 0; 
end_W(37, 72) <= 1; end_W(37, 73) <= 1; end_W(37, 74) <= 1; end_W(37, 75) <= 1; end_W(37, 76) <= 1; end_W(37, 77) <= 1; end_W(37, 78) <= 1; end_W(37, 79) <= 1; 
end_W(37, 80) <= 0; end_W(37, 81) <= 0; end_W(37, 82) <= 0; end_W(37, 83) <= 0; end_W(37, 84) <= 0; end_W(37, 85) <= 0; end_W(37, 86) <= 0; end_W(37, 87) <= 0; 
end_W(37, 88) <= 0; end_W(37, 89) <= 0; end_W(37, 90) <= 0; end_W(37, 91) <= 0; end_W(37, 92) <= 0; end_W(37, 93) <= 0; end_W(37, 94) <= 0; end_W(37, 95) <= 0; 
end_W(37, 96) <= 1; end_W(37, 97) <= 1; end_W(37, 98) <= 1; end_W(37, 99) <= 1; end_W(37, 100) <= 1; end_W(37, 101) <= 1; end_W(37, 102) <= 1; end_W(37, 103) <= 1; 
end_W(37, 104) <= 0; end_W(37, 105) <= 0; end_W(37, 106) <= 0; end_W(37, 107) <= 0; end_W(37, 108) <= 1; end_W(37, 109) <= 1; end_W(37, 110) <= 1; end_W(37, 111) <= 1; 
end_W(37, 112) <= 1; end_W(37, 113) <= 1; end_W(37, 114) <= 1; end_W(37, 115) <= 1; end_W(37, 116) <= 1; end_W(37, 117) <= 1; end_W(37, 118) <= 1; end_W(37, 119) <= 1; 
end_W(37, 120) <= 1; end_W(37, 121) <= 1; end_W(37, 122) <= 1; end_W(37, 123) <= 1; end_W(37, 124) <= 1; end_W(37, 125) <= 1; end_W(37, 126) <= 1; end_W(37, 127) <= 1; 
end_W(37, 128) <= 1; end_W(37, 129) <= 1; end_W(37, 130) <= 1; end_W(37, 131) <= 1; end_W(37, 132) <= 1; end_W(37, 133) <= 1; end_W(37, 134) <= 1; end_W(37, 135) <= 1; 
end_W(37, 136) <= 0; end_W(37, 137) <= 0; end_W(37, 138) <= 0; end_W(37, 139) <= 0; end_W(37, 140) <= 0; end_W(37, 141) <= 0; end_W(37, 142) <= 0; end_W(37, 143) <= 0; 
end_W(37, 144) <= 0; end_W(37, 145) <= 0; end_W(37, 146) <= 0; end_W(37, 147) <= 0; end_W(37, 148) <= 0; end_W(37, 149) <= 0; end_W(37, 150) <= 0; end_W(37, 151) <= 0; 
end_W(37, 152) <= 0; end_W(37, 153) <= 0; end_W(37, 154) <= 0; end_W(37, 155) <= 0; end_W(37, 156) <= 0; end_W(37, 157) <= 0; end_W(37, 158) <= 0; end_W(37, 159) <= 0; 
end_W(37, 160) <= 0; end_W(37, 161) <= 0; end_W(37, 162) <= 0; end_W(37, 163) <= 0; end_W(37, 164) <= 0; end_W(37, 165) <= 0; end_W(37, 166) <= 0; end_W(37, 167) <= 0; 
end_W(37, 168) <= 0; end_W(37, 169) <= 0; end_W(37, 170) <= 0; end_W(37, 171) <= 0; end_W(37, 172) <= 0; end_W(37, 173) <= 0; end_W(37, 174) <= 0; end_W(37, 175) <= 0; 
end_W(37, 176) <= 0; end_W(37, 177) <= 0; end_W(37, 178) <= 0; end_W(37, 179) <= 0; end_W(37, 180) <= 0; end_W(37, 181) <= 0; end_W(37, 182) <= 0; end_W(37, 183) <= 0; 
end_W(37, 184) <= 1; end_W(37, 185) <= 1; end_W(37, 186) <= 1; end_W(37, 187) <= 1; end_W(37, 188) <= 1; end_W(37, 189) <= 1; end_W(37, 190) <= 1; end_W(37, 191) <= 1; 
end_W(37, 192) <= 1; end_W(37, 193) <= 1; end_W(37, 194) <= 1; end_W(37, 195) <= 1; end_W(37, 196) <= 1; end_W(37, 197) <= 1; end_W(37, 198) <= 1; end_W(37, 199) <= 1; 
end_W(37, 200) <= 1; end_W(37, 201) <= 1; end_W(37, 202) <= 1; end_W(37, 203) <= 1; end_W(37, 204) <= 0; end_W(37, 205) <= 0; end_W(37, 206) <= 0; end_W(37, 207) <= 0; 
end_W(37, 208) <= 0; end_W(37, 209) <= 0; end_W(37, 210) <= 0; end_W(37, 211) <= 0; end_W(37, 212) <= 0; end_W(37, 213) <= 0; end_W(37, 214) <= 0; end_W(37, 215) <= 0; 
end_W(37, 216) <= 0; end_W(37, 217) <= 0; end_W(37, 218) <= 0; end_W(37, 219) <= 0; end_W(37, 220) <= 0; end_W(37, 221) <= 0; end_W(37, 222) <= 0; end_W(37, 223) <= 0; 
end_W(37, 224) <= 0; end_W(37, 225) <= 0; end_W(37, 226) <= 0; end_W(37, 227) <= 0; end_W(37, 228) <= 1; end_W(37, 229) <= 1; end_W(37, 230) <= 1; end_W(37, 231) <= 1; 
end_W(37, 232) <= 1; end_W(37, 233) <= 1; end_W(37, 234) <= 1; end_W(37, 235) <= 1; end_W(37, 236) <= 0; end_W(37, 237) <= 0; end_W(37, 238) <= 0; end_W(37, 239) <= 0; 
end_W(37, 240) <= 0; end_W(37, 241) <= 0; end_W(37, 242) <= 0; end_W(37, 243) <= 0; end_W(37, 244) <= 0; end_W(37, 245) <= 0; end_W(37, 246) <= 0; end_W(37, 247) <= 0; 
end_W(37, 248) <= 0; end_W(37, 249) <= 0; end_W(37, 250) <= 0; end_W(37, 251) <= 0; end_W(37, 252) <= 1; end_W(37, 253) <= 1; end_W(37, 254) <= 1; end_W(37, 255) <= 1; 
end_W(37, 256) <= 1; end_W(37, 257) <= 1; end_W(37, 258) <= 1; end_W(37, 259) <= 1; end_W(37, 260) <= 1; end_W(37, 261) <= 1; end_W(37, 262) <= 1; end_W(37, 263) <= 1; 
end_W(37, 264) <= 1; end_W(37, 265) <= 1; end_W(37, 266) <= 1; end_W(37, 267) <= 1; end_W(37, 268) <= 1; end_W(37, 269) <= 1; end_W(37, 270) <= 1; end_W(37, 271) <= 1; 
end_W(37, 272) <= 1; end_W(37, 273) <= 1; end_W(37, 274) <= 1; end_W(37, 275) <= 1; end_W(37, 276) <= 1; end_W(37, 277) <= 1; end_W(37, 278) <= 1; end_W(37, 279) <= 1; 
end_W(37, 280) <= 0; end_W(37, 281) <= 0; end_W(37, 282) <= 0; end_W(37, 283) <= 0; end_W(37, 284) <= 0; end_W(37, 285) <= 0; end_W(37, 286) <= 0; end_W(37, 287) <= 0; 
end_W(37, 288) <= 1; end_W(37, 289) <= 1; end_W(37, 290) <= 1; end_W(37, 291) <= 1; end_W(37, 292) <= 1; end_W(37, 293) <= 1; end_W(37, 294) <= 1; end_W(37, 295) <= 1; 
end_W(37, 296) <= 1; end_W(37, 297) <= 1; end_W(37, 298) <= 1; end_W(37, 299) <= 1; end_W(37, 300) <= 0; end_W(37, 301) <= 0; end_W(37, 302) <= 0; end_W(37, 303) <= 0; 
end_W(37, 304) <= 0; end_W(37, 305) <= 0; end_W(37, 306) <= 0; end_W(37, 307) <= 0; end_W(37, 308) <= 1; end_W(37, 309) <= 1; end_W(37, 310) <= 1; end_W(37, 311) <= 1; 
end_W(37, 312) <= 1; end_W(37, 313) <= 1; end_W(37, 314) <= 1; end_W(37, 315) <= 1; end_W(37, 316) <= 0; end_W(37, 317) <= 0; end_W(37, 318) <= 0; end_W(37, 319) <= 0; 
end_W(37, 320) <= 0; end_W(37, 321) <= 0; end_W(37, 322) <= 0; end_W(37, 323) <= 0; end_W(38, 0) <= 0; end_W(38, 1) <= 0; end_W(38, 2) <= 0; end_W(38, 3) <= 0; end_W(38, 4) <= 0; end_W(38, 5) <= 0; end_W(38, 6) <= 0; end_W(38, 7) <= 0; 
end_W(38, 8) <= 1; end_W(38, 9) <= 1; end_W(38, 10) <= 1; end_W(38, 11) <= 1; end_W(38, 12) <= 1; end_W(38, 13) <= 1; end_W(38, 14) <= 1; end_W(38, 15) <= 1; 
end_W(38, 16) <= 1; end_W(38, 17) <= 1; end_W(38, 18) <= 1; end_W(38, 19) <= 1; end_W(38, 20) <= 0; end_W(38, 21) <= 0; end_W(38, 22) <= 0; end_W(38, 23) <= 0; 
end_W(38, 24) <= 1; end_W(38, 25) <= 1; end_W(38, 26) <= 1; end_W(38, 27) <= 1; end_W(38, 28) <= 0; end_W(38, 29) <= 0; end_W(38, 30) <= 0; end_W(38, 31) <= 0; 
end_W(38, 32) <= 0; end_W(38, 33) <= 0; end_W(38, 34) <= 0; end_W(38, 35) <= 0; end_W(38, 36) <= 1; end_W(38, 37) <= 1; end_W(38, 38) <= 1; end_W(38, 39) <= 1; 
end_W(38, 40) <= 1; end_W(38, 41) <= 1; end_W(38, 42) <= 1; end_W(38, 43) <= 1; end_W(38, 44) <= 0; end_W(38, 45) <= 0; end_W(38, 46) <= 0; end_W(38, 47) <= 0; 
end_W(38, 48) <= 0; end_W(38, 49) <= 0; end_W(38, 50) <= 0; end_W(38, 51) <= 0; end_W(38, 52) <= 0; end_W(38, 53) <= 0; end_W(38, 54) <= 0; end_W(38, 55) <= 0; 
end_W(38, 56) <= 1; end_W(38, 57) <= 1; end_W(38, 58) <= 1; end_W(38, 59) <= 1; end_W(38, 60) <= 1; end_W(38, 61) <= 1; end_W(38, 62) <= 1; end_W(38, 63) <= 1; 
end_W(38, 64) <= 0; end_W(38, 65) <= 0; end_W(38, 66) <= 0; end_W(38, 67) <= 0; end_W(38, 68) <= 0; end_W(38, 69) <= 0; end_W(38, 70) <= 0; end_W(38, 71) <= 0; 
end_W(38, 72) <= 1; end_W(38, 73) <= 1; end_W(38, 74) <= 1; end_W(38, 75) <= 1; end_W(38, 76) <= 1; end_W(38, 77) <= 1; end_W(38, 78) <= 1; end_W(38, 79) <= 1; 
end_W(38, 80) <= 0; end_W(38, 81) <= 0; end_W(38, 82) <= 0; end_W(38, 83) <= 0; end_W(38, 84) <= 0; end_W(38, 85) <= 0; end_W(38, 86) <= 0; end_W(38, 87) <= 0; 
end_W(38, 88) <= 0; end_W(38, 89) <= 0; end_W(38, 90) <= 0; end_W(38, 91) <= 0; end_W(38, 92) <= 0; end_W(38, 93) <= 0; end_W(38, 94) <= 0; end_W(38, 95) <= 0; 
end_W(38, 96) <= 1; end_W(38, 97) <= 1; end_W(38, 98) <= 1; end_W(38, 99) <= 1; end_W(38, 100) <= 1; end_W(38, 101) <= 1; end_W(38, 102) <= 1; end_W(38, 103) <= 1; 
end_W(38, 104) <= 0; end_W(38, 105) <= 0; end_W(38, 106) <= 0; end_W(38, 107) <= 0; end_W(38, 108) <= 1; end_W(38, 109) <= 1; end_W(38, 110) <= 1; end_W(38, 111) <= 1; 
end_W(38, 112) <= 1; end_W(38, 113) <= 1; end_W(38, 114) <= 1; end_W(38, 115) <= 1; end_W(38, 116) <= 1; end_W(38, 117) <= 1; end_W(38, 118) <= 1; end_W(38, 119) <= 1; 
end_W(38, 120) <= 1; end_W(38, 121) <= 1; end_W(38, 122) <= 1; end_W(38, 123) <= 1; end_W(38, 124) <= 1; end_W(38, 125) <= 1; end_W(38, 126) <= 1; end_W(38, 127) <= 1; 
end_W(38, 128) <= 1; end_W(38, 129) <= 1; end_W(38, 130) <= 1; end_W(38, 131) <= 1; end_W(38, 132) <= 1; end_W(38, 133) <= 1; end_W(38, 134) <= 1; end_W(38, 135) <= 1; 
end_W(38, 136) <= 0; end_W(38, 137) <= 0; end_W(38, 138) <= 0; end_W(38, 139) <= 0; end_W(38, 140) <= 0; end_W(38, 141) <= 0; end_W(38, 142) <= 0; end_W(38, 143) <= 0; 
end_W(38, 144) <= 0; end_W(38, 145) <= 0; end_W(38, 146) <= 0; end_W(38, 147) <= 0; end_W(38, 148) <= 0; end_W(38, 149) <= 0; end_W(38, 150) <= 0; end_W(38, 151) <= 0; 
end_W(38, 152) <= 0; end_W(38, 153) <= 0; end_W(38, 154) <= 0; end_W(38, 155) <= 0; end_W(38, 156) <= 0; end_W(38, 157) <= 0; end_W(38, 158) <= 0; end_W(38, 159) <= 0; 
end_W(38, 160) <= 0; end_W(38, 161) <= 0; end_W(38, 162) <= 0; end_W(38, 163) <= 0; end_W(38, 164) <= 0; end_W(38, 165) <= 0; end_W(38, 166) <= 0; end_W(38, 167) <= 0; 
end_W(38, 168) <= 0; end_W(38, 169) <= 0; end_W(38, 170) <= 0; end_W(38, 171) <= 0; end_W(38, 172) <= 0; end_W(38, 173) <= 0; end_W(38, 174) <= 0; end_W(38, 175) <= 0; 
end_W(38, 176) <= 0; end_W(38, 177) <= 0; end_W(38, 178) <= 0; end_W(38, 179) <= 0; end_W(38, 180) <= 0; end_W(38, 181) <= 0; end_W(38, 182) <= 0; end_W(38, 183) <= 0; 
end_W(38, 184) <= 1; end_W(38, 185) <= 1; end_W(38, 186) <= 1; end_W(38, 187) <= 1; end_W(38, 188) <= 1; end_W(38, 189) <= 1; end_W(38, 190) <= 1; end_W(38, 191) <= 1; 
end_W(38, 192) <= 1; end_W(38, 193) <= 1; end_W(38, 194) <= 1; end_W(38, 195) <= 1; end_W(38, 196) <= 1; end_W(38, 197) <= 1; end_W(38, 198) <= 1; end_W(38, 199) <= 1; 
end_W(38, 200) <= 1; end_W(38, 201) <= 1; end_W(38, 202) <= 1; end_W(38, 203) <= 1; end_W(38, 204) <= 0; end_W(38, 205) <= 0; end_W(38, 206) <= 0; end_W(38, 207) <= 0; 
end_W(38, 208) <= 0; end_W(38, 209) <= 0; end_W(38, 210) <= 0; end_W(38, 211) <= 0; end_W(38, 212) <= 0; end_W(38, 213) <= 0; end_W(38, 214) <= 0; end_W(38, 215) <= 0; 
end_W(38, 216) <= 0; end_W(38, 217) <= 0; end_W(38, 218) <= 0; end_W(38, 219) <= 0; end_W(38, 220) <= 0; end_W(38, 221) <= 0; end_W(38, 222) <= 0; end_W(38, 223) <= 0; 
end_W(38, 224) <= 0; end_W(38, 225) <= 0; end_W(38, 226) <= 0; end_W(38, 227) <= 0; end_W(38, 228) <= 1; end_W(38, 229) <= 1; end_W(38, 230) <= 1; end_W(38, 231) <= 1; 
end_W(38, 232) <= 1; end_W(38, 233) <= 1; end_W(38, 234) <= 1; end_W(38, 235) <= 1; end_W(38, 236) <= 0; end_W(38, 237) <= 0; end_W(38, 238) <= 0; end_W(38, 239) <= 0; 
end_W(38, 240) <= 0; end_W(38, 241) <= 0; end_W(38, 242) <= 0; end_W(38, 243) <= 0; end_W(38, 244) <= 0; end_W(38, 245) <= 0; end_W(38, 246) <= 0; end_W(38, 247) <= 0; 
end_W(38, 248) <= 0; end_W(38, 249) <= 0; end_W(38, 250) <= 0; end_W(38, 251) <= 0; end_W(38, 252) <= 1; end_W(38, 253) <= 1; end_W(38, 254) <= 1; end_W(38, 255) <= 1; 
end_W(38, 256) <= 1; end_W(38, 257) <= 1; end_W(38, 258) <= 1; end_W(38, 259) <= 1; end_W(38, 260) <= 1; end_W(38, 261) <= 1; end_W(38, 262) <= 1; end_W(38, 263) <= 1; 
end_W(38, 264) <= 1; end_W(38, 265) <= 1; end_W(38, 266) <= 1; end_W(38, 267) <= 1; end_W(38, 268) <= 1; end_W(38, 269) <= 1; end_W(38, 270) <= 1; end_W(38, 271) <= 1; 
end_W(38, 272) <= 1; end_W(38, 273) <= 1; end_W(38, 274) <= 1; end_W(38, 275) <= 1; end_W(38, 276) <= 1; end_W(38, 277) <= 1; end_W(38, 278) <= 1; end_W(38, 279) <= 1; 
end_W(38, 280) <= 0; end_W(38, 281) <= 0; end_W(38, 282) <= 0; end_W(38, 283) <= 0; end_W(38, 284) <= 0; end_W(38, 285) <= 0; end_W(38, 286) <= 0; end_W(38, 287) <= 0; 
end_W(38, 288) <= 1; end_W(38, 289) <= 1; end_W(38, 290) <= 1; end_W(38, 291) <= 1; end_W(38, 292) <= 1; end_W(38, 293) <= 1; end_W(38, 294) <= 1; end_W(38, 295) <= 1; 
end_W(38, 296) <= 1; end_W(38, 297) <= 1; end_W(38, 298) <= 1; end_W(38, 299) <= 1; end_W(38, 300) <= 0; end_W(38, 301) <= 0; end_W(38, 302) <= 0; end_W(38, 303) <= 0; 
end_W(38, 304) <= 0; end_W(38, 305) <= 0; end_W(38, 306) <= 0; end_W(38, 307) <= 0; end_W(38, 308) <= 1; end_W(38, 309) <= 1; end_W(38, 310) <= 1; end_W(38, 311) <= 1; 
end_W(38, 312) <= 1; end_W(38, 313) <= 1; end_W(38, 314) <= 1; end_W(38, 315) <= 1; end_W(38, 316) <= 0; end_W(38, 317) <= 0; end_W(38, 318) <= 0; end_W(38, 319) <= 0; 
end_W(38, 320) <= 0; end_W(38, 321) <= 0; end_W(38, 322) <= 0; end_W(38, 323) <= 0; end_W(39, 0) <= 0; end_W(39, 1) <= 0; end_W(39, 2) <= 0; end_W(39, 3) <= 0; end_W(39, 4) <= 0; end_W(39, 5) <= 0; end_W(39, 6) <= 0; end_W(39, 7) <= 0; 
end_W(39, 8) <= 1; end_W(39, 9) <= 1; end_W(39, 10) <= 1; end_W(39, 11) <= 1; end_W(39, 12) <= 1; end_W(39, 13) <= 1; end_W(39, 14) <= 1; end_W(39, 15) <= 1; 
end_W(39, 16) <= 1; end_W(39, 17) <= 1; end_W(39, 18) <= 1; end_W(39, 19) <= 1; end_W(39, 20) <= 0; end_W(39, 21) <= 0; end_W(39, 22) <= 0; end_W(39, 23) <= 0; 
end_W(39, 24) <= 1; end_W(39, 25) <= 1; end_W(39, 26) <= 1; end_W(39, 27) <= 1; end_W(39, 28) <= 0; end_W(39, 29) <= 0; end_W(39, 30) <= 0; end_W(39, 31) <= 0; 
end_W(39, 32) <= 0; end_W(39, 33) <= 0; end_W(39, 34) <= 0; end_W(39, 35) <= 0; end_W(39, 36) <= 1; end_W(39, 37) <= 1; end_W(39, 38) <= 1; end_W(39, 39) <= 1; 
end_W(39, 40) <= 1; end_W(39, 41) <= 1; end_W(39, 42) <= 1; end_W(39, 43) <= 1; end_W(39, 44) <= 0; end_W(39, 45) <= 0; end_W(39, 46) <= 0; end_W(39, 47) <= 0; 
end_W(39, 48) <= 0; end_W(39, 49) <= 0; end_W(39, 50) <= 0; end_W(39, 51) <= 0; end_W(39, 52) <= 0; end_W(39, 53) <= 0; end_W(39, 54) <= 0; end_W(39, 55) <= 0; 
end_W(39, 56) <= 1; end_W(39, 57) <= 1; end_W(39, 58) <= 1; end_W(39, 59) <= 1; end_W(39, 60) <= 1; end_W(39, 61) <= 1; end_W(39, 62) <= 1; end_W(39, 63) <= 1; 
end_W(39, 64) <= 0; end_W(39, 65) <= 0; end_W(39, 66) <= 0; end_W(39, 67) <= 0; end_W(39, 68) <= 0; end_W(39, 69) <= 0; end_W(39, 70) <= 0; end_W(39, 71) <= 0; 
end_W(39, 72) <= 1; end_W(39, 73) <= 1; end_W(39, 74) <= 1; end_W(39, 75) <= 1; end_W(39, 76) <= 1; end_W(39, 77) <= 1; end_W(39, 78) <= 1; end_W(39, 79) <= 1; 
end_W(39, 80) <= 0; end_W(39, 81) <= 0; end_W(39, 82) <= 0; end_W(39, 83) <= 0; end_W(39, 84) <= 0; end_W(39, 85) <= 0; end_W(39, 86) <= 0; end_W(39, 87) <= 0; 
end_W(39, 88) <= 0; end_W(39, 89) <= 0; end_W(39, 90) <= 0; end_W(39, 91) <= 0; end_W(39, 92) <= 0; end_W(39, 93) <= 0; end_W(39, 94) <= 0; end_W(39, 95) <= 0; 
end_W(39, 96) <= 1; end_W(39, 97) <= 1; end_W(39, 98) <= 1; end_W(39, 99) <= 1; end_W(39, 100) <= 1; end_W(39, 101) <= 1; end_W(39, 102) <= 1; end_W(39, 103) <= 1; 
end_W(39, 104) <= 0; end_W(39, 105) <= 0; end_W(39, 106) <= 0; end_W(39, 107) <= 0; end_W(39, 108) <= 1; end_W(39, 109) <= 1; end_W(39, 110) <= 1; end_W(39, 111) <= 1; 
end_W(39, 112) <= 1; end_W(39, 113) <= 1; end_W(39, 114) <= 1; end_W(39, 115) <= 1; end_W(39, 116) <= 1; end_W(39, 117) <= 1; end_W(39, 118) <= 1; end_W(39, 119) <= 1; 
end_W(39, 120) <= 1; end_W(39, 121) <= 1; end_W(39, 122) <= 1; end_W(39, 123) <= 1; end_W(39, 124) <= 1; end_W(39, 125) <= 1; end_W(39, 126) <= 1; end_W(39, 127) <= 1; 
end_W(39, 128) <= 1; end_W(39, 129) <= 1; end_W(39, 130) <= 1; end_W(39, 131) <= 1; end_W(39, 132) <= 1; end_W(39, 133) <= 1; end_W(39, 134) <= 1; end_W(39, 135) <= 1; 
end_W(39, 136) <= 0; end_W(39, 137) <= 0; end_W(39, 138) <= 0; end_W(39, 139) <= 0; end_W(39, 140) <= 0; end_W(39, 141) <= 0; end_W(39, 142) <= 0; end_W(39, 143) <= 0; 
end_W(39, 144) <= 0; end_W(39, 145) <= 0; end_W(39, 146) <= 0; end_W(39, 147) <= 0; end_W(39, 148) <= 0; end_W(39, 149) <= 0; end_W(39, 150) <= 0; end_W(39, 151) <= 0; 
end_W(39, 152) <= 0; end_W(39, 153) <= 0; end_W(39, 154) <= 0; end_W(39, 155) <= 0; end_W(39, 156) <= 0; end_W(39, 157) <= 0; end_W(39, 158) <= 0; end_W(39, 159) <= 0; 
end_W(39, 160) <= 0; end_W(39, 161) <= 0; end_W(39, 162) <= 0; end_W(39, 163) <= 0; end_W(39, 164) <= 0; end_W(39, 165) <= 0; end_W(39, 166) <= 0; end_W(39, 167) <= 0; 
end_W(39, 168) <= 0; end_W(39, 169) <= 0; end_W(39, 170) <= 0; end_W(39, 171) <= 0; end_W(39, 172) <= 0; end_W(39, 173) <= 0; end_W(39, 174) <= 0; end_W(39, 175) <= 0; 
end_W(39, 176) <= 0; end_W(39, 177) <= 0; end_W(39, 178) <= 0; end_W(39, 179) <= 0; end_W(39, 180) <= 0; end_W(39, 181) <= 0; end_W(39, 182) <= 0; end_W(39, 183) <= 0; 
end_W(39, 184) <= 1; end_W(39, 185) <= 1; end_W(39, 186) <= 1; end_W(39, 187) <= 1; end_W(39, 188) <= 1; end_W(39, 189) <= 1; end_W(39, 190) <= 1; end_W(39, 191) <= 1; 
end_W(39, 192) <= 1; end_W(39, 193) <= 1; end_W(39, 194) <= 1; end_W(39, 195) <= 1; end_W(39, 196) <= 1; end_W(39, 197) <= 1; end_W(39, 198) <= 1; end_W(39, 199) <= 1; 
end_W(39, 200) <= 1; end_W(39, 201) <= 1; end_W(39, 202) <= 1; end_W(39, 203) <= 1; end_W(39, 204) <= 0; end_W(39, 205) <= 0; end_W(39, 206) <= 0; end_W(39, 207) <= 0; 
end_W(39, 208) <= 0; end_W(39, 209) <= 0; end_W(39, 210) <= 0; end_W(39, 211) <= 0; end_W(39, 212) <= 0; end_W(39, 213) <= 0; end_W(39, 214) <= 0; end_W(39, 215) <= 0; 
end_W(39, 216) <= 0; end_W(39, 217) <= 0; end_W(39, 218) <= 0; end_W(39, 219) <= 0; end_W(39, 220) <= 0; end_W(39, 221) <= 0; end_W(39, 222) <= 0; end_W(39, 223) <= 0; 
end_W(39, 224) <= 0; end_W(39, 225) <= 0; end_W(39, 226) <= 0; end_W(39, 227) <= 0; end_W(39, 228) <= 1; end_W(39, 229) <= 1; end_W(39, 230) <= 1; end_W(39, 231) <= 1; 
end_W(39, 232) <= 1; end_W(39, 233) <= 1; end_W(39, 234) <= 1; end_W(39, 235) <= 1; end_W(39, 236) <= 0; end_W(39, 237) <= 0; end_W(39, 238) <= 0; end_W(39, 239) <= 0; 
end_W(39, 240) <= 0; end_W(39, 241) <= 0; end_W(39, 242) <= 0; end_W(39, 243) <= 0; end_W(39, 244) <= 0; end_W(39, 245) <= 0; end_W(39, 246) <= 0; end_W(39, 247) <= 0; 
end_W(39, 248) <= 0; end_W(39, 249) <= 0; end_W(39, 250) <= 0; end_W(39, 251) <= 0; end_W(39, 252) <= 1; end_W(39, 253) <= 1; end_W(39, 254) <= 1; end_W(39, 255) <= 1; 
end_W(39, 256) <= 1; end_W(39, 257) <= 1; end_W(39, 258) <= 1; end_W(39, 259) <= 1; end_W(39, 260) <= 1; end_W(39, 261) <= 1; end_W(39, 262) <= 1; end_W(39, 263) <= 1; 
end_W(39, 264) <= 1; end_W(39, 265) <= 1; end_W(39, 266) <= 1; end_W(39, 267) <= 1; end_W(39, 268) <= 1; end_W(39, 269) <= 1; end_W(39, 270) <= 1; end_W(39, 271) <= 1; 
end_W(39, 272) <= 1; end_W(39, 273) <= 1; end_W(39, 274) <= 1; end_W(39, 275) <= 1; end_W(39, 276) <= 1; end_W(39, 277) <= 1; end_W(39, 278) <= 1; end_W(39, 279) <= 1; 
end_W(39, 280) <= 0; end_W(39, 281) <= 0; end_W(39, 282) <= 0; end_W(39, 283) <= 0; end_W(39, 284) <= 0; end_W(39, 285) <= 0; end_W(39, 286) <= 0; end_W(39, 287) <= 0; 
end_W(39, 288) <= 1; end_W(39, 289) <= 1; end_W(39, 290) <= 1; end_W(39, 291) <= 1; end_W(39, 292) <= 1; end_W(39, 293) <= 1; end_W(39, 294) <= 1; end_W(39, 295) <= 1; 
end_W(39, 296) <= 1; end_W(39, 297) <= 1; end_W(39, 298) <= 1; end_W(39, 299) <= 1; end_W(39, 300) <= 0; end_W(39, 301) <= 0; end_W(39, 302) <= 0; end_W(39, 303) <= 0; 
end_W(39, 304) <= 0; end_W(39, 305) <= 0; end_W(39, 306) <= 0; end_W(39, 307) <= 0; end_W(39, 308) <= 1; end_W(39, 309) <= 1; end_W(39, 310) <= 1; end_W(39, 311) <= 1; 
end_W(39, 312) <= 1; end_W(39, 313) <= 1; end_W(39, 314) <= 1; end_W(39, 315) <= 1; end_W(39, 316) <= 0; end_W(39, 317) <= 0; end_W(39, 318) <= 0; end_W(39, 319) <= 0; 
end_W(39, 320) <= 0; end_W(39, 321) <= 0; end_W(39, 322) <= 0; end_W(39, 323) <= 0; 

end Behavioral;
