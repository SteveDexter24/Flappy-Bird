

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package flappypkg is
    type flappyWord is array (0 to 59, 0 to 593) of integer;
end package;

use work.flappypkg.all;

entity flappy is
    Port (flappy_W: out flappyWord );
end flappy;

architecture Behavioral of flappy is

begin


flappy_W(0, 0) <= 1; flappy_W(0, 1) <= 1; flappy_W(0, 2) <= 1; flappy_W(0, 3) <= 1; flappy_W(0, 4) <= 1; flappy_W(0, 5) <= 1; flappy_W(0, 6) <= 1; flappy_W(0, 7) <= 1; flappy_W(0, 8) <= 1; flappy_W(0, 9) <= 1; flappy_W(0, 10) <= 1; flappy_W(0, 11) <= 1; flappy_W(0, 12) <= 1; flappy_W(0, 13) <= 1; flappy_W(0, 14) <= 1; flappy_W(0, 15) <= 1; flappy_W(0, 16) <= 1; flappy_W(0, 17) <= 1; flappy_W(0, 18) <= 1; flappy_W(0, 19) <= 1; flappy_W(0, 20) <= 1; flappy_W(0, 21) <= 1; flappy_W(0, 22) <= 1; flappy_W(0, 23) <= 1; flappy_W(0, 24) <= 1; flappy_W(0, 25) <= 1; flappy_W(0, 26) <= 1; flappy_W(0, 27) <= 1; flappy_W(0, 28) <= 1; flappy_W(0, 29) <= 1; flappy_W(0, 30) <= 1; flappy_W(0, 31) <= 1; flappy_W(0, 32) <= 1; flappy_W(0, 33) <= 1; flappy_W(0, 34) <= 1; flappy_W(0, 35) <= 1; flappy_W(0, 36) <= 1; flappy_W(0, 37) <= 1; flappy_W(0, 38) <= 1; flappy_W(0, 39) <= 1; flappy_W(0, 40) <= 1; flappy_W(0, 41) <= 1; flappy_W(0, 42) <= 0; flappy_W(0, 43) <= 0; flappy_W(0, 44) <= 0; flappy_W(0, 45) <= 0; flappy_W(0, 46) <= 0; flappy_W(0, 47) <= 0; flappy_W(0, 48) <= 0; flappy_W(0, 49) <= 0; flappy_W(0, 50) <= 0; flappy_W(0, 51) <= 0; flappy_W(0, 52) <= 0; flappy_W(0, 53) <= 0; flappy_W(0, 54) <= 1; flappy_W(0, 55) <= 1; flappy_W(0, 56) <= 1; flappy_W(0, 57) <= 1; flappy_W(0, 58) <= 1; flappy_W(0, 59) <= 1; flappy_W(0, 60) <= 1; flappy_W(0, 61) <= 1; flappy_W(0, 62) <= 1; flappy_W(0, 63) <= 1; flappy_W(0, 64) <= 1; flappy_W(0, 65) <= 1; flappy_W(0, 66) <= 1; flappy_W(0, 67) <= 1; flappy_W(0, 68) <= 1; flappy_W(0, 69) <= 1; flappy_W(0, 70) <= 1; flappy_W(0, 71) <= 1; flappy_W(0, 72) <= 1; flappy_W(0, 73) <= 1; flappy_W(0, 74) <= 1; flappy_W(0, 75) <= 1; flappy_W(0, 76) <= 1; flappy_W(0, 77) <= 1; flappy_W(0, 78) <= 0; flappy_W(0, 79) <= 0; flappy_W(0, 80) <= 0; flappy_W(0, 81) <= 0; flappy_W(0, 82) <= 0; flappy_W(0, 83) <= 0; flappy_W(0, 84) <= 0; flappy_W(0, 85) <= 0; flappy_W(0, 86) <= 0; flappy_W(0, 87) <= 0; flappy_W(0, 88) <= 0; flappy_W(0, 89) <= 0; flappy_W(0, 90) <= 0; flappy_W(0, 91) <= 0; flappy_W(0, 92) <= 0; flappy_W(0, 93) <= 0; flappy_W(0, 94) <= 0; flappy_W(0, 95) <= 0; flappy_W(0, 96) <= 0; flappy_W(0, 97) <= 0; flappy_W(0, 98) <= 0; flappy_W(0, 99) <= 0; flappy_W(0, 100) <= 0; flappy_W(0, 101) <= 0; flappy_W(0, 102) <= 0; flappy_W(0, 103) <= 0; flappy_W(0, 104) <= 0; flappy_W(0, 105) <= 0; flappy_W(0, 106) <= 0; flappy_W(0, 107) <= 0; flappy_W(0, 108) <= 0; flappy_W(0, 109) <= 0; flappy_W(0, 110) <= 0; flappy_W(0, 111) <= 0; flappy_W(0, 112) <= 0; flappy_W(0, 113) <= 0; flappy_W(0, 114) <= 0; flappy_W(0, 115) <= 0; flappy_W(0, 116) <= 0; flappy_W(0, 117) <= 0; flappy_W(0, 118) <= 0; flappy_W(0, 119) <= 0; flappy_W(0, 120) <= 0; flappy_W(0, 121) <= 0; flappy_W(0, 122) <= 0; flappy_W(0, 123) <= 0; flappy_W(0, 124) <= 0; flappy_W(0, 125) <= 0; flappy_W(0, 126) <= 1; flappy_W(0, 127) <= 1; flappy_W(0, 128) <= 1; flappy_W(0, 129) <= 1; flappy_W(0, 130) <= 1; flappy_W(0, 131) <= 1; flappy_W(0, 132) <= 0; flappy_W(0, 133) <= 0; flappy_W(0, 134) <= 0; flappy_W(0, 135) <= 0; flappy_W(0, 136) <= 0; flappy_W(0, 137) <= 0; flappy_W(0, 138) <= 0; flappy_W(0, 139) <= 0; flappy_W(0, 140) <= 0; flappy_W(0, 141) <= 0; flappy_W(0, 142) <= 0; flappy_W(0, 143) <= 0; flappy_W(0, 144) <= 0; flappy_W(0, 145) <= 0; flappy_W(0, 146) <= 0; flappy_W(0, 147) <= 0; flappy_W(0, 148) <= 0; flappy_W(0, 149) <= 0; flappy_W(0, 150) <= 0; flappy_W(0, 151) <= 0; flappy_W(0, 152) <= 0; flappy_W(0, 153) <= 0; flappy_W(0, 154) <= 0; flappy_W(0, 155) <= 0; flappy_W(0, 156) <= 0; flappy_W(0, 157) <= 0; flappy_W(0, 158) <= 0; flappy_W(0, 159) <= 0; flappy_W(0, 160) <= 0; flappy_W(0, 161) <= 0; flappy_W(0, 162) <= 1; flappy_W(0, 163) <= 1; flappy_W(0, 164) <= 1; flappy_W(0, 165) <= 1; flappy_W(0, 166) <= 1; flappy_W(0, 167) <= 1; flappy_W(0, 168) <= 1; flappy_W(0, 169) <= 1; flappy_W(0, 170) <= 1; flappy_W(0, 171) <= 1; flappy_W(0, 172) <= 1; flappy_W(0, 173) <= 1; flappy_W(0, 174) <= 1; flappy_W(0, 175) <= 1; flappy_W(0, 176) <= 1; flappy_W(0, 177) <= 1; flappy_W(0, 178) <= 1; flappy_W(0, 179) <= 1; flappy_W(0, 180) <= 1; flappy_W(0, 181) <= 1; flappy_W(0, 182) <= 1; flappy_W(0, 183) <= 1; flappy_W(0, 184) <= 1; flappy_W(0, 185) <= 1; flappy_W(0, 186) <= 1; flappy_W(0, 187) <= 1; flappy_W(0, 188) <= 1; flappy_W(0, 189) <= 1; flappy_W(0, 190) <= 1; flappy_W(0, 191) <= 1; flappy_W(0, 192) <= 1; flappy_W(0, 193) <= 1; flappy_W(0, 194) <= 1; flappy_W(0, 195) <= 1; flappy_W(0, 196) <= 1; flappy_W(0, 197) <= 1; flappy_W(0, 198) <= 0; flappy_W(0, 199) <= 0; flappy_W(0, 200) <= 0; flappy_W(0, 201) <= 0; flappy_W(0, 202) <= 0; flappy_W(0, 203) <= 0; flappy_W(0, 204) <= 0; flappy_W(0, 205) <= 0; flappy_W(0, 206) <= 0; flappy_W(0, 207) <= 0; flappy_W(0, 208) <= 0; flappy_W(0, 209) <= 0; flappy_W(0, 210) <= 0; flappy_W(0, 211) <= 0; flappy_W(0, 212) <= 0; flappy_W(0, 213) <= 0; flappy_W(0, 214) <= 0; flappy_W(0, 215) <= 0; flappy_W(0, 216) <= 1; flappy_W(0, 217) <= 1; flappy_W(0, 218) <= 1; flappy_W(0, 219) <= 1; flappy_W(0, 220) <= 1; flappy_W(0, 221) <= 1; flappy_W(0, 222) <= 1; flappy_W(0, 223) <= 1; flappy_W(0, 224) <= 1; flappy_W(0, 225) <= 1; flappy_W(0, 226) <= 1; flappy_W(0, 227) <= 1; flappy_W(0, 228) <= 1; flappy_W(0, 229) <= 1; flappy_W(0, 230) <= 1; flappy_W(0, 231) <= 1; flappy_W(0, 232) <= 1; flappy_W(0, 233) <= 1; flappy_W(0, 234) <= 1; flappy_W(0, 235) <= 1; flappy_W(0, 236) <= 1; flappy_W(0, 237) <= 1; flappy_W(0, 238) <= 1; flappy_W(0, 239) <= 1; flappy_W(0, 240) <= 1; flappy_W(0, 241) <= 1; flappy_W(0, 242) <= 1; flappy_W(0, 243) <= 1; flappy_W(0, 244) <= 1; flappy_W(0, 245) <= 1; flappy_W(0, 246) <= 1; flappy_W(0, 247) <= 1; flappy_W(0, 248) <= 1; flappy_W(0, 249) <= 1; flappy_W(0, 250) <= 1; flappy_W(0, 251) <= 1; flappy_W(0, 252) <= 0; flappy_W(0, 253) <= 0; flappy_W(0, 254) <= 0; flappy_W(0, 255) <= 0; flappy_W(0, 256) <= 0; flappy_W(0, 257) <= 0; flappy_W(0, 258) <= 0; flappy_W(0, 259) <= 0; flappy_W(0, 260) <= 0; flappy_W(0, 261) <= 0; flappy_W(0, 262) <= 0; flappy_W(0, 263) <= 0; flappy_W(0, 264) <= 0; flappy_W(0, 265) <= 0; flappy_W(0, 266) <= 0; flappy_W(0, 267) <= 0; flappy_W(0, 268) <= 0; flappy_W(0, 269) <= 0; flappy_W(0, 270) <= 1; flappy_W(0, 271) <= 1; flappy_W(0, 272) <= 1; flappy_W(0, 273) <= 1; flappy_W(0, 274) <= 1; flappy_W(0, 275) <= 1; flappy_W(0, 276) <= 1; flappy_W(0, 277) <= 1; flappy_W(0, 278) <= 1; flappy_W(0, 279) <= 1; flappy_W(0, 280) <= 1; flappy_W(0, 281) <= 1; flappy_W(0, 282) <= 0; flappy_W(0, 283) <= 0; flappy_W(0, 284) <= 0; flappy_W(0, 285) <= 0; flappy_W(0, 286) <= 0; flappy_W(0, 287) <= 0; flappy_W(0, 288) <= 0; flappy_W(0, 289) <= 0; flappy_W(0, 290) <= 0; flappy_W(0, 291) <= 0; flappy_W(0, 292) <= 0; flappy_W(0, 293) <= 0; flappy_W(0, 294) <= 0; flappy_W(0, 295) <= 0; flappy_W(0, 296) <= 0; flappy_W(0, 297) <= 0; flappy_W(0, 298) <= 0; flappy_W(0, 299) <= 0; flappy_W(0, 300) <= 0; flappy_W(0, 301) <= 0; flappy_W(0, 302) <= 0; flappy_W(0, 303) <= 0; flappy_W(0, 304) <= 0; flappy_W(0, 305) <= 0; flappy_W(0, 306) <= 1; flappy_W(0, 307) <= 1; flappy_W(0, 308) <= 1; flappy_W(0, 309) <= 1; flappy_W(0, 310) <= 1; flappy_W(0, 311) <= 1; flappy_W(0, 312) <= 1; flappy_W(0, 313) <= 1; flappy_W(0, 314) <= 1; flappy_W(0, 315) <= 1; flappy_W(0, 316) <= 1; flappy_W(0, 317) <= 1; flappy_W(0, 318) <= 0; flappy_W(0, 319) <= 0; flappy_W(0, 320) <= 0; flappy_W(0, 321) <= 0; flappy_W(0, 322) <= 0; flappy_W(0, 323) <= 0; flappy_W(0, 324) <= 0; flappy_W(0, 325) <= 0; flappy_W(0, 326) <= 0; flappy_W(0, 327) <= 0; flappy_W(0, 328) <= 0; flappy_W(0, 329) <= 0; flappy_W(0, 330) <= 0; flappy_W(0, 331) <= 0; flappy_W(0, 332) <= 0; flappy_W(0, 333) <= 0; flappy_W(0, 334) <= 0; flappy_W(0, 335) <= 0; flappy_W(0, 336) <= 0; flappy_W(0, 337) <= 0; flappy_W(0, 338) <= 0; flappy_W(0, 339) <= 0; flappy_W(0, 340) <= 0; flappy_W(0, 341) <= 0; flappy_W(0, 342) <= 0; flappy_W(0, 343) <= 0; flappy_W(0, 344) <= 0; flappy_W(0, 345) <= 0; flappy_W(0, 346) <= 0; flappy_W(0, 347) <= 0; flappy_W(0, 348) <= 0; flappy_W(0, 349) <= 0; flappy_W(0, 350) <= 0; flappy_W(0, 351) <= 0; flappy_W(0, 352) <= 0; flappy_W(0, 353) <= 0; flappy_W(0, 354) <= 0; flappy_W(0, 355) <= 0; flappy_W(0, 356) <= 0; flappy_W(0, 357) <= 0; flappy_W(0, 358) <= 0; flappy_W(0, 359) <= 0; flappy_W(0, 360) <= 0; flappy_W(0, 361) <= 0; flappy_W(0, 362) <= 0; flappy_W(0, 363) <= 0; flappy_W(0, 364) <= 0; flappy_W(0, 365) <= 0; flappy_W(0, 366) <= 0; flappy_W(0, 367) <= 0; flappy_W(0, 368) <= 0; flappy_W(0, 369) <= 0; flappy_W(0, 370) <= 0; flappy_W(0, 371) <= 0; flappy_W(0, 372) <= 0; flappy_W(0, 373) <= 0; flappy_W(0, 374) <= 0; flappy_W(0, 375) <= 0; flappy_W(0, 376) <= 0; flappy_W(0, 377) <= 0; flappy_W(0, 378) <= 0; flappy_W(0, 379) <= 0; flappy_W(0, 380) <= 0; flappy_W(0, 381) <= 0; flappy_W(0, 382) <= 0; flappy_W(0, 383) <= 0; flappy_W(0, 384) <= 0; flappy_W(0, 385) <= 0; flappy_W(0, 386) <= 0; flappy_W(0, 387) <= 0; flappy_W(0, 388) <= 0; flappy_W(0, 389) <= 0; flappy_W(0, 390) <= 0; flappy_W(0, 391) <= 0; flappy_W(0, 392) <= 0; flappy_W(0, 393) <= 0; flappy_W(0, 394) <= 0; flappy_W(0, 395) <= 0; flappy_W(0, 396) <= 1; flappy_W(0, 397) <= 1; flappy_W(0, 398) <= 1; flappy_W(0, 399) <= 1; flappy_W(0, 400) <= 1; flappy_W(0, 401) <= 1; flappy_W(0, 402) <= 1; flappy_W(0, 403) <= 1; flappy_W(0, 404) <= 1; flappy_W(0, 405) <= 1; flappy_W(0, 406) <= 1; flappy_W(0, 407) <= 1; flappy_W(0, 408) <= 1; flappy_W(0, 409) <= 1; flappy_W(0, 410) <= 1; flappy_W(0, 411) <= 1; flappy_W(0, 412) <= 1; flappy_W(0, 413) <= 1; flappy_W(0, 414) <= 1; flappy_W(0, 415) <= 1; flappy_W(0, 416) <= 1; flappy_W(0, 417) <= 1; flappy_W(0, 418) <= 1; flappy_W(0, 419) <= 1; flappy_W(0, 420) <= 1; flappy_W(0, 421) <= 1; flappy_W(0, 422) <= 1; flappy_W(0, 423) <= 1; flappy_W(0, 424) <= 1; flappy_W(0, 425) <= 1; flappy_W(0, 426) <= 1; flappy_W(0, 427) <= 1; flappy_W(0, 428) <= 1; flappy_W(0, 429) <= 1; flappy_W(0, 430) <= 1; flappy_W(0, 431) <= 1; flappy_W(0, 432) <= 0; flappy_W(0, 433) <= 0; flappy_W(0, 434) <= 0; flappy_W(0, 435) <= 0; flappy_W(0, 436) <= 0; flappy_W(0, 437) <= 0; flappy_W(0, 438) <= 0; flappy_W(0, 439) <= 0; flappy_W(0, 440) <= 0; flappy_W(0, 441) <= 0; flappy_W(0, 442) <= 0; flappy_W(0, 443) <= 0; flappy_W(0, 444) <= 0; flappy_W(0, 445) <= 0; flappy_W(0, 446) <= 0; flappy_W(0, 447) <= 0; flappy_W(0, 448) <= 0; flappy_W(0, 449) <= 0; flappy_W(0, 450) <= 0; flappy_W(0, 451) <= 0; flappy_W(0, 452) <= 0; flappy_W(0, 453) <= 0; flappy_W(0, 454) <= 0; flappy_W(0, 455) <= 0; flappy_W(0, 456) <= 0; flappy_W(0, 457) <= 0; flappy_W(0, 458) <= 0; flappy_W(0, 459) <= 0; flappy_W(0, 460) <= 0; flappy_W(0, 461) <= 0; flappy_W(0, 462) <= 1; flappy_W(0, 463) <= 1; flappy_W(0, 464) <= 1; flappy_W(0, 465) <= 1; flappy_W(0, 466) <= 1; flappy_W(0, 467) <= 1; flappy_W(0, 468) <= 1; flappy_W(0, 469) <= 1; flappy_W(0, 470) <= 1; flappy_W(0, 471) <= 1; flappy_W(0, 472) <= 1; flappy_W(0, 473) <= 1; flappy_W(0, 474) <= 1; flappy_W(0, 475) <= 1; flappy_W(0, 476) <= 1; flappy_W(0, 477) <= 1; flappy_W(0, 478) <= 1; flappy_W(0, 479) <= 1; flappy_W(0, 480) <= 1; flappy_W(0, 481) <= 1; flappy_W(0, 482) <= 1; flappy_W(0, 483) <= 1; flappy_W(0, 484) <= 1; flappy_W(0, 485) <= 1; flappy_W(0, 486) <= 0; flappy_W(0, 487) <= 0; flappy_W(0, 488) <= 0; flappy_W(0, 489) <= 0; flappy_W(0, 490) <= 0; flappy_W(0, 491) <= 0; flappy_W(0, 492) <= 0; flappy_W(0, 493) <= 0; flappy_W(0, 494) <= 0; flappy_W(0, 495) <= 0; flappy_W(0, 496) <= 0; flappy_W(0, 497) <= 0; flappy_W(0, 498) <= 0; flappy_W(0, 499) <= 0; flappy_W(0, 500) <= 0; flappy_W(0, 501) <= 0; flappy_W(0, 502) <= 0; flappy_W(0, 503) <= 0; flappy_W(0, 504) <= 1; flappy_W(0, 505) <= 1; flappy_W(0, 506) <= 1; flappy_W(0, 507) <= 1; flappy_W(0, 508) <= 1; flappy_W(0, 509) <= 1; flappy_W(0, 510) <= 1; flappy_W(0, 511) <= 1; flappy_W(0, 512) <= 1; flappy_W(0, 513) <= 1; flappy_W(0, 514) <= 1; flappy_W(0, 515) <= 1; flappy_W(0, 516) <= 1; flappy_W(0, 517) <= 1; flappy_W(0, 518) <= 1; flappy_W(0, 519) <= 1; flappy_W(0, 520) <= 1; flappy_W(0, 521) <= 1; flappy_W(0, 522) <= 1; flappy_W(0, 523) <= 1; flappy_W(0, 524) <= 1; flappy_W(0, 525) <= 1; flappy_W(0, 526) <= 1; flappy_W(0, 527) <= 1; flappy_W(0, 528) <= 1; flappy_W(0, 529) <= 1; flappy_W(0, 530) <= 1; flappy_W(0, 531) <= 1; flappy_W(0, 532) <= 1; flappy_W(0, 533) <= 1; flappy_W(0, 534) <= 1; flappy_W(0, 535) <= 1; flappy_W(0, 536) <= 1; flappy_W(0, 537) <= 1; flappy_W(0, 538) <= 1; flappy_W(0, 539) <= 1; flappy_W(0, 540) <= 0; flappy_W(0, 541) <= 0; flappy_W(0, 542) <= 0; flappy_W(0, 543) <= 0; flappy_W(0, 544) <= 0; flappy_W(0, 545) <= 0; flappy_W(0, 546) <= 0; flappy_W(0, 547) <= 0; flappy_W(0, 548) <= 0; flappy_W(0, 549) <= 0; flappy_W(0, 550) <= 0; flappy_W(0, 551) <= 0; flappy_W(0, 552) <= 0; flappy_W(0, 553) <= 0; flappy_W(0, 554) <= 0; flappy_W(0, 555) <= 0; flappy_W(0, 556) <= 0; flappy_W(0, 557) <= 0; flappy_W(0, 558) <= 1; flappy_W(0, 559) <= 1; flappy_W(0, 560) <= 1; flappy_W(0, 561) <= 1; flappy_W(0, 562) <= 1; flappy_W(0, 563) <= 1; flappy_W(0, 564) <= 1; flappy_W(0, 565) <= 1; flappy_W(0, 566) <= 1; flappy_W(0, 567) <= 1; flappy_W(0, 568) <= 1; flappy_W(0, 569) <= 1; flappy_W(0, 570) <= 1; flappy_W(0, 571) <= 1; flappy_W(0, 572) <= 1; flappy_W(0, 573) <= 1; flappy_W(0, 574) <= 1; flappy_W(0, 575) <= 1; flappy_W(0, 576) <= 1; flappy_W(0, 577) <= 1; flappy_W(0, 578) <= 1; flappy_W(0, 579) <= 1; flappy_W(0, 580) <= 1; flappy_W(0, 581) <= 1; flappy_W(0, 582) <= 1; flappy_W(0, 583) <= 1; flappy_W(0, 584) <= 1; flappy_W(0, 585) <= 1; flappy_W(0, 586) <= 1; flappy_W(0, 587) <= 1; flappy_W(0, 588) <= 0; flappy_W(0, 589) <= 0; flappy_W(0, 590) <= 0; flappy_W(0, 591) <= 0; flappy_W(0, 592) <= 0; flappy_W(0, 593) <= 0; 
flappy_W(1, 0) <= 1; flappy_W(1, 1) <= 1; flappy_W(1, 2) <= 1; flappy_W(1, 3) <= 1; flappy_W(1, 4) <= 1; flappy_W(1, 5) <= 1; flappy_W(1, 6) <= 1; flappy_W(1, 7) <= 1; flappy_W(1, 8) <= 1; flappy_W(1, 9) <= 1; flappy_W(1, 10) <= 1; flappy_W(1, 11) <= 1; flappy_W(1, 12) <= 1; flappy_W(1, 13) <= 1; flappy_W(1, 14) <= 1; flappy_W(1, 15) <= 1; flappy_W(1, 16) <= 1; flappy_W(1, 17) <= 1; flappy_W(1, 18) <= 1; flappy_W(1, 19) <= 1; flappy_W(1, 20) <= 1; flappy_W(1, 21) <= 1; flappy_W(1, 22) <= 1; flappy_W(1, 23) <= 1; flappy_W(1, 24) <= 1; flappy_W(1, 25) <= 1; flappy_W(1, 26) <= 1; flappy_W(1, 27) <= 1; flappy_W(1, 28) <= 1; flappy_W(1, 29) <= 1; flappy_W(1, 30) <= 1; flappy_W(1, 31) <= 1; flappy_W(1, 32) <= 1; flappy_W(1, 33) <= 1; flappy_W(1, 34) <= 1; flappy_W(1, 35) <= 1; flappy_W(1, 36) <= 1; flappy_W(1, 37) <= 1; flappy_W(1, 38) <= 1; flappy_W(1, 39) <= 1; flappy_W(1, 40) <= 1; flappy_W(1, 41) <= 1; flappy_W(1, 42) <= 0; flappy_W(1, 43) <= 0; flappy_W(1, 44) <= 0; flappy_W(1, 45) <= 0; flappy_W(1, 46) <= 0; flappy_W(1, 47) <= 0; flappy_W(1, 48) <= 0; flappy_W(1, 49) <= 0; flappy_W(1, 50) <= 0; flappy_W(1, 51) <= 0; flappy_W(1, 52) <= 0; flappy_W(1, 53) <= 0; flappy_W(1, 54) <= 1; flappy_W(1, 55) <= 1; flappy_W(1, 56) <= 1; flappy_W(1, 57) <= 1; flappy_W(1, 58) <= 1; flappy_W(1, 59) <= 1; flappy_W(1, 60) <= 1; flappy_W(1, 61) <= 1; flappy_W(1, 62) <= 1; flappy_W(1, 63) <= 1; flappy_W(1, 64) <= 1; flappy_W(1, 65) <= 1; flappy_W(1, 66) <= 1; flappy_W(1, 67) <= 1; flappy_W(1, 68) <= 1; flappy_W(1, 69) <= 1; flappy_W(1, 70) <= 1; flappy_W(1, 71) <= 1; flappy_W(1, 72) <= 1; flappy_W(1, 73) <= 1; flappy_W(1, 74) <= 1; flappy_W(1, 75) <= 1; flappy_W(1, 76) <= 1; flappy_W(1, 77) <= 1; flappy_W(1, 78) <= 0; flappy_W(1, 79) <= 0; flappy_W(1, 80) <= 0; flappy_W(1, 81) <= 0; flappy_W(1, 82) <= 0; flappy_W(1, 83) <= 0; flappy_W(1, 84) <= 0; flappy_W(1, 85) <= 0; flappy_W(1, 86) <= 0; flappy_W(1, 87) <= 0; flappy_W(1, 88) <= 0; flappy_W(1, 89) <= 0; flappy_W(1, 90) <= 0; flappy_W(1, 91) <= 0; flappy_W(1, 92) <= 0; flappy_W(1, 93) <= 0; flappy_W(1, 94) <= 0; flappy_W(1, 95) <= 0; flappy_W(1, 96) <= 0; flappy_W(1, 97) <= 0; flappy_W(1, 98) <= 0; flappy_W(1, 99) <= 0; flappy_W(1, 100) <= 0; flappy_W(1, 101) <= 0; flappy_W(1, 102) <= 0; flappy_W(1, 103) <= 0; flappy_W(1, 104) <= 0; flappy_W(1, 105) <= 0; flappy_W(1, 106) <= 0; flappy_W(1, 107) <= 0; flappy_W(1, 108) <= 0; flappy_W(1, 109) <= 0; flappy_W(1, 110) <= 0; flappy_W(1, 111) <= 0; flappy_W(1, 112) <= 0; flappy_W(1, 113) <= 0; flappy_W(1, 114) <= 0; flappy_W(1, 115) <= 0; flappy_W(1, 116) <= 0; flappy_W(1, 117) <= 0; flappy_W(1, 118) <= 0; flappy_W(1, 119) <= 0; flappy_W(1, 120) <= 0; flappy_W(1, 121) <= 0; flappy_W(1, 122) <= 0; flappy_W(1, 123) <= 0; flappy_W(1, 124) <= 0; flappy_W(1, 125) <= 0; flappy_W(1, 126) <= 1; flappy_W(1, 127) <= 1; flappy_W(1, 128) <= 1; flappy_W(1, 129) <= 1; flappy_W(1, 130) <= 1; flappy_W(1, 131) <= 1; flappy_W(1, 132) <= 0; flappy_W(1, 133) <= 0; flappy_W(1, 134) <= 0; flappy_W(1, 135) <= 0; flappy_W(1, 136) <= 0; flappy_W(1, 137) <= 0; flappy_W(1, 138) <= 0; flappy_W(1, 139) <= 0; flappy_W(1, 140) <= 0; flappy_W(1, 141) <= 0; flappy_W(1, 142) <= 0; flappy_W(1, 143) <= 0; flappy_W(1, 144) <= 0; flappy_W(1, 145) <= 0; flappy_W(1, 146) <= 0; flappy_W(1, 147) <= 0; flappy_W(1, 148) <= 0; flappy_W(1, 149) <= 0; flappy_W(1, 150) <= 0; flappy_W(1, 151) <= 0; flappy_W(1, 152) <= 0; flappy_W(1, 153) <= 0; flappy_W(1, 154) <= 0; flappy_W(1, 155) <= 0; flappy_W(1, 156) <= 0; flappy_W(1, 157) <= 0; flappy_W(1, 158) <= 0; flappy_W(1, 159) <= 0; flappy_W(1, 160) <= 0; flappy_W(1, 161) <= 0; flappy_W(1, 162) <= 1; flappy_W(1, 163) <= 1; flappy_W(1, 164) <= 1; flappy_W(1, 165) <= 1; flappy_W(1, 166) <= 1; flappy_W(1, 167) <= 1; flappy_W(1, 168) <= 1; flappy_W(1, 169) <= 1; flappy_W(1, 170) <= 1; flappy_W(1, 171) <= 1; flappy_W(1, 172) <= 1; flappy_W(1, 173) <= 1; flappy_W(1, 174) <= 1; flappy_W(1, 175) <= 1; flappy_W(1, 176) <= 1; flappy_W(1, 177) <= 1; flappy_W(1, 178) <= 1; flappy_W(1, 179) <= 1; flappy_W(1, 180) <= 1; flappy_W(1, 181) <= 1; flappy_W(1, 182) <= 1; flappy_W(1, 183) <= 1; flappy_W(1, 184) <= 1; flappy_W(1, 185) <= 1; flappy_W(1, 186) <= 1; flappy_W(1, 187) <= 1; flappy_W(1, 188) <= 1; flappy_W(1, 189) <= 1; flappy_W(1, 190) <= 1; flappy_W(1, 191) <= 1; flappy_W(1, 192) <= 1; flappy_W(1, 193) <= 1; flappy_W(1, 194) <= 1; flappy_W(1, 195) <= 1; flappy_W(1, 196) <= 1; flappy_W(1, 197) <= 1; flappy_W(1, 198) <= 0; flappy_W(1, 199) <= 0; flappy_W(1, 200) <= 0; flappy_W(1, 201) <= 0; flappy_W(1, 202) <= 0; flappy_W(1, 203) <= 0; flappy_W(1, 204) <= 0; flappy_W(1, 205) <= 0; flappy_W(1, 206) <= 0; flappy_W(1, 207) <= 0; flappy_W(1, 208) <= 0; flappy_W(1, 209) <= 0; flappy_W(1, 210) <= 0; flappy_W(1, 211) <= 0; flappy_W(1, 212) <= 0; flappy_W(1, 213) <= 0; flappy_W(1, 214) <= 0; flappy_W(1, 215) <= 0; flappy_W(1, 216) <= 1; flappy_W(1, 217) <= 1; flappy_W(1, 218) <= 1; flappy_W(1, 219) <= 1; flappy_W(1, 220) <= 1; flappy_W(1, 221) <= 1; flappy_W(1, 222) <= 1; flappy_W(1, 223) <= 1; flappy_W(1, 224) <= 1; flappy_W(1, 225) <= 1; flappy_W(1, 226) <= 1; flappy_W(1, 227) <= 1; flappy_W(1, 228) <= 1; flappy_W(1, 229) <= 1; flappy_W(1, 230) <= 1; flappy_W(1, 231) <= 1; flappy_W(1, 232) <= 1; flappy_W(1, 233) <= 1; flappy_W(1, 234) <= 1; flappy_W(1, 235) <= 1; flappy_W(1, 236) <= 1; flappy_W(1, 237) <= 1; flappy_W(1, 238) <= 1; flappy_W(1, 239) <= 1; flappy_W(1, 240) <= 1; flappy_W(1, 241) <= 1; flappy_W(1, 242) <= 1; flappy_W(1, 243) <= 1; flappy_W(1, 244) <= 1; flappy_W(1, 245) <= 1; flappy_W(1, 246) <= 1; flappy_W(1, 247) <= 1; flappy_W(1, 248) <= 1; flappy_W(1, 249) <= 1; flappy_W(1, 250) <= 1; flappy_W(1, 251) <= 1; flappy_W(1, 252) <= 0; flappy_W(1, 253) <= 0; flappy_W(1, 254) <= 0; flappy_W(1, 255) <= 0; flappy_W(1, 256) <= 0; flappy_W(1, 257) <= 0; flappy_W(1, 258) <= 0; flappy_W(1, 259) <= 0; flappy_W(1, 260) <= 0; flappy_W(1, 261) <= 0; flappy_W(1, 262) <= 0; flappy_W(1, 263) <= 0; flappy_W(1, 264) <= 0; flappy_W(1, 265) <= 0; flappy_W(1, 266) <= 0; flappy_W(1, 267) <= 0; flappy_W(1, 268) <= 0; flappy_W(1, 269) <= 0; flappy_W(1, 270) <= 1; flappy_W(1, 271) <= 1; flappy_W(1, 272) <= 1; flappy_W(1, 273) <= 1; flappy_W(1, 274) <= 1; flappy_W(1, 275) <= 1; flappy_W(1, 276) <= 1; flappy_W(1, 277) <= 1; flappy_W(1, 278) <= 1; flappy_W(1, 279) <= 1; flappy_W(1, 280) <= 1; flappy_W(1, 281) <= 1; flappy_W(1, 282) <= 0; flappy_W(1, 283) <= 0; flappy_W(1, 284) <= 0; flappy_W(1, 285) <= 0; flappy_W(1, 286) <= 0; flappy_W(1, 287) <= 0; flappy_W(1, 288) <= 0; flappy_W(1, 289) <= 0; flappy_W(1, 290) <= 0; flappy_W(1, 291) <= 0; flappy_W(1, 292) <= 0; flappy_W(1, 293) <= 0; flappy_W(1, 294) <= 0; flappy_W(1, 295) <= 0; flappy_W(1, 296) <= 0; flappy_W(1, 297) <= 0; flappy_W(1, 298) <= 0; flappy_W(1, 299) <= 0; flappy_W(1, 300) <= 0; flappy_W(1, 301) <= 0; flappy_W(1, 302) <= 0; flappy_W(1, 303) <= 0; flappy_W(1, 304) <= 0; flappy_W(1, 305) <= 0; flappy_W(1, 306) <= 1; flappy_W(1, 307) <= 1; flappy_W(1, 308) <= 1; flappy_W(1, 309) <= 1; flappy_W(1, 310) <= 1; flappy_W(1, 311) <= 1; flappy_W(1, 312) <= 1; flappy_W(1, 313) <= 1; flappy_W(1, 314) <= 1; flappy_W(1, 315) <= 1; flappy_W(1, 316) <= 1; flappy_W(1, 317) <= 1; flappy_W(1, 318) <= 0; flappy_W(1, 319) <= 0; flappy_W(1, 320) <= 0; flappy_W(1, 321) <= 0; flappy_W(1, 322) <= 0; flappy_W(1, 323) <= 0; flappy_W(1, 324) <= 0; flappy_W(1, 325) <= 0; flappy_W(1, 326) <= 0; flappy_W(1, 327) <= 0; flappy_W(1, 328) <= 0; flappy_W(1, 329) <= 0; flappy_W(1, 330) <= 0; flappy_W(1, 331) <= 0; flappy_W(1, 332) <= 0; flappy_W(1, 333) <= 0; flappy_W(1, 334) <= 0; flappy_W(1, 335) <= 0; flappy_W(1, 336) <= 0; flappy_W(1, 337) <= 0; flappy_W(1, 338) <= 0; flappy_W(1, 339) <= 0; flappy_W(1, 340) <= 0; flappy_W(1, 341) <= 0; flappy_W(1, 342) <= 0; flappy_W(1, 343) <= 0; flappy_W(1, 344) <= 0; flappy_W(1, 345) <= 0; flappy_W(1, 346) <= 0; flappy_W(1, 347) <= 0; flappy_W(1, 348) <= 0; flappy_W(1, 349) <= 0; flappy_W(1, 350) <= 0; flappy_W(1, 351) <= 0; flappy_W(1, 352) <= 0; flappy_W(1, 353) <= 0; flappy_W(1, 354) <= 0; flappy_W(1, 355) <= 0; flappy_W(1, 356) <= 0; flappy_W(1, 357) <= 0; flappy_W(1, 358) <= 0; flappy_W(1, 359) <= 0; flappy_W(1, 360) <= 0; flappy_W(1, 361) <= 0; flappy_W(1, 362) <= 0; flappy_W(1, 363) <= 0; flappy_W(1, 364) <= 0; flappy_W(1, 365) <= 0; flappy_W(1, 366) <= 0; flappy_W(1, 367) <= 0; flappy_W(1, 368) <= 0; flappy_W(1, 369) <= 0; flappy_W(1, 370) <= 0; flappy_W(1, 371) <= 0; flappy_W(1, 372) <= 0; flappy_W(1, 373) <= 0; flappy_W(1, 374) <= 0; flappy_W(1, 375) <= 0; flappy_W(1, 376) <= 0; flappy_W(1, 377) <= 0; flappy_W(1, 378) <= 0; flappy_W(1, 379) <= 0; flappy_W(1, 380) <= 0; flappy_W(1, 381) <= 0; flappy_W(1, 382) <= 0; flappy_W(1, 383) <= 0; flappy_W(1, 384) <= 0; flappy_W(1, 385) <= 0; flappy_W(1, 386) <= 0; flappy_W(1, 387) <= 0; flappy_W(1, 388) <= 0; flappy_W(1, 389) <= 0; flappy_W(1, 390) <= 0; flappy_W(1, 391) <= 0; flappy_W(1, 392) <= 0; flappy_W(1, 393) <= 0; flappy_W(1, 394) <= 0; flappy_W(1, 395) <= 0; flappy_W(1, 396) <= 1; flappy_W(1, 397) <= 1; flappy_W(1, 398) <= 1; flappy_W(1, 399) <= 1; flappy_W(1, 400) <= 1; flappy_W(1, 401) <= 1; flappy_W(1, 402) <= 1; flappy_W(1, 403) <= 1; flappy_W(1, 404) <= 1; flappy_W(1, 405) <= 1; flappy_W(1, 406) <= 1; flappy_W(1, 407) <= 1; flappy_W(1, 408) <= 1; flappy_W(1, 409) <= 1; flappy_W(1, 410) <= 1; flappy_W(1, 411) <= 1; flappy_W(1, 412) <= 1; flappy_W(1, 413) <= 1; flappy_W(1, 414) <= 1; flappy_W(1, 415) <= 1; flappy_W(1, 416) <= 1; flappy_W(1, 417) <= 1; flappy_W(1, 418) <= 1; flappy_W(1, 419) <= 1; flappy_W(1, 420) <= 1; flappy_W(1, 421) <= 1; flappy_W(1, 422) <= 1; flappy_W(1, 423) <= 1; flappy_W(1, 424) <= 1; flappy_W(1, 425) <= 1; flappy_W(1, 426) <= 1; flappy_W(1, 427) <= 1; flappy_W(1, 428) <= 1; flappy_W(1, 429) <= 1; flappy_W(1, 430) <= 1; flappy_W(1, 431) <= 1; flappy_W(1, 432) <= 0; flappy_W(1, 433) <= 0; flappy_W(1, 434) <= 0; flappy_W(1, 435) <= 0; flappy_W(1, 436) <= 0; flappy_W(1, 437) <= 0; flappy_W(1, 438) <= 0; flappy_W(1, 439) <= 0; flappy_W(1, 440) <= 0; flappy_W(1, 441) <= 0; flappy_W(1, 442) <= 0; flappy_W(1, 443) <= 0; flappy_W(1, 444) <= 0; flappy_W(1, 445) <= 0; flappy_W(1, 446) <= 0; flappy_W(1, 447) <= 0; flappy_W(1, 448) <= 0; flappy_W(1, 449) <= 0; flappy_W(1, 450) <= 0; flappy_W(1, 451) <= 0; flappy_W(1, 452) <= 0; flappy_W(1, 453) <= 0; flappy_W(1, 454) <= 0; flappy_W(1, 455) <= 0; flappy_W(1, 456) <= 0; flappy_W(1, 457) <= 0; flappy_W(1, 458) <= 0; flappy_W(1, 459) <= 0; flappy_W(1, 460) <= 0; flappy_W(1, 461) <= 0; flappy_W(1, 462) <= 1; flappy_W(1, 463) <= 1; flappy_W(1, 464) <= 1; flappy_W(1, 465) <= 1; flappy_W(1, 466) <= 1; flappy_W(1, 467) <= 1; flappy_W(1, 468) <= 1; flappy_W(1, 469) <= 1; flappy_W(1, 470) <= 1; flappy_W(1, 471) <= 1; flappy_W(1, 472) <= 1; flappy_W(1, 473) <= 1; flappy_W(1, 474) <= 1; flappy_W(1, 475) <= 1; flappy_W(1, 476) <= 1; flappy_W(1, 477) <= 1; flappy_W(1, 478) <= 1; flappy_W(1, 479) <= 1; flappy_W(1, 480) <= 1; flappy_W(1, 481) <= 1; flappy_W(1, 482) <= 1; flappy_W(1, 483) <= 1; flappy_W(1, 484) <= 1; flappy_W(1, 485) <= 1; flappy_W(1, 486) <= 0; flappy_W(1, 487) <= 0; flappy_W(1, 488) <= 0; flappy_W(1, 489) <= 0; flappy_W(1, 490) <= 0; flappy_W(1, 491) <= 0; flappy_W(1, 492) <= 0; flappy_W(1, 493) <= 0; flappy_W(1, 494) <= 0; flappy_W(1, 495) <= 0; flappy_W(1, 496) <= 0; flappy_W(1, 497) <= 0; flappy_W(1, 498) <= 0; flappy_W(1, 499) <= 0; flappy_W(1, 500) <= 0; flappy_W(1, 501) <= 0; flappy_W(1, 502) <= 0; flappy_W(1, 503) <= 0; flappy_W(1, 504) <= 1; flappy_W(1, 505) <= 1; flappy_W(1, 506) <= 1; flappy_W(1, 507) <= 1; flappy_W(1, 508) <= 1; flappy_W(1, 509) <= 1; flappy_W(1, 510) <= 1; flappy_W(1, 511) <= 1; flappy_W(1, 512) <= 1; flappy_W(1, 513) <= 1; flappy_W(1, 514) <= 1; flappy_W(1, 515) <= 1; flappy_W(1, 516) <= 1; flappy_W(1, 517) <= 1; flappy_W(1, 518) <= 1; flappy_W(1, 519) <= 1; flappy_W(1, 520) <= 1; flappy_W(1, 521) <= 1; flappy_W(1, 522) <= 1; flappy_W(1, 523) <= 1; flappy_W(1, 524) <= 1; flappy_W(1, 525) <= 1; flappy_W(1, 526) <= 1; flappy_W(1, 527) <= 1; flappy_W(1, 528) <= 1; flappy_W(1, 529) <= 1; flappy_W(1, 530) <= 1; flappy_W(1, 531) <= 1; flappy_W(1, 532) <= 1; flappy_W(1, 533) <= 1; flappy_W(1, 534) <= 1; flappy_W(1, 535) <= 1; flappy_W(1, 536) <= 1; flappy_W(1, 537) <= 1; flappy_W(1, 538) <= 1; flappy_W(1, 539) <= 1; flappy_W(1, 540) <= 0; flappy_W(1, 541) <= 0; flappy_W(1, 542) <= 0; flappy_W(1, 543) <= 0; flappy_W(1, 544) <= 0; flappy_W(1, 545) <= 0; flappy_W(1, 546) <= 0; flappy_W(1, 547) <= 0; flappy_W(1, 548) <= 0; flappy_W(1, 549) <= 0; flappy_W(1, 550) <= 0; flappy_W(1, 551) <= 0; flappy_W(1, 552) <= 0; flappy_W(1, 553) <= 0; flappy_W(1, 554) <= 0; flappy_W(1, 555) <= 0; flappy_W(1, 556) <= 0; flappy_W(1, 557) <= 0; flappy_W(1, 558) <= 1; flappy_W(1, 559) <= 1; flappy_W(1, 560) <= 1; flappy_W(1, 561) <= 1; flappy_W(1, 562) <= 1; flappy_W(1, 563) <= 1; flappy_W(1, 564) <= 1; flappy_W(1, 565) <= 1; flappy_W(1, 566) <= 1; flappy_W(1, 567) <= 1; flappy_W(1, 568) <= 1; flappy_W(1, 569) <= 1; flappy_W(1, 570) <= 1; flappy_W(1, 571) <= 1; flappy_W(1, 572) <= 1; flappy_W(1, 573) <= 1; flappy_W(1, 574) <= 1; flappy_W(1, 575) <= 1; flappy_W(1, 576) <= 1; flappy_W(1, 577) <= 1; flappy_W(1, 578) <= 1; flappy_W(1, 579) <= 1; flappy_W(1, 580) <= 1; flappy_W(1, 581) <= 1; flappy_W(1, 582) <= 1; flappy_W(1, 583) <= 1; flappy_W(1, 584) <= 1; flappy_W(1, 585) <= 1; flappy_W(1, 586) <= 1; flappy_W(1, 587) <= 1; flappy_W(1, 588) <= 0; flappy_W(1, 589) <= 0; flappy_W(1, 590) <= 0; flappy_W(1, 591) <= 0; flappy_W(1, 592) <= 0; flappy_W(1, 593) <= 0; 
flappy_W(2, 0) <= 1; flappy_W(2, 1) <= 1; flappy_W(2, 2) <= 1; flappy_W(2, 3) <= 1; flappy_W(2, 4) <= 1; flappy_W(2, 5) <= 1; flappy_W(2, 6) <= 1; flappy_W(2, 7) <= 1; flappy_W(2, 8) <= 1; flappy_W(2, 9) <= 1; flappy_W(2, 10) <= 1; flappy_W(2, 11) <= 1; flappy_W(2, 12) <= 1; flappy_W(2, 13) <= 1; flappy_W(2, 14) <= 1; flappy_W(2, 15) <= 1; flappy_W(2, 16) <= 1; flappy_W(2, 17) <= 1; flappy_W(2, 18) <= 1; flappy_W(2, 19) <= 1; flappy_W(2, 20) <= 1; flappy_W(2, 21) <= 1; flappy_W(2, 22) <= 1; flappy_W(2, 23) <= 1; flappy_W(2, 24) <= 1; flappy_W(2, 25) <= 1; flappy_W(2, 26) <= 1; flappy_W(2, 27) <= 1; flappy_W(2, 28) <= 1; flappy_W(2, 29) <= 1; flappy_W(2, 30) <= 1; flappy_W(2, 31) <= 1; flappy_W(2, 32) <= 1; flappy_W(2, 33) <= 1; flappy_W(2, 34) <= 1; flappy_W(2, 35) <= 1; flappy_W(2, 36) <= 1; flappy_W(2, 37) <= 1; flappy_W(2, 38) <= 1; flappy_W(2, 39) <= 1; flappy_W(2, 40) <= 1; flappy_W(2, 41) <= 1; flappy_W(2, 42) <= 0; flappy_W(2, 43) <= 0; flappy_W(2, 44) <= 0; flappy_W(2, 45) <= 0; flappy_W(2, 46) <= 0; flappy_W(2, 47) <= 0; flappy_W(2, 48) <= 0; flappy_W(2, 49) <= 0; flappy_W(2, 50) <= 0; flappy_W(2, 51) <= 0; flappy_W(2, 52) <= 0; flappy_W(2, 53) <= 0; flappy_W(2, 54) <= 1; flappy_W(2, 55) <= 1; flappy_W(2, 56) <= 1; flappy_W(2, 57) <= 1; flappy_W(2, 58) <= 1; flappy_W(2, 59) <= 1; flappy_W(2, 60) <= 1; flappy_W(2, 61) <= 1; flappy_W(2, 62) <= 1; flappy_W(2, 63) <= 1; flappy_W(2, 64) <= 1; flappy_W(2, 65) <= 1; flappy_W(2, 66) <= 1; flappy_W(2, 67) <= 1; flappy_W(2, 68) <= 1; flappy_W(2, 69) <= 1; flappy_W(2, 70) <= 1; flappy_W(2, 71) <= 1; flappy_W(2, 72) <= 1; flappy_W(2, 73) <= 1; flappy_W(2, 74) <= 1; flappy_W(2, 75) <= 1; flappy_W(2, 76) <= 1; flappy_W(2, 77) <= 1; flappy_W(2, 78) <= 0; flappy_W(2, 79) <= 0; flappy_W(2, 80) <= 0; flappy_W(2, 81) <= 0; flappy_W(2, 82) <= 0; flappy_W(2, 83) <= 0; flappy_W(2, 84) <= 0; flappy_W(2, 85) <= 0; flappy_W(2, 86) <= 0; flappy_W(2, 87) <= 0; flappy_W(2, 88) <= 0; flappy_W(2, 89) <= 0; flappy_W(2, 90) <= 0; flappy_W(2, 91) <= 0; flappy_W(2, 92) <= 0; flappy_W(2, 93) <= 0; flappy_W(2, 94) <= 0; flappy_W(2, 95) <= 0; flappy_W(2, 96) <= 0; flappy_W(2, 97) <= 0; flappy_W(2, 98) <= 0; flappy_W(2, 99) <= 0; flappy_W(2, 100) <= 0; flappy_W(2, 101) <= 0; flappy_W(2, 102) <= 0; flappy_W(2, 103) <= 0; flappy_W(2, 104) <= 0; flappy_W(2, 105) <= 0; flappy_W(2, 106) <= 0; flappy_W(2, 107) <= 0; flappy_W(2, 108) <= 0; flappy_W(2, 109) <= 0; flappy_W(2, 110) <= 0; flappy_W(2, 111) <= 0; flappy_W(2, 112) <= 0; flappy_W(2, 113) <= 0; flappy_W(2, 114) <= 0; flappy_W(2, 115) <= 0; flappy_W(2, 116) <= 0; flappy_W(2, 117) <= 0; flappy_W(2, 118) <= 0; flappy_W(2, 119) <= 0; flappy_W(2, 120) <= 0; flappy_W(2, 121) <= 0; flappy_W(2, 122) <= 0; flappy_W(2, 123) <= 0; flappy_W(2, 124) <= 0; flappy_W(2, 125) <= 0; flappy_W(2, 126) <= 1; flappy_W(2, 127) <= 1; flappy_W(2, 128) <= 1; flappy_W(2, 129) <= 1; flappy_W(2, 130) <= 1; flappy_W(2, 131) <= 1; flappy_W(2, 132) <= 0; flappy_W(2, 133) <= 0; flappy_W(2, 134) <= 0; flappy_W(2, 135) <= 0; flappy_W(2, 136) <= 0; flappy_W(2, 137) <= 0; flappy_W(2, 138) <= 0; flappy_W(2, 139) <= 0; flappy_W(2, 140) <= 0; flappy_W(2, 141) <= 0; flappy_W(2, 142) <= 0; flappy_W(2, 143) <= 0; flappy_W(2, 144) <= 0; flappy_W(2, 145) <= 0; flappy_W(2, 146) <= 0; flappy_W(2, 147) <= 0; flappy_W(2, 148) <= 0; flappy_W(2, 149) <= 0; flappy_W(2, 150) <= 0; flappy_W(2, 151) <= 0; flappy_W(2, 152) <= 0; flappy_W(2, 153) <= 0; flappy_W(2, 154) <= 0; flappy_W(2, 155) <= 0; flappy_W(2, 156) <= 0; flappy_W(2, 157) <= 0; flappy_W(2, 158) <= 0; flappy_W(2, 159) <= 0; flappy_W(2, 160) <= 0; flappy_W(2, 161) <= 0; flappy_W(2, 162) <= 1; flappy_W(2, 163) <= 1; flappy_W(2, 164) <= 1; flappy_W(2, 165) <= 1; flappy_W(2, 166) <= 1; flappy_W(2, 167) <= 1; flappy_W(2, 168) <= 1; flappy_W(2, 169) <= 1; flappy_W(2, 170) <= 1; flappy_W(2, 171) <= 1; flappy_W(2, 172) <= 1; flappy_W(2, 173) <= 1; flappy_W(2, 174) <= 1; flappy_W(2, 175) <= 1; flappy_W(2, 176) <= 1; flappy_W(2, 177) <= 1; flappy_W(2, 178) <= 1; flappy_W(2, 179) <= 1; flappy_W(2, 180) <= 1; flappy_W(2, 181) <= 1; flappy_W(2, 182) <= 1; flappy_W(2, 183) <= 1; flappy_W(2, 184) <= 1; flappy_W(2, 185) <= 1; flappy_W(2, 186) <= 1; flappy_W(2, 187) <= 1; flappy_W(2, 188) <= 1; flappy_W(2, 189) <= 1; flappy_W(2, 190) <= 1; flappy_W(2, 191) <= 1; flappy_W(2, 192) <= 1; flappy_W(2, 193) <= 1; flappy_W(2, 194) <= 1; flappy_W(2, 195) <= 1; flappy_W(2, 196) <= 1; flappy_W(2, 197) <= 1; flappy_W(2, 198) <= 0; flappy_W(2, 199) <= 0; flappy_W(2, 200) <= 0; flappy_W(2, 201) <= 0; flappy_W(2, 202) <= 0; flappy_W(2, 203) <= 0; flappy_W(2, 204) <= 0; flappy_W(2, 205) <= 0; flappy_W(2, 206) <= 0; flappy_W(2, 207) <= 0; flappy_W(2, 208) <= 0; flappy_W(2, 209) <= 0; flappy_W(2, 210) <= 0; flappy_W(2, 211) <= 0; flappy_W(2, 212) <= 0; flappy_W(2, 213) <= 0; flappy_W(2, 214) <= 0; flappy_W(2, 215) <= 0; flappy_W(2, 216) <= 1; flappy_W(2, 217) <= 1; flappy_W(2, 218) <= 1; flappy_W(2, 219) <= 1; flappy_W(2, 220) <= 1; flappy_W(2, 221) <= 1; flappy_W(2, 222) <= 1; flappy_W(2, 223) <= 1; flappy_W(2, 224) <= 1; flappy_W(2, 225) <= 1; flappy_W(2, 226) <= 1; flappy_W(2, 227) <= 1; flappy_W(2, 228) <= 1; flappy_W(2, 229) <= 1; flappy_W(2, 230) <= 1; flappy_W(2, 231) <= 1; flappy_W(2, 232) <= 1; flappy_W(2, 233) <= 1; flappy_W(2, 234) <= 1; flappy_W(2, 235) <= 1; flappy_W(2, 236) <= 1; flappy_W(2, 237) <= 1; flappy_W(2, 238) <= 1; flappy_W(2, 239) <= 1; flappy_W(2, 240) <= 1; flappy_W(2, 241) <= 1; flappy_W(2, 242) <= 1; flappy_W(2, 243) <= 1; flappy_W(2, 244) <= 1; flappy_W(2, 245) <= 1; flappy_W(2, 246) <= 1; flappy_W(2, 247) <= 1; flappy_W(2, 248) <= 1; flappy_W(2, 249) <= 1; flappy_W(2, 250) <= 1; flappy_W(2, 251) <= 1; flappy_W(2, 252) <= 0; flappy_W(2, 253) <= 0; flappy_W(2, 254) <= 0; flappy_W(2, 255) <= 0; flappy_W(2, 256) <= 0; flappy_W(2, 257) <= 0; flappy_W(2, 258) <= 0; flappy_W(2, 259) <= 0; flappy_W(2, 260) <= 0; flappy_W(2, 261) <= 0; flappy_W(2, 262) <= 0; flappy_W(2, 263) <= 0; flappy_W(2, 264) <= 0; flappy_W(2, 265) <= 0; flappy_W(2, 266) <= 0; flappy_W(2, 267) <= 0; flappy_W(2, 268) <= 0; flappy_W(2, 269) <= 0; flappy_W(2, 270) <= 1; flappy_W(2, 271) <= 1; flappy_W(2, 272) <= 1; flappy_W(2, 273) <= 1; flappy_W(2, 274) <= 1; flappy_W(2, 275) <= 1; flappy_W(2, 276) <= 1; flappy_W(2, 277) <= 1; flappy_W(2, 278) <= 1; flappy_W(2, 279) <= 1; flappy_W(2, 280) <= 1; flappy_W(2, 281) <= 1; flappy_W(2, 282) <= 0; flappy_W(2, 283) <= 0; flappy_W(2, 284) <= 0; flappy_W(2, 285) <= 0; flappy_W(2, 286) <= 0; flappy_W(2, 287) <= 0; flappy_W(2, 288) <= 0; flappy_W(2, 289) <= 0; flappy_W(2, 290) <= 0; flappy_W(2, 291) <= 0; flappy_W(2, 292) <= 0; flappy_W(2, 293) <= 0; flappy_W(2, 294) <= 0; flappy_W(2, 295) <= 0; flappy_W(2, 296) <= 0; flappy_W(2, 297) <= 0; flappy_W(2, 298) <= 0; flappy_W(2, 299) <= 0; flappy_W(2, 300) <= 0; flappy_W(2, 301) <= 0; flappy_W(2, 302) <= 0; flappy_W(2, 303) <= 0; flappy_W(2, 304) <= 0; flappy_W(2, 305) <= 0; flappy_W(2, 306) <= 1; flappy_W(2, 307) <= 1; flappy_W(2, 308) <= 1; flappy_W(2, 309) <= 1; flappy_W(2, 310) <= 1; flappy_W(2, 311) <= 1; flappy_W(2, 312) <= 1; flappy_W(2, 313) <= 1; flappy_W(2, 314) <= 1; flappy_W(2, 315) <= 1; flappy_W(2, 316) <= 1; flappy_W(2, 317) <= 1; flappy_W(2, 318) <= 0; flappy_W(2, 319) <= 0; flappy_W(2, 320) <= 0; flappy_W(2, 321) <= 0; flappy_W(2, 322) <= 0; flappy_W(2, 323) <= 0; flappy_W(2, 324) <= 0; flappy_W(2, 325) <= 0; flappy_W(2, 326) <= 0; flappy_W(2, 327) <= 0; flappy_W(2, 328) <= 0; flappy_W(2, 329) <= 0; flappy_W(2, 330) <= 0; flappy_W(2, 331) <= 0; flappy_W(2, 332) <= 0; flappy_W(2, 333) <= 0; flappy_W(2, 334) <= 0; flappy_W(2, 335) <= 0; flappy_W(2, 336) <= 0; flappy_W(2, 337) <= 0; flappy_W(2, 338) <= 0; flappy_W(2, 339) <= 0; flappy_W(2, 340) <= 0; flappy_W(2, 341) <= 0; flappy_W(2, 342) <= 0; flappy_W(2, 343) <= 0; flappy_W(2, 344) <= 0; flappy_W(2, 345) <= 0; flappy_W(2, 346) <= 0; flappy_W(2, 347) <= 0; flappy_W(2, 348) <= 0; flappy_W(2, 349) <= 0; flappy_W(2, 350) <= 0; flappy_W(2, 351) <= 0; flappy_W(2, 352) <= 0; flappy_W(2, 353) <= 0; flappy_W(2, 354) <= 0; flappy_W(2, 355) <= 0; flappy_W(2, 356) <= 0; flappy_W(2, 357) <= 0; flappy_W(2, 358) <= 0; flappy_W(2, 359) <= 0; flappy_W(2, 360) <= 0; flappy_W(2, 361) <= 0; flappy_W(2, 362) <= 0; flappy_W(2, 363) <= 0; flappy_W(2, 364) <= 0; flappy_W(2, 365) <= 0; flappy_W(2, 366) <= 0; flappy_W(2, 367) <= 0; flappy_W(2, 368) <= 0; flappy_W(2, 369) <= 0; flappy_W(2, 370) <= 0; flappy_W(2, 371) <= 0; flappy_W(2, 372) <= 0; flappy_W(2, 373) <= 0; flappy_W(2, 374) <= 0; flappy_W(2, 375) <= 0; flappy_W(2, 376) <= 0; flappy_W(2, 377) <= 0; flappy_W(2, 378) <= 0; flappy_W(2, 379) <= 0; flappy_W(2, 380) <= 0; flappy_W(2, 381) <= 0; flappy_W(2, 382) <= 0; flappy_W(2, 383) <= 0; flappy_W(2, 384) <= 0; flappy_W(2, 385) <= 0; flappy_W(2, 386) <= 0; flappy_W(2, 387) <= 0; flappy_W(2, 388) <= 0; flappy_W(2, 389) <= 0; flappy_W(2, 390) <= 0; flappy_W(2, 391) <= 0; flappy_W(2, 392) <= 0; flappy_W(2, 393) <= 0; flappy_W(2, 394) <= 0; flappy_W(2, 395) <= 0; flappy_W(2, 396) <= 1; flappy_W(2, 397) <= 1; flappy_W(2, 398) <= 1; flappy_W(2, 399) <= 1; flappy_W(2, 400) <= 1; flappy_W(2, 401) <= 1; flappy_W(2, 402) <= 1; flappy_W(2, 403) <= 1; flappy_W(2, 404) <= 1; flappy_W(2, 405) <= 1; flappy_W(2, 406) <= 1; flappy_W(2, 407) <= 1; flappy_W(2, 408) <= 1; flappy_W(2, 409) <= 1; flappy_W(2, 410) <= 1; flappy_W(2, 411) <= 1; flappy_W(2, 412) <= 1; flappy_W(2, 413) <= 1; flappy_W(2, 414) <= 1; flappy_W(2, 415) <= 1; flappy_W(2, 416) <= 1; flappy_W(2, 417) <= 1; flappy_W(2, 418) <= 1; flappy_W(2, 419) <= 1; flappy_W(2, 420) <= 1; flappy_W(2, 421) <= 1; flappy_W(2, 422) <= 1; flappy_W(2, 423) <= 1; flappy_W(2, 424) <= 1; flappy_W(2, 425) <= 1; flappy_W(2, 426) <= 1; flappy_W(2, 427) <= 1; flappy_W(2, 428) <= 1; flappy_W(2, 429) <= 1; flappy_W(2, 430) <= 1; flappy_W(2, 431) <= 1; flappy_W(2, 432) <= 0; flappy_W(2, 433) <= 0; flappy_W(2, 434) <= 0; flappy_W(2, 435) <= 0; flappy_W(2, 436) <= 0; flappy_W(2, 437) <= 0; flappy_W(2, 438) <= 0; flappy_W(2, 439) <= 0; flappy_W(2, 440) <= 0; flappy_W(2, 441) <= 0; flappy_W(2, 442) <= 0; flappy_W(2, 443) <= 0; flappy_W(2, 444) <= 0; flappy_W(2, 445) <= 0; flappy_W(2, 446) <= 0; flappy_W(2, 447) <= 0; flappy_W(2, 448) <= 0; flappy_W(2, 449) <= 0; flappy_W(2, 450) <= 0; flappy_W(2, 451) <= 0; flappy_W(2, 452) <= 0; flappy_W(2, 453) <= 0; flappy_W(2, 454) <= 0; flappy_W(2, 455) <= 0; flappy_W(2, 456) <= 0; flappy_W(2, 457) <= 0; flappy_W(2, 458) <= 0; flappy_W(2, 459) <= 0; flappy_W(2, 460) <= 0; flappy_W(2, 461) <= 0; flappy_W(2, 462) <= 1; flappy_W(2, 463) <= 1; flappy_W(2, 464) <= 1; flappy_W(2, 465) <= 1; flappy_W(2, 466) <= 1; flappy_W(2, 467) <= 1; flappy_W(2, 468) <= 1; flappy_W(2, 469) <= 1; flappy_W(2, 470) <= 1; flappy_W(2, 471) <= 1; flappy_W(2, 472) <= 1; flappy_W(2, 473) <= 1; flappy_W(2, 474) <= 1; flappy_W(2, 475) <= 1; flappy_W(2, 476) <= 1; flappy_W(2, 477) <= 1; flappy_W(2, 478) <= 1; flappy_W(2, 479) <= 1; flappy_W(2, 480) <= 1; flappy_W(2, 481) <= 1; flappy_W(2, 482) <= 1; flappy_W(2, 483) <= 1; flappy_W(2, 484) <= 1; flappy_W(2, 485) <= 1; flappy_W(2, 486) <= 0; flappy_W(2, 487) <= 0; flappy_W(2, 488) <= 0; flappy_W(2, 489) <= 0; flappy_W(2, 490) <= 0; flappy_W(2, 491) <= 0; flappy_W(2, 492) <= 0; flappy_W(2, 493) <= 0; flappy_W(2, 494) <= 0; flappy_W(2, 495) <= 0; flappy_W(2, 496) <= 0; flappy_W(2, 497) <= 0; flappy_W(2, 498) <= 0; flappy_W(2, 499) <= 0; flappy_W(2, 500) <= 0; flappy_W(2, 501) <= 0; flappy_W(2, 502) <= 0; flappy_W(2, 503) <= 0; flappy_W(2, 504) <= 1; flappy_W(2, 505) <= 1; flappy_W(2, 506) <= 1; flappy_W(2, 507) <= 1; flappy_W(2, 508) <= 1; flappy_W(2, 509) <= 1; flappy_W(2, 510) <= 1; flappy_W(2, 511) <= 1; flappy_W(2, 512) <= 1; flappy_W(2, 513) <= 1; flappy_W(2, 514) <= 1; flappy_W(2, 515) <= 1; flappy_W(2, 516) <= 1; flappy_W(2, 517) <= 1; flappy_W(2, 518) <= 1; flappy_W(2, 519) <= 1; flappy_W(2, 520) <= 1; flappy_W(2, 521) <= 1; flappy_W(2, 522) <= 1; flappy_W(2, 523) <= 1; flappy_W(2, 524) <= 1; flappy_W(2, 525) <= 1; flappy_W(2, 526) <= 1; flappy_W(2, 527) <= 1; flappy_W(2, 528) <= 1; flappy_W(2, 529) <= 1; flappy_W(2, 530) <= 1; flappy_W(2, 531) <= 1; flappy_W(2, 532) <= 1; flappy_W(2, 533) <= 1; flappy_W(2, 534) <= 1; flappy_W(2, 535) <= 1; flappy_W(2, 536) <= 1; flappy_W(2, 537) <= 1; flappy_W(2, 538) <= 1; flappy_W(2, 539) <= 1; flappy_W(2, 540) <= 0; flappy_W(2, 541) <= 0; flappy_W(2, 542) <= 0; flappy_W(2, 543) <= 0; flappy_W(2, 544) <= 0; flappy_W(2, 545) <= 0; flappy_W(2, 546) <= 0; flappy_W(2, 547) <= 0; flappy_W(2, 548) <= 0; flappy_W(2, 549) <= 0; flappy_W(2, 550) <= 0; flappy_W(2, 551) <= 0; flappy_W(2, 552) <= 0; flappy_W(2, 553) <= 0; flappy_W(2, 554) <= 0; flappy_W(2, 555) <= 0; flappy_W(2, 556) <= 0; flappy_W(2, 557) <= 0; flappy_W(2, 558) <= 1; flappy_W(2, 559) <= 1; flappy_W(2, 560) <= 1; flappy_W(2, 561) <= 1; flappy_W(2, 562) <= 1; flappy_W(2, 563) <= 1; flappy_W(2, 564) <= 1; flappy_W(2, 565) <= 1; flappy_W(2, 566) <= 1; flappy_W(2, 567) <= 1; flappy_W(2, 568) <= 1; flappy_W(2, 569) <= 1; flappy_W(2, 570) <= 1; flappy_W(2, 571) <= 1; flappy_W(2, 572) <= 1; flappy_W(2, 573) <= 1; flappy_W(2, 574) <= 1; flappy_W(2, 575) <= 1; flappy_W(2, 576) <= 1; flappy_W(2, 577) <= 1; flappy_W(2, 578) <= 1; flappy_W(2, 579) <= 1; flappy_W(2, 580) <= 1; flappy_W(2, 581) <= 1; flappy_W(2, 582) <= 1; flappy_W(2, 583) <= 1; flappy_W(2, 584) <= 1; flappy_W(2, 585) <= 1; flappy_W(2, 586) <= 1; flappy_W(2, 587) <= 1; flappy_W(2, 588) <= 0; flappy_W(2, 589) <= 0; flappy_W(2, 590) <= 0; flappy_W(2, 591) <= 0; flappy_W(2, 592) <= 0; flappy_W(2, 593) <= 0; 
flappy_W(3, 0) <= 1; flappy_W(3, 1) <= 1; flappy_W(3, 2) <= 1; flappy_W(3, 3) <= 1; flappy_W(3, 4) <= 1; flappy_W(3, 5) <= 1; flappy_W(3, 6) <= 1; flappy_W(3, 7) <= 1; flappy_W(3, 8) <= 1; flappy_W(3, 9) <= 1; flappy_W(3, 10) <= 1; flappy_W(3, 11) <= 1; flappy_W(3, 12) <= 1; flappy_W(3, 13) <= 1; flappy_W(3, 14) <= 1; flappy_W(3, 15) <= 1; flappy_W(3, 16) <= 1; flappy_W(3, 17) <= 1; flappy_W(3, 18) <= 1; flappy_W(3, 19) <= 1; flappy_W(3, 20) <= 1; flappy_W(3, 21) <= 1; flappy_W(3, 22) <= 1; flappy_W(3, 23) <= 1; flappy_W(3, 24) <= 1; flappy_W(3, 25) <= 1; flappy_W(3, 26) <= 1; flappy_W(3, 27) <= 1; flappy_W(3, 28) <= 1; flappy_W(3, 29) <= 1; flappy_W(3, 30) <= 1; flappy_W(3, 31) <= 1; flappy_W(3, 32) <= 1; flappy_W(3, 33) <= 1; flappy_W(3, 34) <= 1; flappy_W(3, 35) <= 1; flappy_W(3, 36) <= 1; flappy_W(3, 37) <= 1; flappy_W(3, 38) <= 1; flappy_W(3, 39) <= 1; flappy_W(3, 40) <= 1; flappy_W(3, 41) <= 1; flappy_W(3, 42) <= 0; flappy_W(3, 43) <= 0; flappy_W(3, 44) <= 0; flappy_W(3, 45) <= 0; flappy_W(3, 46) <= 0; flappy_W(3, 47) <= 0; flappy_W(3, 48) <= 0; flappy_W(3, 49) <= 0; flappy_W(3, 50) <= 0; flappy_W(3, 51) <= 0; flappy_W(3, 52) <= 0; flappy_W(3, 53) <= 0; flappy_W(3, 54) <= 1; flappy_W(3, 55) <= 1; flappy_W(3, 56) <= 1; flappy_W(3, 57) <= 1; flappy_W(3, 58) <= 1; flappy_W(3, 59) <= 1; flappy_W(3, 60) <= 1; flappy_W(3, 61) <= 1; flappy_W(3, 62) <= 1; flappy_W(3, 63) <= 1; flappy_W(3, 64) <= 1; flappy_W(3, 65) <= 1; flappy_W(3, 66) <= 1; flappy_W(3, 67) <= 1; flappy_W(3, 68) <= 1; flappy_W(3, 69) <= 1; flappy_W(3, 70) <= 1; flappy_W(3, 71) <= 1; flappy_W(3, 72) <= 1; flappy_W(3, 73) <= 1; flappy_W(3, 74) <= 1; flappy_W(3, 75) <= 1; flappy_W(3, 76) <= 1; flappy_W(3, 77) <= 1; flappy_W(3, 78) <= 0; flappy_W(3, 79) <= 0; flappy_W(3, 80) <= 0; flappy_W(3, 81) <= 0; flappy_W(3, 82) <= 0; flappy_W(3, 83) <= 0; flappy_W(3, 84) <= 0; flappy_W(3, 85) <= 0; flappy_W(3, 86) <= 0; flappy_W(3, 87) <= 0; flappy_W(3, 88) <= 0; flappy_W(3, 89) <= 0; flappy_W(3, 90) <= 0; flappy_W(3, 91) <= 0; flappy_W(3, 92) <= 0; flappy_W(3, 93) <= 0; flappy_W(3, 94) <= 0; flappy_W(3, 95) <= 0; flappy_W(3, 96) <= 0; flappy_W(3, 97) <= 0; flappy_W(3, 98) <= 0; flappy_W(3, 99) <= 0; flappy_W(3, 100) <= 0; flappy_W(3, 101) <= 0; flappy_W(3, 102) <= 0; flappy_W(3, 103) <= 0; flappy_W(3, 104) <= 0; flappy_W(3, 105) <= 0; flappy_W(3, 106) <= 0; flappy_W(3, 107) <= 0; flappy_W(3, 108) <= 0; flappy_W(3, 109) <= 0; flappy_W(3, 110) <= 0; flappy_W(3, 111) <= 0; flappy_W(3, 112) <= 0; flappy_W(3, 113) <= 0; flappy_W(3, 114) <= 0; flappy_W(3, 115) <= 0; flappy_W(3, 116) <= 0; flappy_W(3, 117) <= 0; flappy_W(3, 118) <= 0; flappy_W(3, 119) <= 0; flappy_W(3, 120) <= 0; flappy_W(3, 121) <= 0; flappy_W(3, 122) <= 0; flappy_W(3, 123) <= 0; flappy_W(3, 124) <= 0; flappy_W(3, 125) <= 0; flappy_W(3, 126) <= 1; flappy_W(3, 127) <= 1; flappy_W(3, 128) <= 1; flappy_W(3, 129) <= 1; flappy_W(3, 130) <= 1; flappy_W(3, 131) <= 1; flappy_W(3, 132) <= 0; flappy_W(3, 133) <= 0; flappy_W(3, 134) <= 0; flappy_W(3, 135) <= 0; flappy_W(3, 136) <= 0; flappy_W(3, 137) <= 0; flappy_W(3, 138) <= 0; flappy_W(3, 139) <= 0; flappy_W(3, 140) <= 0; flappy_W(3, 141) <= 0; flappy_W(3, 142) <= 0; flappy_W(3, 143) <= 0; flappy_W(3, 144) <= 0; flappy_W(3, 145) <= 0; flappy_W(3, 146) <= 0; flappy_W(3, 147) <= 0; flappy_W(3, 148) <= 0; flappy_W(3, 149) <= 0; flappy_W(3, 150) <= 0; flappy_W(3, 151) <= 0; flappy_W(3, 152) <= 0; flappy_W(3, 153) <= 0; flappy_W(3, 154) <= 0; flappy_W(3, 155) <= 0; flappy_W(3, 156) <= 0; flappy_W(3, 157) <= 0; flappy_W(3, 158) <= 0; flappy_W(3, 159) <= 0; flappy_W(3, 160) <= 0; flappy_W(3, 161) <= 0; flappy_W(3, 162) <= 1; flappy_W(3, 163) <= 1; flappy_W(3, 164) <= 1; flappy_W(3, 165) <= 1; flappy_W(3, 166) <= 1; flappy_W(3, 167) <= 1; flappy_W(3, 168) <= 1; flappy_W(3, 169) <= 1; flappy_W(3, 170) <= 1; flappy_W(3, 171) <= 1; flappy_W(3, 172) <= 1; flappy_W(3, 173) <= 1; flappy_W(3, 174) <= 1; flappy_W(3, 175) <= 1; flappy_W(3, 176) <= 1; flappy_W(3, 177) <= 1; flappy_W(3, 178) <= 1; flappy_W(3, 179) <= 1; flappy_W(3, 180) <= 1; flappy_W(3, 181) <= 1; flappy_W(3, 182) <= 1; flappy_W(3, 183) <= 1; flappy_W(3, 184) <= 1; flappy_W(3, 185) <= 1; flappy_W(3, 186) <= 1; flappy_W(3, 187) <= 1; flappy_W(3, 188) <= 1; flappy_W(3, 189) <= 1; flappy_W(3, 190) <= 1; flappy_W(3, 191) <= 1; flappy_W(3, 192) <= 1; flappy_W(3, 193) <= 1; flappy_W(3, 194) <= 1; flappy_W(3, 195) <= 1; flappy_W(3, 196) <= 1; flappy_W(3, 197) <= 1; flappy_W(3, 198) <= 0; flappy_W(3, 199) <= 0; flappy_W(3, 200) <= 0; flappy_W(3, 201) <= 0; flappy_W(3, 202) <= 0; flappy_W(3, 203) <= 0; flappy_W(3, 204) <= 0; flappy_W(3, 205) <= 0; flappy_W(3, 206) <= 0; flappy_W(3, 207) <= 0; flappy_W(3, 208) <= 0; flappy_W(3, 209) <= 0; flappy_W(3, 210) <= 0; flappy_W(3, 211) <= 0; flappy_W(3, 212) <= 0; flappy_W(3, 213) <= 0; flappy_W(3, 214) <= 0; flappy_W(3, 215) <= 0; flappy_W(3, 216) <= 1; flappy_W(3, 217) <= 1; flappy_W(3, 218) <= 1; flappy_W(3, 219) <= 1; flappy_W(3, 220) <= 1; flappy_W(3, 221) <= 1; flappy_W(3, 222) <= 1; flappy_W(3, 223) <= 1; flappy_W(3, 224) <= 1; flappy_W(3, 225) <= 1; flappy_W(3, 226) <= 1; flappy_W(3, 227) <= 1; flappy_W(3, 228) <= 1; flappy_W(3, 229) <= 1; flappy_W(3, 230) <= 1; flappy_W(3, 231) <= 1; flappy_W(3, 232) <= 1; flappy_W(3, 233) <= 1; flappy_W(3, 234) <= 1; flappy_W(3, 235) <= 1; flappy_W(3, 236) <= 1; flappy_W(3, 237) <= 1; flappy_W(3, 238) <= 1; flappy_W(3, 239) <= 1; flappy_W(3, 240) <= 1; flappy_W(3, 241) <= 1; flappy_W(3, 242) <= 1; flappy_W(3, 243) <= 1; flappy_W(3, 244) <= 1; flappy_W(3, 245) <= 1; flappy_W(3, 246) <= 1; flappy_W(3, 247) <= 1; flappy_W(3, 248) <= 1; flappy_W(3, 249) <= 1; flappy_W(3, 250) <= 1; flappy_W(3, 251) <= 1; flappy_W(3, 252) <= 0; flappy_W(3, 253) <= 0; flappy_W(3, 254) <= 0; flappy_W(3, 255) <= 0; flappy_W(3, 256) <= 0; flappy_W(3, 257) <= 0; flappy_W(3, 258) <= 0; flappy_W(3, 259) <= 0; flappy_W(3, 260) <= 0; flappy_W(3, 261) <= 0; flappy_W(3, 262) <= 0; flappy_W(3, 263) <= 0; flappy_W(3, 264) <= 0; flappy_W(3, 265) <= 0; flappy_W(3, 266) <= 0; flappy_W(3, 267) <= 0; flappy_W(3, 268) <= 0; flappy_W(3, 269) <= 0; flappy_W(3, 270) <= 1; flappy_W(3, 271) <= 1; flappy_W(3, 272) <= 1; flappy_W(3, 273) <= 1; flappy_W(3, 274) <= 1; flappy_W(3, 275) <= 1; flappy_W(3, 276) <= 1; flappy_W(3, 277) <= 1; flappy_W(3, 278) <= 1; flappy_W(3, 279) <= 1; flappy_W(3, 280) <= 1; flappy_W(3, 281) <= 1; flappy_W(3, 282) <= 0; flappy_W(3, 283) <= 0; flappy_W(3, 284) <= 0; flappy_W(3, 285) <= 0; flappy_W(3, 286) <= 0; flappy_W(3, 287) <= 0; flappy_W(3, 288) <= 0; flappy_W(3, 289) <= 0; flappy_W(3, 290) <= 0; flappy_W(3, 291) <= 0; flappy_W(3, 292) <= 0; flappy_W(3, 293) <= 0; flappy_W(3, 294) <= 0; flappy_W(3, 295) <= 0; flappy_W(3, 296) <= 0; flappy_W(3, 297) <= 0; flappy_W(3, 298) <= 0; flappy_W(3, 299) <= 0; flappy_W(3, 300) <= 0; flappy_W(3, 301) <= 0; flappy_W(3, 302) <= 0; flappy_W(3, 303) <= 0; flappy_W(3, 304) <= 0; flappy_W(3, 305) <= 0; flappy_W(3, 306) <= 1; flappy_W(3, 307) <= 1; flappy_W(3, 308) <= 1; flappy_W(3, 309) <= 1; flappy_W(3, 310) <= 1; flappy_W(3, 311) <= 1; flappy_W(3, 312) <= 1; flappy_W(3, 313) <= 1; flappy_W(3, 314) <= 1; flappy_W(3, 315) <= 1; flappy_W(3, 316) <= 1; flappy_W(3, 317) <= 1; flappy_W(3, 318) <= 0; flappy_W(3, 319) <= 0; flappy_W(3, 320) <= 0; flappy_W(3, 321) <= 0; flappy_W(3, 322) <= 0; flappy_W(3, 323) <= 0; flappy_W(3, 324) <= 0; flappy_W(3, 325) <= 0; flappy_W(3, 326) <= 0; flappy_W(3, 327) <= 0; flappy_W(3, 328) <= 0; flappy_W(3, 329) <= 0; flappy_W(3, 330) <= 0; flappy_W(3, 331) <= 0; flappy_W(3, 332) <= 0; flappy_W(3, 333) <= 0; flappy_W(3, 334) <= 0; flappy_W(3, 335) <= 0; flappy_W(3, 336) <= 0; flappy_W(3, 337) <= 0; flappy_W(3, 338) <= 0; flappy_W(3, 339) <= 0; flappy_W(3, 340) <= 0; flappy_W(3, 341) <= 0; flappy_W(3, 342) <= 0; flappy_W(3, 343) <= 0; flappy_W(3, 344) <= 0; flappy_W(3, 345) <= 0; flappy_W(3, 346) <= 0; flappy_W(3, 347) <= 0; flappy_W(3, 348) <= 0; flappy_W(3, 349) <= 0; flappy_W(3, 350) <= 0; flappy_W(3, 351) <= 0; flappy_W(3, 352) <= 0; flappy_W(3, 353) <= 0; flappy_W(3, 354) <= 0; flappy_W(3, 355) <= 0; flappy_W(3, 356) <= 0; flappy_W(3, 357) <= 0; flappy_W(3, 358) <= 0; flappy_W(3, 359) <= 0; flappy_W(3, 360) <= 0; flappy_W(3, 361) <= 0; flappy_W(3, 362) <= 0; flappy_W(3, 363) <= 0; flappy_W(3, 364) <= 0; flappy_W(3, 365) <= 0; flappy_W(3, 366) <= 0; flappy_W(3, 367) <= 0; flappy_W(3, 368) <= 0; flappy_W(3, 369) <= 0; flappy_W(3, 370) <= 0; flappy_W(3, 371) <= 0; flappy_W(3, 372) <= 0; flappy_W(3, 373) <= 0; flappy_W(3, 374) <= 0; flappy_W(3, 375) <= 0; flappy_W(3, 376) <= 0; flappy_W(3, 377) <= 0; flappy_W(3, 378) <= 0; flappy_W(3, 379) <= 0; flappy_W(3, 380) <= 0; flappy_W(3, 381) <= 0; flappy_W(3, 382) <= 0; flappy_W(3, 383) <= 0; flappy_W(3, 384) <= 0; flappy_W(3, 385) <= 0; flappy_W(3, 386) <= 0; flappy_W(3, 387) <= 0; flappy_W(3, 388) <= 0; flappy_W(3, 389) <= 0; flappy_W(3, 390) <= 0; flappy_W(3, 391) <= 0; flappy_W(3, 392) <= 0; flappy_W(3, 393) <= 0; flappy_W(3, 394) <= 0; flappy_W(3, 395) <= 0; flappy_W(3, 396) <= 1; flappy_W(3, 397) <= 1; flappy_W(3, 398) <= 1; flappy_W(3, 399) <= 1; flappy_W(3, 400) <= 1; flappy_W(3, 401) <= 1; flappy_W(3, 402) <= 1; flappy_W(3, 403) <= 1; flappy_W(3, 404) <= 1; flappy_W(3, 405) <= 1; flappy_W(3, 406) <= 1; flappy_W(3, 407) <= 1; flappy_W(3, 408) <= 1; flappy_W(3, 409) <= 1; flappy_W(3, 410) <= 1; flappy_W(3, 411) <= 1; flappy_W(3, 412) <= 1; flappy_W(3, 413) <= 1; flappy_W(3, 414) <= 1; flappy_W(3, 415) <= 1; flappy_W(3, 416) <= 1; flappy_W(3, 417) <= 1; flappy_W(3, 418) <= 1; flappy_W(3, 419) <= 1; flappy_W(3, 420) <= 1; flappy_W(3, 421) <= 1; flappy_W(3, 422) <= 1; flappy_W(3, 423) <= 1; flappy_W(3, 424) <= 1; flappy_W(3, 425) <= 1; flappy_W(3, 426) <= 1; flappy_W(3, 427) <= 1; flappy_W(3, 428) <= 1; flappy_W(3, 429) <= 1; flappy_W(3, 430) <= 1; flappy_W(3, 431) <= 1; flappy_W(3, 432) <= 0; flappy_W(3, 433) <= 0; flappy_W(3, 434) <= 0; flappy_W(3, 435) <= 0; flappy_W(3, 436) <= 0; flappy_W(3, 437) <= 0; flappy_W(3, 438) <= 0; flappy_W(3, 439) <= 0; flappy_W(3, 440) <= 0; flappy_W(3, 441) <= 0; flappy_W(3, 442) <= 0; flappy_W(3, 443) <= 0; flappy_W(3, 444) <= 0; flappy_W(3, 445) <= 0; flappy_W(3, 446) <= 0; flappy_W(3, 447) <= 0; flappy_W(3, 448) <= 0; flappy_W(3, 449) <= 0; flappy_W(3, 450) <= 0; flappy_W(3, 451) <= 0; flappy_W(3, 452) <= 0; flappy_W(3, 453) <= 0; flappy_W(3, 454) <= 0; flappy_W(3, 455) <= 0; flappy_W(3, 456) <= 0; flappy_W(3, 457) <= 0; flappy_W(3, 458) <= 0; flappy_W(3, 459) <= 0; flappy_W(3, 460) <= 0; flappy_W(3, 461) <= 0; flappy_W(3, 462) <= 1; flappy_W(3, 463) <= 1; flappy_W(3, 464) <= 1; flappy_W(3, 465) <= 1; flappy_W(3, 466) <= 1; flappy_W(3, 467) <= 1; flappy_W(3, 468) <= 1; flappy_W(3, 469) <= 1; flappy_W(3, 470) <= 1; flappy_W(3, 471) <= 1; flappy_W(3, 472) <= 1; flappy_W(3, 473) <= 1; flappy_W(3, 474) <= 1; flappy_W(3, 475) <= 1; flappy_W(3, 476) <= 1; flappy_W(3, 477) <= 1; flappy_W(3, 478) <= 1; flappy_W(3, 479) <= 1; flappy_W(3, 480) <= 1; flappy_W(3, 481) <= 1; flappy_W(3, 482) <= 1; flappy_W(3, 483) <= 1; flappy_W(3, 484) <= 1; flappy_W(3, 485) <= 1; flappy_W(3, 486) <= 0; flappy_W(3, 487) <= 0; flappy_W(3, 488) <= 0; flappy_W(3, 489) <= 0; flappy_W(3, 490) <= 0; flappy_W(3, 491) <= 0; flappy_W(3, 492) <= 0; flappy_W(3, 493) <= 0; flappy_W(3, 494) <= 0; flappy_W(3, 495) <= 0; flappy_W(3, 496) <= 0; flappy_W(3, 497) <= 0; flappy_W(3, 498) <= 0; flappy_W(3, 499) <= 0; flappy_W(3, 500) <= 0; flappy_W(3, 501) <= 0; flappy_W(3, 502) <= 0; flappy_W(3, 503) <= 0; flappy_W(3, 504) <= 1; flappy_W(3, 505) <= 1; flappy_W(3, 506) <= 1; flappy_W(3, 507) <= 1; flappy_W(3, 508) <= 1; flappy_W(3, 509) <= 1; flappy_W(3, 510) <= 1; flappy_W(3, 511) <= 1; flappy_W(3, 512) <= 1; flappy_W(3, 513) <= 1; flappy_W(3, 514) <= 1; flappy_W(3, 515) <= 1; flappy_W(3, 516) <= 1; flappy_W(3, 517) <= 1; flappy_W(3, 518) <= 1; flappy_W(3, 519) <= 1; flappy_W(3, 520) <= 1; flappy_W(3, 521) <= 1; flappy_W(3, 522) <= 1; flappy_W(3, 523) <= 1; flappy_W(3, 524) <= 1; flappy_W(3, 525) <= 1; flappy_W(3, 526) <= 1; flappy_W(3, 527) <= 1; flappy_W(3, 528) <= 1; flappy_W(3, 529) <= 1; flappy_W(3, 530) <= 1; flappy_W(3, 531) <= 1; flappy_W(3, 532) <= 1; flappy_W(3, 533) <= 1; flappy_W(3, 534) <= 1; flappy_W(3, 535) <= 1; flappy_W(3, 536) <= 1; flappy_W(3, 537) <= 1; flappy_W(3, 538) <= 1; flappy_W(3, 539) <= 1; flappy_W(3, 540) <= 0; flappy_W(3, 541) <= 0; flappy_W(3, 542) <= 0; flappy_W(3, 543) <= 0; flappy_W(3, 544) <= 0; flappy_W(3, 545) <= 0; flappy_W(3, 546) <= 0; flappy_W(3, 547) <= 0; flappy_W(3, 548) <= 0; flappy_W(3, 549) <= 0; flappy_W(3, 550) <= 0; flappy_W(3, 551) <= 0; flappy_W(3, 552) <= 0; flappy_W(3, 553) <= 0; flappy_W(3, 554) <= 0; flappy_W(3, 555) <= 0; flappy_W(3, 556) <= 0; flappy_W(3, 557) <= 0; flappy_W(3, 558) <= 1; flappy_W(3, 559) <= 1; flappy_W(3, 560) <= 1; flappy_W(3, 561) <= 1; flappy_W(3, 562) <= 1; flappy_W(3, 563) <= 1; flappy_W(3, 564) <= 1; flappy_W(3, 565) <= 1; flappy_W(3, 566) <= 1; flappy_W(3, 567) <= 1; flappy_W(3, 568) <= 1; flappy_W(3, 569) <= 1; flappy_W(3, 570) <= 1; flappy_W(3, 571) <= 1; flappy_W(3, 572) <= 1; flappy_W(3, 573) <= 1; flappy_W(3, 574) <= 1; flappy_W(3, 575) <= 1; flappy_W(3, 576) <= 1; flappy_W(3, 577) <= 1; flappy_W(3, 578) <= 1; flappy_W(3, 579) <= 1; flappy_W(3, 580) <= 1; flappy_W(3, 581) <= 1; flappy_W(3, 582) <= 1; flappy_W(3, 583) <= 1; flappy_W(3, 584) <= 1; flappy_W(3, 585) <= 1; flappy_W(3, 586) <= 1; flappy_W(3, 587) <= 1; flappy_W(3, 588) <= 0; flappy_W(3, 589) <= 0; flappy_W(3, 590) <= 0; flappy_W(3, 591) <= 0; flappy_W(3, 592) <= 0; flappy_W(3, 593) <= 0; 
flappy_W(4, 0) <= 1; flappy_W(4, 1) <= 1; flappy_W(4, 2) <= 1; flappy_W(4, 3) <= 1; flappy_W(4, 4) <= 1; flappy_W(4, 5) <= 1; flappy_W(4, 6) <= 1; flappy_W(4, 7) <= 1; flappy_W(4, 8) <= 1; flappy_W(4, 9) <= 1; flappy_W(4, 10) <= 1; flappy_W(4, 11) <= 1; flappy_W(4, 12) <= 1; flappy_W(4, 13) <= 1; flappy_W(4, 14) <= 1; flappy_W(4, 15) <= 1; flappy_W(4, 16) <= 1; flappy_W(4, 17) <= 1; flappy_W(4, 18) <= 1; flappy_W(4, 19) <= 1; flappy_W(4, 20) <= 1; flappy_W(4, 21) <= 1; flappy_W(4, 22) <= 1; flappy_W(4, 23) <= 1; flappy_W(4, 24) <= 1; flappy_W(4, 25) <= 1; flappy_W(4, 26) <= 1; flappy_W(4, 27) <= 1; flappy_W(4, 28) <= 1; flappy_W(4, 29) <= 1; flappy_W(4, 30) <= 1; flappy_W(4, 31) <= 1; flappy_W(4, 32) <= 1; flappy_W(4, 33) <= 1; flappy_W(4, 34) <= 1; flappy_W(4, 35) <= 1; flappy_W(4, 36) <= 1; flappy_W(4, 37) <= 1; flappy_W(4, 38) <= 1; flappy_W(4, 39) <= 1; flappy_W(4, 40) <= 1; flappy_W(4, 41) <= 1; flappy_W(4, 42) <= 0; flappy_W(4, 43) <= 0; flappy_W(4, 44) <= 0; flappy_W(4, 45) <= 0; flappy_W(4, 46) <= 0; flappy_W(4, 47) <= 0; flappy_W(4, 48) <= 0; flappy_W(4, 49) <= 0; flappy_W(4, 50) <= 0; flappy_W(4, 51) <= 0; flappy_W(4, 52) <= 0; flappy_W(4, 53) <= 0; flappy_W(4, 54) <= 1; flappy_W(4, 55) <= 1; flappy_W(4, 56) <= 1; flappy_W(4, 57) <= 1; flappy_W(4, 58) <= 1; flappy_W(4, 59) <= 1; flappy_W(4, 60) <= 1; flappy_W(4, 61) <= 1; flappy_W(4, 62) <= 1; flappy_W(4, 63) <= 1; flappy_W(4, 64) <= 1; flappy_W(4, 65) <= 1; flappy_W(4, 66) <= 1; flappy_W(4, 67) <= 1; flappy_W(4, 68) <= 1; flappy_W(4, 69) <= 1; flappy_W(4, 70) <= 1; flappy_W(4, 71) <= 1; flappy_W(4, 72) <= 1; flappy_W(4, 73) <= 1; flappy_W(4, 74) <= 1; flappy_W(4, 75) <= 1; flappy_W(4, 76) <= 1; flappy_W(4, 77) <= 1; flappy_W(4, 78) <= 0; flappy_W(4, 79) <= 0; flappy_W(4, 80) <= 0; flappy_W(4, 81) <= 0; flappy_W(4, 82) <= 0; flappy_W(4, 83) <= 0; flappy_W(4, 84) <= 0; flappy_W(4, 85) <= 0; flappy_W(4, 86) <= 0; flappy_W(4, 87) <= 0; flappy_W(4, 88) <= 0; flappy_W(4, 89) <= 0; flappy_W(4, 90) <= 0; flappy_W(4, 91) <= 0; flappy_W(4, 92) <= 0; flappy_W(4, 93) <= 0; flappy_W(4, 94) <= 0; flappy_W(4, 95) <= 0; flappy_W(4, 96) <= 0; flappy_W(4, 97) <= 0; flappy_W(4, 98) <= 0; flappy_W(4, 99) <= 0; flappy_W(4, 100) <= 0; flappy_W(4, 101) <= 0; flappy_W(4, 102) <= 0; flappy_W(4, 103) <= 0; flappy_W(4, 104) <= 0; flappy_W(4, 105) <= 0; flappy_W(4, 106) <= 0; flappy_W(4, 107) <= 0; flappy_W(4, 108) <= 0; flappy_W(4, 109) <= 0; flappy_W(4, 110) <= 0; flappy_W(4, 111) <= 0; flappy_W(4, 112) <= 0; flappy_W(4, 113) <= 0; flappy_W(4, 114) <= 0; flappy_W(4, 115) <= 0; flappy_W(4, 116) <= 0; flappy_W(4, 117) <= 0; flappy_W(4, 118) <= 0; flappy_W(4, 119) <= 0; flappy_W(4, 120) <= 0; flappy_W(4, 121) <= 0; flappy_W(4, 122) <= 0; flappy_W(4, 123) <= 0; flappy_W(4, 124) <= 0; flappy_W(4, 125) <= 0; flappy_W(4, 126) <= 1; flappy_W(4, 127) <= 1; flappy_W(4, 128) <= 1; flappy_W(4, 129) <= 1; flappy_W(4, 130) <= 1; flappy_W(4, 131) <= 1; flappy_W(4, 132) <= 0; flappy_W(4, 133) <= 0; flappy_W(4, 134) <= 0; flappy_W(4, 135) <= 0; flappy_W(4, 136) <= 0; flappy_W(4, 137) <= 0; flappy_W(4, 138) <= 0; flappy_W(4, 139) <= 0; flappy_W(4, 140) <= 0; flappy_W(4, 141) <= 0; flappy_W(4, 142) <= 0; flappy_W(4, 143) <= 0; flappy_W(4, 144) <= 0; flappy_W(4, 145) <= 0; flappy_W(4, 146) <= 0; flappy_W(4, 147) <= 0; flappy_W(4, 148) <= 0; flappy_W(4, 149) <= 0; flappy_W(4, 150) <= 0; flappy_W(4, 151) <= 0; flappy_W(4, 152) <= 0; flappy_W(4, 153) <= 0; flappy_W(4, 154) <= 0; flappy_W(4, 155) <= 0; flappy_W(4, 156) <= 0; flappy_W(4, 157) <= 0; flappy_W(4, 158) <= 0; flappy_W(4, 159) <= 0; flappy_W(4, 160) <= 0; flappy_W(4, 161) <= 0; flappy_W(4, 162) <= 1; flappy_W(4, 163) <= 1; flappy_W(4, 164) <= 1; flappy_W(4, 165) <= 1; flappy_W(4, 166) <= 1; flappy_W(4, 167) <= 1; flappy_W(4, 168) <= 1; flappy_W(4, 169) <= 1; flappy_W(4, 170) <= 1; flappy_W(4, 171) <= 1; flappy_W(4, 172) <= 1; flappy_W(4, 173) <= 1; flappy_W(4, 174) <= 1; flappy_W(4, 175) <= 1; flappy_W(4, 176) <= 1; flappy_W(4, 177) <= 1; flappy_W(4, 178) <= 1; flappy_W(4, 179) <= 1; flappy_W(4, 180) <= 1; flappy_W(4, 181) <= 1; flappy_W(4, 182) <= 1; flappy_W(4, 183) <= 1; flappy_W(4, 184) <= 1; flappy_W(4, 185) <= 1; flappy_W(4, 186) <= 1; flappy_W(4, 187) <= 1; flappy_W(4, 188) <= 1; flappy_W(4, 189) <= 1; flappy_W(4, 190) <= 1; flappy_W(4, 191) <= 1; flappy_W(4, 192) <= 1; flappy_W(4, 193) <= 1; flappy_W(4, 194) <= 1; flappy_W(4, 195) <= 1; flappy_W(4, 196) <= 1; flappy_W(4, 197) <= 1; flappy_W(4, 198) <= 0; flappy_W(4, 199) <= 0; flappy_W(4, 200) <= 0; flappy_W(4, 201) <= 0; flappy_W(4, 202) <= 0; flappy_W(4, 203) <= 0; flappy_W(4, 204) <= 0; flappy_W(4, 205) <= 0; flappy_W(4, 206) <= 0; flappy_W(4, 207) <= 0; flappy_W(4, 208) <= 0; flappy_W(4, 209) <= 0; flappy_W(4, 210) <= 0; flappy_W(4, 211) <= 0; flappy_W(4, 212) <= 0; flappy_W(4, 213) <= 0; flappy_W(4, 214) <= 0; flappy_W(4, 215) <= 0; flappy_W(4, 216) <= 1; flappy_W(4, 217) <= 1; flappy_W(4, 218) <= 1; flappy_W(4, 219) <= 1; flappy_W(4, 220) <= 1; flappy_W(4, 221) <= 1; flappy_W(4, 222) <= 1; flappy_W(4, 223) <= 1; flappy_W(4, 224) <= 1; flappy_W(4, 225) <= 1; flappy_W(4, 226) <= 1; flappy_W(4, 227) <= 1; flappy_W(4, 228) <= 1; flappy_W(4, 229) <= 1; flappy_W(4, 230) <= 1; flappy_W(4, 231) <= 1; flappy_W(4, 232) <= 1; flappy_W(4, 233) <= 1; flappy_W(4, 234) <= 1; flappy_W(4, 235) <= 1; flappy_W(4, 236) <= 1; flappy_W(4, 237) <= 1; flappy_W(4, 238) <= 1; flappy_W(4, 239) <= 1; flappy_W(4, 240) <= 1; flappy_W(4, 241) <= 1; flappy_W(4, 242) <= 1; flappy_W(4, 243) <= 1; flappy_W(4, 244) <= 1; flappy_W(4, 245) <= 1; flappy_W(4, 246) <= 1; flappy_W(4, 247) <= 1; flappy_W(4, 248) <= 1; flappy_W(4, 249) <= 1; flappy_W(4, 250) <= 1; flappy_W(4, 251) <= 1; flappy_W(4, 252) <= 0; flappy_W(4, 253) <= 0; flappy_W(4, 254) <= 0; flappy_W(4, 255) <= 0; flappy_W(4, 256) <= 0; flappy_W(4, 257) <= 0; flappy_W(4, 258) <= 0; flappy_W(4, 259) <= 0; flappy_W(4, 260) <= 0; flappy_W(4, 261) <= 0; flappy_W(4, 262) <= 0; flappy_W(4, 263) <= 0; flappy_W(4, 264) <= 0; flappy_W(4, 265) <= 0; flappy_W(4, 266) <= 0; flappy_W(4, 267) <= 0; flappy_W(4, 268) <= 0; flappy_W(4, 269) <= 0; flappy_W(4, 270) <= 1; flappy_W(4, 271) <= 1; flappy_W(4, 272) <= 1; flappy_W(4, 273) <= 1; flappy_W(4, 274) <= 1; flappy_W(4, 275) <= 1; flappy_W(4, 276) <= 1; flappy_W(4, 277) <= 1; flappy_W(4, 278) <= 1; flappy_W(4, 279) <= 1; flappy_W(4, 280) <= 1; flappy_W(4, 281) <= 1; flappy_W(4, 282) <= 0; flappy_W(4, 283) <= 0; flappy_W(4, 284) <= 0; flappy_W(4, 285) <= 0; flappy_W(4, 286) <= 0; flappy_W(4, 287) <= 0; flappy_W(4, 288) <= 0; flappy_W(4, 289) <= 0; flappy_W(4, 290) <= 0; flappy_W(4, 291) <= 0; flappy_W(4, 292) <= 0; flappy_W(4, 293) <= 0; flappy_W(4, 294) <= 0; flappy_W(4, 295) <= 0; flappy_W(4, 296) <= 0; flappy_W(4, 297) <= 0; flappy_W(4, 298) <= 0; flappy_W(4, 299) <= 0; flappy_W(4, 300) <= 0; flappy_W(4, 301) <= 0; flappy_W(4, 302) <= 0; flappy_W(4, 303) <= 0; flappy_W(4, 304) <= 0; flappy_W(4, 305) <= 0; flappy_W(4, 306) <= 1; flappy_W(4, 307) <= 1; flappy_W(4, 308) <= 1; flappy_W(4, 309) <= 1; flappy_W(4, 310) <= 1; flappy_W(4, 311) <= 1; flappy_W(4, 312) <= 1; flappy_W(4, 313) <= 1; flappy_W(4, 314) <= 1; flappy_W(4, 315) <= 1; flappy_W(4, 316) <= 1; flappy_W(4, 317) <= 1; flappy_W(4, 318) <= 0; flappy_W(4, 319) <= 0; flappy_W(4, 320) <= 0; flappy_W(4, 321) <= 0; flappy_W(4, 322) <= 0; flappy_W(4, 323) <= 0; flappy_W(4, 324) <= 0; flappy_W(4, 325) <= 0; flappy_W(4, 326) <= 0; flappy_W(4, 327) <= 0; flappy_W(4, 328) <= 0; flappy_W(4, 329) <= 0; flappy_W(4, 330) <= 0; flappy_W(4, 331) <= 0; flappy_W(4, 332) <= 0; flappy_W(4, 333) <= 0; flappy_W(4, 334) <= 0; flappy_W(4, 335) <= 0; flappy_W(4, 336) <= 0; flappy_W(4, 337) <= 0; flappy_W(4, 338) <= 0; flappy_W(4, 339) <= 0; flappy_W(4, 340) <= 0; flappy_W(4, 341) <= 0; flappy_W(4, 342) <= 0; flappy_W(4, 343) <= 0; flappy_W(4, 344) <= 0; flappy_W(4, 345) <= 0; flappy_W(4, 346) <= 0; flappy_W(4, 347) <= 0; flappy_W(4, 348) <= 0; flappy_W(4, 349) <= 0; flappy_W(4, 350) <= 0; flappy_W(4, 351) <= 0; flappy_W(4, 352) <= 0; flappy_W(4, 353) <= 0; flappy_W(4, 354) <= 0; flappy_W(4, 355) <= 0; flappy_W(4, 356) <= 0; flappy_W(4, 357) <= 0; flappy_W(4, 358) <= 0; flappy_W(4, 359) <= 0; flappy_W(4, 360) <= 0; flappy_W(4, 361) <= 0; flappy_W(4, 362) <= 0; flappy_W(4, 363) <= 0; flappy_W(4, 364) <= 0; flappy_W(4, 365) <= 0; flappy_W(4, 366) <= 0; flappy_W(4, 367) <= 0; flappy_W(4, 368) <= 0; flappy_W(4, 369) <= 0; flappy_W(4, 370) <= 0; flappy_W(4, 371) <= 0; flappy_W(4, 372) <= 0; flappy_W(4, 373) <= 0; flappy_W(4, 374) <= 0; flappy_W(4, 375) <= 0; flappy_W(4, 376) <= 0; flappy_W(4, 377) <= 0; flappy_W(4, 378) <= 0; flappy_W(4, 379) <= 0; flappy_W(4, 380) <= 0; flappy_W(4, 381) <= 0; flappy_W(4, 382) <= 0; flappy_W(4, 383) <= 0; flappy_W(4, 384) <= 0; flappy_W(4, 385) <= 0; flappy_W(4, 386) <= 0; flappy_W(4, 387) <= 0; flappy_W(4, 388) <= 0; flappy_W(4, 389) <= 0; flappy_W(4, 390) <= 0; flappy_W(4, 391) <= 0; flappy_W(4, 392) <= 0; flappy_W(4, 393) <= 0; flappy_W(4, 394) <= 0; flappy_W(4, 395) <= 0; flappy_W(4, 396) <= 1; flappy_W(4, 397) <= 1; flappy_W(4, 398) <= 1; flappy_W(4, 399) <= 1; flappy_W(4, 400) <= 1; flappy_W(4, 401) <= 1; flappy_W(4, 402) <= 1; flappy_W(4, 403) <= 1; flappy_W(4, 404) <= 1; flappy_W(4, 405) <= 1; flappy_W(4, 406) <= 1; flappy_W(4, 407) <= 1; flappy_W(4, 408) <= 1; flappy_W(4, 409) <= 1; flappy_W(4, 410) <= 1; flappy_W(4, 411) <= 1; flappy_W(4, 412) <= 1; flappy_W(4, 413) <= 1; flappy_W(4, 414) <= 1; flappy_W(4, 415) <= 1; flappy_W(4, 416) <= 1; flappy_W(4, 417) <= 1; flappy_W(4, 418) <= 1; flappy_W(4, 419) <= 1; flappy_W(4, 420) <= 1; flappy_W(4, 421) <= 1; flappy_W(4, 422) <= 1; flappy_W(4, 423) <= 1; flappy_W(4, 424) <= 1; flappy_W(4, 425) <= 1; flappy_W(4, 426) <= 1; flappy_W(4, 427) <= 1; flappy_W(4, 428) <= 1; flappy_W(4, 429) <= 1; flappy_W(4, 430) <= 1; flappy_W(4, 431) <= 1; flappy_W(4, 432) <= 0; flappy_W(4, 433) <= 0; flappy_W(4, 434) <= 0; flappy_W(4, 435) <= 0; flappy_W(4, 436) <= 0; flappy_W(4, 437) <= 0; flappy_W(4, 438) <= 0; flappy_W(4, 439) <= 0; flappy_W(4, 440) <= 0; flappy_W(4, 441) <= 0; flappy_W(4, 442) <= 0; flappy_W(4, 443) <= 0; flappy_W(4, 444) <= 0; flappy_W(4, 445) <= 0; flappy_W(4, 446) <= 0; flappy_W(4, 447) <= 0; flappy_W(4, 448) <= 0; flappy_W(4, 449) <= 0; flappy_W(4, 450) <= 0; flappy_W(4, 451) <= 0; flappy_W(4, 452) <= 0; flappy_W(4, 453) <= 0; flappy_W(4, 454) <= 0; flappy_W(4, 455) <= 0; flappy_W(4, 456) <= 0; flappy_W(4, 457) <= 0; flappy_W(4, 458) <= 0; flappy_W(4, 459) <= 0; flappy_W(4, 460) <= 0; flappy_W(4, 461) <= 0; flappy_W(4, 462) <= 1; flappy_W(4, 463) <= 1; flappy_W(4, 464) <= 1; flappy_W(4, 465) <= 1; flappy_W(4, 466) <= 1; flappy_W(4, 467) <= 1; flappy_W(4, 468) <= 1; flappy_W(4, 469) <= 1; flappy_W(4, 470) <= 1; flappy_W(4, 471) <= 1; flappy_W(4, 472) <= 1; flappy_W(4, 473) <= 1; flappy_W(4, 474) <= 1; flappy_W(4, 475) <= 1; flappy_W(4, 476) <= 1; flappy_W(4, 477) <= 1; flappy_W(4, 478) <= 1; flappy_W(4, 479) <= 1; flappy_W(4, 480) <= 1; flappy_W(4, 481) <= 1; flappy_W(4, 482) <= 1; flappy_W(4, 483) <= 1; flappy_W(4, 484) <= 1; flappy_W(4, 485) <= 1; flappy_W(4, 486) <= 0; flappy_W(4, 487) <= 0; flappy_W(4, 488) <= 0; flappy_W(4, 489) <= 0; flappy_W(4, 490) <= 0; flappy_W(4, 491) <= 0; flappy_W(4, 492) <= 0; flappy_W(4, 493) <= 0; flappy_W(4, 494) <= 0; flappy_W(4, 495) <= 0; flappy_W(4, 496) <= 0; flappy_W(4, 497) <= 0; flappy_W(4, 498) <= 0; flappy_W(4, 499) <= 0; flappy_W(4, 500) <= 0; flappy_W(4, 501) <= 0; flappy_W(4, 502) <= 0; flappy_W(4, 503) <= 0; flappy_W(4, 504) <= 1; flappy_W(4, 505) <= 1; flappy_W(4, 506) <= 1; flappy_W(4, 507) <= 1; flappy_W(4, 508) <= 1; flappy_W(4, 509) <= 1; flappy_W(4, 510) <= 1; flappy_W(4, 511) <= 1; flappy_W(4, 512) <= 1; flappy_W(4, 513) <= 1; flappy_W(4, 514) <= 1; flappy_W(4, 515) <= 1; flappy_W(4, 516) <= 1; flappy_W(4, 517) <= 1; flappy_W(4, 518) <= 1; flappy_W(4, 519) <= 1; flappy_W(4, 520) <= 1; flappy_W(4, 521) <= 1; flappy_W(4, 522) <= 1; flappy_W(4, 523) <= 1; flappy_W(4, 524) <= 1; flappy_W(4, 525) <= 1; flappy_W(4, 526) <= 1; flappy_W(4, 527) <= 1; flappy_W(4, 528) <= 1; flappy_W(4, 529) <= 1; flappy_W(4, 530) <= 1; flappy_W(4, 531) <= 1; flappy_W(4, 532) <= 1; flappy_W(4, 533) <= 1; flappy_W(4, 534) <= 1; flappy_W(4, 535) <= 1; flappy_W(4, 536) <= 1; flappy_W(4, 537) <= 1; flappy_W(4, 538) <= 1; flappy_W(4, 539) <= 1; flappy_W(4, 540) <= 0; flappy_W(4, 541) <= 0; flappy_W(4, 542) <= 0; flappy_W(4, 543) <= 0; flappy_W(4, 544) <= 0; flappy_W(4, 545) <= 0; flappy_W(4, 546) <= 0; flappy_W(4, 547) <= 0; flappy_W(4, 548) <= 0; flappy_W(4, 549) <= 0; flappy_W(4, 550) <= 0; flappy_W(4, 551) <= 0; flappy_W(4, 552) <= 0; flappy_W(4, 553) <= 0; flappy_W(4, 554) <= 0; flappy_W(4, 555) <= 0; flappy_W(4, 556) <= 0; flappy_W(4, 557) <= 0; flappy_W(4, 558) <= 1; flappy_W(4, 559) <= 1; flappy_W(4, 560) <= 1; flappy_W(4, 561) <= 1; flappy_W(4, 562) <= 1; flappy_W(4, 563) <= 1; flappy_W(4, 564) <= 1; flappy_W(4, 565) <= 1; flappy_W(4, 566) <= 1; flappy_W(4, 567) <= 1; flappy_W(4, 568) <= 1; flappy_W(4, 569) <= 1; flappy_W(4, 570) <= 1; flappy_W(4, 571) <= 1; flappy_W(4, 572) <= 1; flappy_W(4, 573) <= 1; flappy_W(4, 574) <= 1; flappy_W(4, 575) <= 1; flappy_W(4, 576) <= 1; flappy_W(4, 577) <= 1; flappy_W(4, 578) <= 1; flappy_W(4, 579) <= 1; flappy_W(4, 580) <= 1; flappy_W(4, 581) <= 1; flappy_W(4, 582) <= 1; flappy_W(4, 583) <= 1; flappy_W(4, 584) <= 1; flappy_W(4, 585) <= 1; flappy_W(4, 586) <= 1; flappy_W(4, 587) <= 1; flappy_W(4, 588) <= 0; flappy_W(4, 589) <= 0; flappy_W(4, 590) <= 0; flappy_W(4, 591) <= 0; flappy_W(4, 592) <= 0; flappy_W(4, 593) <= 0; 
flappy_W(5, 0) <= 1; flappy_W(5, 1) <= 1; flappy_W(5, 2) <= 1; flappy_W(5, 3) <= 1; flappy_W(5, 4) <= 1; flappy_W(5, 5) <= 1; flappy_W(5, 6) <= 1; flappy_W(5, 7) <= 1; flappy_W(5, 8) <= 1; flappy_W(5, 9) <= 1; flappy_W(5, 10) <= 1; flappy_W(5, 11) <= 1; flappy_W(5, 12) <= 1; flappy_W(5, 13) <= 1; flappy_W(5, 14) <= 1; flappy_W(5, 15) <= 1; flappy_W(5, 16) <= 1; flappy_W(5, 17) <= 1; flappy_W(5, 18) <= 1; flappy_W(5, 19) <= 1; flappy_W(5, 20) <= 1; flappy_W(5, 21) <= 1; flappy_W(5, 22) <= 1; flappy_W(5, 23) <= 1; flappy_W(5, 24) <= 1; flappy_W(5, 25) <= 1; flappy_W(5, 26) <= 1; flappy_W(5, 27) <= 1; flappy_W(5, 28) <= 1; flappy_W(5, 29) <= 1; flappy_W(5, 30) <= 1; flappy_W(5, 31) <= 1; flappy_W(5, 32) <= 1; flappy_W(5, 33) <= 1; flappy_W(5, 34) <= 1; flappy_W(5, 35) <= 1; flappy_W(5, 36) <= 1; flappy_W(5, 37) <= 1; flappy_W(5, 38) <= 1; flappy_W(5, 39) <= 1; flappy_W(5, 40) <= 1; flappy_W(5, 41) <= 1; flappy_W(5, 42) <= 0; flappy_W(5, 43) <= 0; flappy_W(5, 44) <= 0; flappy_W(5, 45) <= 0; flappy_W(5, 46) <= 0; flappy_W(5, 47) <= 0; flappy_W(5, 48) <= 0; flappy_W(5, 49) <= 0; flappy_W(5, 50) <= 0; flappy_W(5, 51) <= 0; flappy_W(5, 52) <= 0; flappy_W(5, 53) <= 0; flappy_W(5, 54) <= 1; flappy_W(5, 55) <= 1; flappy_W(5, 56) <= 1; flappy_W(5, 57) <= 1; flappy_W(5, 58) <= 1; flappy_W(5, 59) <= 1; flappy_W(5, 60) <= 1; flappy_W(5, 61) <= 1; flappy_W(5, 62) <= 1; flappy_W(5, 63) <= 1; flappy_W(5, 64) <= 1; flappy_W(5, 65) <= 1; flappy_W(5, 66) <= 1; flappy_W(5, 67) <= 1; flappy_W(5, 68) <= 1; flappy_W(5, 69) <= 1; flappy_W(5, 70) <= 1; flappy_W(5, 71) <= 1; flappy_W(5, 72) <= 1; flappy_W(5, 73) <= 1; flappy_W(5, 74) <= 1; flappy_W(5, 75) <= 1; flappy_W(5, 76) <= 1; flappy_W(5, 77) <= 1; flappy_W(5, 78) <= 0; flappy_W(5, 79) <= 0; flappy_W(5, 80) <= 0; flappy_W(5, 81) <= 0; flappy_W(5, 82) <= 0; flappy_W(5, 83) <= 0; flappy_W(5, 84) <= 0; flappy_W(5, 85) <= 0; flappy_W(5, 86) <= 0; flappy_W(5, 87) <= 0; flappy_W(5, 88) <= 0; flappy_W(5, 89) <= 0; flappy_W(5, 90) <= 0; flappy_W(5, 91) <= 0; flappy_W(5, 92) <= 0; flappy_W(5, 93) <= 0; flappy_W(5, 94) <= 0; flappy_W(5, 95) <= 0; flappy_W(5, 96) <= 0; flappy_W(5, 97) <= 0; flappy_W(5, 98) <= 0; flappy_W(5, 99) <= 0; flappy_W(5, 100) <= 0; flappy_W(5, 101) <= 0; flappy_W(5, 102) <= 0; flappy_W(5, 103) <= 0; flappy_W(5, 104) <= 0; flappy_W(5, 105) <= 0; flappy_W(5, 106) <= 0; flappy_W(5, 107) <= 0; flappy_W(5, 108) <= 0; flappy_W(5, 109) <= 0; flappy_W(5, 110) <= 0; flappy_W(5, 111) <= 0; flappy_W(5, 112) <= 0; flappy_W(5, 113) <= 0; flappy_W(5, 114) <= 0; flappy_W(5, 115) <= 0; flappy_W(5, 116) <= 0; flappy_W(5, 117) <= 0; flappy_W(5, 118) <= 0; flappy_W(5, 119) <= 0; flappy_W(5, 120) <= 0; flappy_W(5, 121) <= 0; flappy_W(5, 122) <= 0; flappy_W(5, 123) <= 0; flappy_W(5, 124) <= 0; flappy_W(5, 125) <= 0; flappy_W(5, 126) <= 1; flappy_W(5, 127) <= 1; flappy_W(5, 128) <= 1; flappy_W(5, 129) <= 1; flappy_W(5, 130) <= 1; flappy_W(5, 131) <= 1; flappy_W(5, 132) <= 0; flappy_W(5, 133) <= 0; flappy_W(5, 134) <= 0; flappy_W(5, 135) <= 0; flappy_W(5, 136) <= 0; flappy_W(5, 137) <= 0; flappy_W(5, 138) <= 0; flappy_W(5, 139) <= 0; flappy_W(5, 140) <= 0; flappy_W(5, 141) <= 0; flappy_W(5, 142) <= 0; flappy_W(5, 143) <= 0; flappy_W(5, 144) <= 0; flappy_W(5, 145) <= 0; flappy_W(5, 146) <= 0; flappy_W(5, 147) <= 0; flappy_W(5, 148) <= 0; flappy_W(5, 149) <= 0; flappy_W(5, 150) <= 0; flappy_W(5, 151) <= 0; flappy_W(5, 152) <= 0; flappy_W(5, 153) <= 0; flappy_W(5, 154) <= 0; flappy_W(5, 155) <= 0; flappy_W(5, 156) <= 0; flappy_W(5, 157) <= 0; flappy_W(5, 158) <= 0; flappy_W(5, 159) <= 0; flappy_W(5, 160) <= 0; flappy_W(5, 161) <= 0; flappy_W(5, 162) <= 1; flappy_W(5, 163) <= 1; flappy_W(5, 164) <= 1; flappy_W(5, 165) <= 1; flappy_W(5, 166) <= 1; flappy_W(5, 167) <= 1; flappy_W(5, 168) <= 1; flappy_W(5, 169) <= 1; flappy_W(5, 170) <= 1; flappy_W(5, 171) <= 1; flappy_W(5, 172) <= 1; flappy_W(5, 173) <= 1; flappy_W(5, 174) <= 1; flappy_W(5, 175) <= 1; flappy_W(5, 176) <= 1; flappy_W(5, 177) <= 1; flappy_W(5, 178) <= 1; flappy_W(5, 179) <= 1; flappy_W(5, 180) <= 1; flappy_W(5, 181) <= 1; flappy_W(5, 182) <= 1; flappy_W(5, 183) <= 1; flappy_W(5, 184) <= 1; flappy_W(5, 185) <= 1; flappy_W(5, 186) <= 1; flappy_W(5, 187) <= 1; flappy_W(5, 188) <= 1; flappy_W(5, 189) <= 1; flappy_W(5, 190) <= 1; flappy_W(5, 191) <= 1; flappy_W(5, 192) <= 1; flappy_W(5, 193) <= 1; flappy_W(5, 194) <= 1; flappy_W(5, 195) <= 1; flappy_W(5, 196) <= 1; flappy_W(5, 197) <= 1; flappy_W(5, 198) <= 0; flappy_W(5, 199) <= 0; flappy_W(5, 200) <= 0; flappy_W(5, 201) <= 0; flappy_W(5, 202) <= 0; flappy_W(5, 203) <= 0; flappy_W(5, 204) <= 0; flappy_W(5, 205) <= 0; flappy_W(5, 206) <= 0; flappy_W(5, 207) <= 0; flappy_W(5, 208) <= 0; flappy_W(5, 209) <= 0; flappy_W(5, 210) <= 0; flappy_W(5, 211) <= 0; flappy_W(5, 212) <= 0; flappy_W(5, 213) <= 0; flappy_W(5, 214) <= 0; flappy_W(5, 215) <= 0; flappy_W(5, 216) <= 1; flappy_W(5, 217) <= 1; flappy_W(5, 218) <= 1; flappy_W(5, 219) <= 1; flappy_W(5, 220) <= 1; flappy_W(5, 221) <= 1; flappy_W(5, 222) <= 1; flappy_W(5, 223) <= 1; flappy_W(5, 224) <= 1; flappy_W(5, 225) <= 1; flappy_W(5, 226) <= 1; flappy_W(5, 227) <= 1; flappy_W(5, 228) <= 1; flappy_W(5, 229) <= 1; flappy_W(5, 230) <= 1; flappy_W(5, 231) <= 1; flappy_W(5, 232) <= 1; flappy_W(5, 233) <= 1; flappy_W(5, 234) <= 1; flappy_W(5, 235) <= 1; flappy_W(5, 236) <= 1; flappy_W(5, 237) <= 1; flappy_W(5, 238) <= 1; flappy_W(5, 239) <= 1; flappy_W(5, 240) <= 1; flappy_W(5, 241) <= 1; flappy_W(5, 242) <= 1; flappy_W(5, 243) <= 1; flappy_W(5, 244) <= 1; flappy_W(5, 245) <= 1; flappy_W(5, 246) <= 1; flappy_W(5, 247) <= 1; flappy_W(5, 248) <= 1; flappy_W(5, 249) <= 1; flappy_W(5, 250) <= 1; flappy_W(5, 251) <= 1; flappy_W(5, 252) <= 0; flappy_W(5, 253) <= 0; flappy_W(5, 254) <= 0; flappy_W(5, 255) <= 0; flappy_W(5, 256) <= 0; flappy_W(5, 257) <= 0; flappy_W(5, 258) <= 0; flappy_W(5, 259) <= 0; flappy_W(5, 260) <= 0; flappy_W(5, 261) <= 0; flappy_W(5, 262) <= 0; flappy_W(5, 263) <= 0; flappy_W(5, 264) <= 0; flappy_W(5, 265) <= 0; flappy_W(5, 266) <= 0; flappy_W(5, 267) <= 0; flappy_W(5, 268) <= 0; flappy_W(5, 269) <= 0; flappy_W(5, 270) <= 1; flappy_W(5, 271) <= 1; flappy_W(5, 272) <= 1; flappy_W(5, 273) <= 1; flappy_W(5, 274) <= 1; flappy_W(5, 275) <= 1; flappy_W(5, 276) <= 1; flappy_W(5, 277) <= 1; flappy_W(5, 278) <= 1; flappy_W(5, 279) <= 1; flappy_W(5, 280) <= 1; flappy_W(5, 281) <= 1; flappy_W(5, 282) <= 0; flappy_W(5, 283) <= 0; flappy_W(5, 284) <= 0; flappy_W(5, 285) <= 0; flappy_W(5, 286) <= 0; flappy_W(5, 287) <= 0; flappy_W(5, 288) <= 0; flappy_W(5, 289) <= 0; flappy_W(5, 290) <= 0; flappy_W(5, 291) <= 0; flappy_W(5, 292) <= 0; flappy_W(5, 293) <= 0; flappy_W(5, 294) <= 0; flappy_W(5, 295) <= 0; flappy_W(5, 296) <= 0; flappy_W(5, 297) <= 0; flappy_W(5, 298) <= 0; flappy_W(5, 299) <= 0; flappy_W(5, 300) <= 0; flappy_W(5, 301) <= 0; flappy_W(5, 302) <= 0; flappy_W(5, 303) <= 0; flappy_W(5, 304) <= 0; flappy_W(5, 305) <= 0; flappy_W(5, 306) <= 1; flappy_W(5, 307) <= 1; flappy_W(5, 308) <= 1; flappy_W(5, 309) <= 1; flappy_W(5, 310) <= 1; flappy_W(5, 311) <= 1; flappy_W(5, 312) <= 1; flappy_W(5, 313) <= 1; flappy_W(5, 314) <= 1; flappy_W(5, 315) <= 1; flappy_W(5, 316) <= 1; flappy_W(5, 317) <= 1; flappy_W(5, 318) <= 0; flappy_W(5, 319) <= 0; flappy_W(5, 320) <= 0; flappy_W(5, 321) <= 0; flappy_W(5, 322) <= 0; flappy_W(5, 323) <= 0; flappy_W(5, 324) <= 0; flappy_W(5, 325) <= 0; flappy_W(5, 326) <= 0; flappy_W(5, 327) <= 0; flappy_W(5, 328) <= 0; flappy_W(5, 329) <= 0; flappy_W(5, 330) <= 0; flappy_W(5, 331) <= 0; flappy_W(5, 332) <= 0; flappy_W(5, 333) <= 0; flappy_W(5, 334) <= 0; flappy_W(5, 335) <= 0; flappy_W(5, 336) <= 0; flappy_W(5, 337) <= 0; flappy_W(5, 338) <= 0; flappy_W(5, 339) <= 0; flappy_W(5, 340) <= 0; flappy_W(5, 341) <= 0; flappy_W(5, 342) <= 0; flappy_W(5, 343) <= 0; flappy_W(5, 344) <= 0; flappy_W(5, 345) <= 0; flappy_W(5, 346) <= 0; flappy_W(5, 347) <= 0; flappy_W(5, 348) <= 0; flappy_W(5, 349) <= 0; flappy_W(5, 350) <= 0; flappy_W(5, 351) <= 0; flappy_W(5, 352) <= 0; flappy_W(5, 353) <= 0; flappy_W(5, 354) <= 0; flappy_W(5, 355) <= 0; flappy_W(5, 356) <= 0; flappy_W(5, 357) <= 0; flappy_W(5, 358) <= 0; flappy_W(5, 359) <= 0; flappy_W(5, 360) <= 0; flappy_W(5, 361) <= 0; flappy_W(5, 362) <= 0; flappy_W(5, 363) <= 0; flappy_W(5, 364) <= 0; flappy_W(5, 365) <= 0; flappy_W(5, 366) <= 0; flappy_W(5, 367) <= 0; flappy_W(5, 368) <= 0; flappy_W(5, 369) <= 0; flappy_W(5, 370) <= 0; flappy_W(5, 371) <= 0; flappy_W(5, 372) <= 0; flappy_W(5, 373) <= 0; flappy_W(5, 374) <= 0; flappy_W(5, 375) <= 0; flappy_W(5, 376) <= 0; flappy_W(5, 377) <= 0; flappy_W(5, 378) <= 0; flappy_W(5, 379) <= 0; flappy_W(5, 380) <= 0; flappy_W(5, 381) <= 0; flappy_W(5, 382) <= 0; flappy_W(5, 383) <= 0; flappy_W(5, 384) <= 0; flappy_W(5, 385) <= 0; flappy_W(5, 386) <= 0; flappy_W(5, 387) <= 0; flappy_W(5, 388) <= 0; flappy_W(5, 389) <= 0; flappy_W(5, 390) <= 0; flappy_W(5, 391) <= 0; flappy_W(5, 392) <= 0; flappy_W(5, 393) <= 0; flappy_W(5, 394) <= 0; flappy_W(5, 395) <= 0; flappy_W(5, 396) <= 1; flappy_W(5, 397) <= 1; flappy_W(5, 398) <= 1; flappy_W(5, 399) <= 1; flappy_W(5, 400) <= 1; flappy_W(5, 401) <= 1; flappy_W(5, 402) <= 1; flappy_W(5, 403) <= 1; flappy_W(5, 404) <= 1; flappy_W(5, 405) <= 1; flappy_W(5, 406) <= 1; flappy_W(5, 407) <= 1; flappy_W(5, 408) <= 1; flappy_W(5, 409) <= 1; flappy_W(5, 410) <= 1; flappy_W(5, 411) <= 1; flappy_W(5, 412) <= 1; flappy_W(5, 413) <= 1; flappy_W(5, 414) <= 1; flappy_W(5, 415) <= 1; flappy_W(5, 416) <= 1; flappy_W(5, 417) <= 1; flappy_W(5, 418) <= 1; flappy_W(5, 419) <= 1; flappy_W(5, 420) <= 1; flappy_W(5, 421) <= 1; flappy_W(5, 422) <= 1; flappy_W(5, 423) <= 1; flappy_W(5, 424) <= 1; flappy_W(5, 425) <= 1; flappy_W(5, 426) <= 1; flappy_W(5, 427) <= 1; flappy_W(5, 428) <= 1; flappy_W(5, 429) <= 1; flappy_W(5, 430) <= 1; flappy_W(5, 431) <= 1; flappy_W(5, 432) <= 0; flappy_W(5, 433) <= 0; flappy_W(5, 434) <= 0; flappy_W(5, 435) <= 0; flappy_W(5, 436) <= 0; flappy_W(5, 437) <= 0; flappy_W(5, 438) <= 0; flappy_W(5, 439) <= 0; flappy_W(5, 440) <= 0; flappy_W(5, 441) <= 0; flappy_W(5, 442) <= 0; flappy_W(5, 443) <= 0; flappy_W(5, 444) <= 0; flappy_W(5, 445) <= 0; flappy_W(5, 446) <= 0; flappy_W(5, 447) <= 0; flappy_W(5, 448) <= 0; flappy_W(5, 449) <= 0; flappy_W(5, 450) <= 0; flappy_W(5, 451) <= 0; flappy_W(5, 452) <= 0; flappy_W(5, 453) <= 0; flappy_W(5, 454) <= 0; flappy_W(5, 455) <= 0; flappy_W(5, 456) <= 0; flappy_W(5, 457) <= 0; flappy_W(5, 458) <= 0; flappy_W(5, 459) <= 0; flappy_W(5, 460) <= 0; flappy_W(5, 461) <= 0; flappy_W(5, 462) <= 1; flappy_W(5, 463) <= 1; flappy_W(5, 464) <= 1; flappy_W(5, 465) <= 1; flappy_W(5, 466) <= 1; flappy_W(5, 467) <= 1; flappy_W(5, 468) <= 1; flappy_W(5, 469) <= 1; flappy_W(5, 470) <= 1; flappy_W(5, 471) <= 1; flappy_W(5, 472) <= 1; flappy_W(5, 473) <= 1; flappy_W(5, 474) <= 1; flappy_W(5, 475) <= 1; flappy_W(5, 476) <= 1; flappy_W(5, 477) <= 1; flappy_W(5, 478) <= 1; flappy_W(5, 479) <= 1; flappy_W(5, 480) <= 1; flappy_W(5, 481) <= 1; flappy_W(5, 482) <= 1; flappy_W(5, 483) <= 1; flappy_W(5, 484) <= 1; flappy_W(5, 485) <= 1; flappy_W(5, 486) <= 0; flappy_W(5, 487) <= 0; flappy_W(5, 488) <= 0; flappy_W(5, 489) <= 0; flappy_W(5, 490) <= 0; flappy_W(5, 491) <= 0; flappy_W(5, 492) <= 0; flappy_W(5, 493) <= 0; flappy_W(5, 494) <= 0; flappy_W(5, 495) <= 0; flappy_W(5, 496) <= 0; flappy_W(5, 497) <= 0; flappy_W(5, 498) <= 0; flappy_W(5, 499) <= 0; flappy_W(5, 500) <= 0; flappy_W(5, 501) <= 0; flappy_W(5, 502) <= 0; flappy_W(5, 503) <= 0; flappy_W(5, 504) <= 1; flappy_W(5, 505) <= 1; flappy_W(5, 506) <= 1; flappy_W(5, 507) <= 1; flappy_W(5, 508) <= 1; flappy_W(5, 509) <= 1; flappy_W(5, 510) <= 1; flappy_W(5, 511) <= 1; flappy_W(5, 512) <= 1; flappy_W(5, 513) <= 1; flappy_W(5, 514) <= 1; flappy_W(5, 515) <= 1; flappy_W(5, 516) <= 1; flappy_W(5, 517) <= 1; flappy_W(5, 518) <= 1; flappy_W(5, 519) <= 1; flappy_W(5, 520) <= 1; flappy_W(5, 521) <= 1; flappy_W(5, 522) <= 1; flappy_W(5, 523) <= 1; flappy_W(5, 524) <= 1; flappy_W(5, 525) <= 1; flappy_W(5, 526) <= 1; flappy_W(5, 527) <= 1; flappy_W(5, 528) <= 1; flappy_W(5, 529) <= 1; flappy_W(5, 530) <= 1; flappy_W(5, 531) <= 1; flappy_W(5, 532) <= 1; flappy_W(5, 533) <= 1; flappy_W(5, 534) <= 1; flappy_W(5, 535) <= 1; flappy_W(5, 536) <= 1; flappy_W(5, 537) <= 1; flappy_W(5, 538) <= 1; flappy_W(5, 539) <= 1; flappy_W(5, 540) <= 0; flappy_W(5, 541) <= 0; flappy_W(5, 542) <= 0; flappy_W(5, 543) <= 0; flappy_W(5, 544) <= 0; flappy_W(5, 545) <= 0; flappy_W(5, 546) <= 0; flappy_W(5, 547) <= 0; flappy_W(5, 548) <= 0; flappy_W(5, 549) <= 0; flappy_W(5, 550) <= 0; flappy_W(5, 551) <= 0; flappy_W(5, 552) <= 0; flappy_W(5, 553) <= 0; flappy_W(5, 554) <= 0; flappy_W(5, 555) <= 0; flappy_W(5, 556) <= 0; flappy_W(5, 557) <= 0; flappy_W(5, 558) <= 1; flappy_W(5, 559) <= 1; flappy_W(5, 560) <= 1; flappy_W(5, 561) <= 1; flappy_W(5, 562) <= 1; flappy_W(5, 563) <= 1; flappy_W(5, 564) <= 1; flappy_W(5, 565) <= 1; flappy_W(5, 566) <= 1; flappy_W(5, 567) <= 1; flappy_W(5, 568) <= 1; flappy_W(5, 569) <= 1; flappy_W(5, 570) <= 1; flappy_W(5, 571) <= 1; flappy_W(5, 572) <= 1; flappy_W(5, 573) <= 1; flappy_W(5, 574) <= 1; flappy_W(5, 575) <= 1; flappy_W(5, 576) <= 1; flappy_W(5, 577) <= 1; flappy_W(5, 578) <= 1; flappy_W(5, 579) <= 1; flappy_W(5, 580) <= 1; flappy_W(5, 581) <= 1; flappy_W(5, 582) <= 1; flappy_W(5, 583) <= 1; flappy_W(5, 584) <= 1; flappy_W(5, 585) <= 1; flappy_W(5, 586) <= 1; flappy_W(5, 587) <= 1; flappy_W(5, 588) <= 0; flappy_W(5, 589) <= 0; flappy_W(5, 590) <= 0; flappy_W(5, 591) <= 0; flappy_W(5, 592) <= 0; flappy_W(5, 593) <= 0; 
flappy_W(6, 0) <= 0; flappy_W(6, 1) <= 0; flappy_W(6, 2) <= 0; flappy_W(6, 3) <= 0; flappy_W(6, 4) <= 0; flappy_W(6, 5) <= 0; flappy_W(6, 6) <= 1; flappy_W(6, 7) <= 1; flappy_W(6, 8) <= 1; flappy_W(6, 9) <= 1; flappy_W(6, 10) <= 1; flappy_W(6, 11) <= 1; flappy_W(6, 12) <= 1; flappy_W(6, 13) <= 1; flappy_W(6, 14) <= 1; flappy_W(6, 15) <= 1; flappy_W(6, 16) <= 1; flappy_W(6, 17) <= 1; flappy_W(6, 18) <= 0; flappy_W(6, 19) <= 0; flappy_W(6, 20) <= 0; flappy_W(6, 21) <= 0; flappy_W(6, 22) <= 0; flappy_W(6, 23) <= 0; flappy_W(6, 24) <= 0; flappy_W(6, 25) <= 0; flappy_W(6, 26) <= 0; flappy_W(6, 27) <= 0; flappy_W(6, 28) <= 0; flappy_W(6, 29) <= 0; flappy_W(6, 30) <= 1; flappy_W(6, 31) <= 1; flappy_W(6, 32) <= 1; flappy_W(6, 33) <= 1; flappy_W(6, 34) <= 1; flappy_W(6, 35) <= 1; flappy_W(6, 36) <= 1; flappy_W(6, 37) <= 1; flappy_W(6, 38) <= 1; flappy_W(6, 39) <= 1; flappy_W(6, 40) <= 1; flappy_W(6, 41) <= 1; flappy_W(6, 42) <= 0; flappy_W(6, 43) <= 0; flappy_W(6, 44) <= 0; flappy_W(6, 45) <= 0; flappy_W(6, 46) <= 0; flappy_W(6, 47) <= 0; flappy_W(6, 48) <= 0; flappy_W(6, 49) <= 0; flappy_W(6, 50) <= 0; flappy_W(6, 51) <= 0; flappy_W(6, 52) <= 0; flappy_W(6, 53) <= 0; flappy_W(6, 54) <= 0; flappy_W(6, 55) <= 0; flappy_W(6, 56) <= 0; flappy_W(6, 57) <= 0; flappy_W(6, 58) <= 0; flappy_W(6, 59) <= 0; flappy_W(6, 60) <= 1; flappy_W(6, 61) <= 1; flappy_W(6, 62) <= 1; flappy_W(6, 63) <= 1; flappy_W(6, 64) <= 1; flappy_W(6, 65) <= 1; flappy_W(6, 66) <= 1; flappy_W(6, 67) <= 1; flappy_W(6, 68) <= 1; flappy_W(6, 69) <= 1; flappy_W(6, 70) <= 1; flappy_W(6, 71) <= 1; flappy_W(6, 72) <= 0; flappy_W(6, 73) <= 0; flappy_W(6, 74) <= 0; flappy_W(6, 75) <= 0; flappy_W(6, 76) <= 0; flappy_W(6, 77) <= 0; flappy_W(6, 78) <= 0; flappy_W(6, 79) <= 0; flappy_W(6, 80) <= 0; flappy_W(6, 81) <= 0; flappy_W(6, 82) <= 0; flappy_W(6, 83) <= 0; flappy_W(6, 84) <= 0; flappy_W(6, 85) <= 0; flappy_W(6, 86) <= 0; flappy_W(6, 87) <= 0; flappy_W(6, 88) <= 0; flappy_W(6, 89) <= 0; flappy_W(6, 90) <= 0; flappy_W(6, 91) <= 0; flappy_W(6, 92) <= 0; flappy_W(6, 93) <= 0; flappy_W(6, 94) <= 0; flappy_W(6, 95) <= 0; flappy_W(6, 96) <= 0; flappy_W(6, 97) <= 0; flappy_W(6, 98) <= 0; flappy_W(6, 99) <= 0; flappy_W(6, 100) <= 0; flappy_W(6, 101) <= 0; flappy_W(6, 102) <= 0; flappy_W(6, 103) <= 0; flappy_W(6, 104) <= 0; flappy_W(6, 105) <= 0; flappy_W(6, 106) <= 0; flappy_W(6, 107) <= 0; flappy_W(6, 108) <= 0; flappy_W(6, 109) <= 0; flappy_W(6, 110) <= 0; flappy_W(6, 111) <= 0; flappy_W(6, 112) <= 0; flappy_W(6, 113) <= 0; flappy_W(6, 114) <= 0; flappy_W(6, 115) <= 0; flappy_W(6, 116) <= 0; flappy_W(6, 117) <= 0; flappy_W(6, 118) <= 0; flappy_W(6, 119) <= 0; flappy_W(6, 120) <= 1; flappy_W(6, 121) <= 1; flappy_W(6, 122) <= 1; flappy_W(6, 123) <= 1; flappy_W(6, 124) <= 1; flappy_W(6, 125) <= 1; flappy_W(6, 126) <= 1; flappy_W(6, 127) <= 1; flappy_W(6, 128) <= 1; flappy_W(6, 129) <= 1; flappy_W(6, 130) <= 1; flappy_W(6, 131) <= 1; flappy_W(6, 132) <= 1; flappy_W(6, 133) <= 1; flappy_W(6, 134) <= 1; flappy_W(6, 135) <= 1; flappy_W(6, 136) <= 1; flappy_W(6, 137) <= 1; flappy_W(6, 138) <= 0; flappy_W(6, 139) <= 0; flappy_W(6, 140) <= 0; flappy_W(6, 141) <= 0; flappy_W(6, 142) <= 0; flappy_W(6, 143) <= 0; flappy_W(6, 144) <= 0; flappy_W(6, 145) <= 0; flappy_W(6, 146) <= 0; flappy_W(6, 147) <= 0; flappy_W(6, 148) <= 0; flappy_W(6, 149) <= 0; flappy_W(6, 150) <= 0; flappy_W(6, 151) <= 0; flappy_W(6, 152) <= 0; flappy_W(6, 153) <= 0; flappy_W(6, 154) <= 0; flappy_W(6, 155) <= 0; flappy_W(6, 156) <= 0; flappy_W(6, 157) <= 0; flappy_W(6, 158) <= 0; flappy_W(6, 159) <= 0; flappy_W(6, 160) <= 0; flappy_W(6, 161) <= 0; flappy_W(6, 162) <= 0; flappy_W(6, 163) <= 0; flappy_W(6, 164) <= 0; flappy_W(6, 165) <= 0; flappy_W(6, 166) <= 0; flappy_W(6, 167) <= 0; flappy_W(6, 168) <= 1; flappy_W(6, 169) <= 1; flappy_W(6, 170) <= 1; flappy_W(6, 171) <= 1; flappy_W(6, 172) <= 1; flappy_W(6, 173) <= 1; flappy_W(6, 174) <= 1; flappy_W(6, 175) <= 1; flappy_W(6, 176) <= 1; flappy_W(6, 177) <= 1; flappy_W(6, 178) <= 1; flappy_W(6, 179) <= 1; flappy_W(6, 180) <= 0; flappy_W(6, 181) <= 0; flappy_W(6, 182) <= 0; flappy_W(6, 183) <= 0; flappy_W(6, 184) <= 0; flappy_W(6, 185) <= 0; flappy_W(6, 186) <= 0; flappy_W(6, 187) <= 0; flappy_W(6, 188) <= 0; flappy_W(6, 189) <= 0; flappy_W(6, 190) <= 0; flappy_W(6, 191) <= 0; flappy_W(6, 192) <= 1; flappy_W(6, 193) <= 1; flappy_W(6, 194) <= 1; flappy_W(6, 195) <= 1; flappy_W(6, 196) <= 1; flappy_W(6, 197) <= 1; flappy_W(6, 198) <= 1; flappy_W(6, 199) <= 1; flappy_W(6, 200) <= 1; flappy_W(6, 201) <= 1; flappy_W(6, 202) <= 1; flappy_W(6, 203) <= 1; flappy_W(6, 204) <= 0; flappy_W(6, 205) <= 0; flappy_W(6, 206) <= 0; flappy_W(6, 207) <= 0; flappy_W(6, 208) <= 0; flappy_W(6, 209) <= 0; flappy_W(6, 210) <= 0; flappy_W(6, 211) <= 0; flappy_W(6, 212) <= 0; flappy_W(6, 213) <= 0; flappy_W(6, 214) <= 0; flappy_W(6, 215) <= 0; flappy_W(6, 216) <= 0; flappy_W(6, 217) <= 0; flappy_W(6, 218) <= 0; flappy_W(6, 219) <= 0; flappy_W(6, 220) <= 0; flappy_W(6, 221) <= 0; flappy_W(6, 222) <= 1; flappy_W(6, 223) <= 1; flappy_W(6, 224) <= 1; flappy_W(6, 225) <= 1; flappy_W(6, 226) <= 1; flappy_W(6, 227) <= 1; flappy_W(6, 228) <= 1; flappy_W(6, 229) <= 1; flappy_W(6, 230) <= 1; flappy_W(6, 231) <= 1; flappy_W(6, 232) <= 1; flappy_W(6, 233) <= 1; flappy_W(6, 234) <= 0; flappy_W(6, 235) <= 0; flappy_W(6, 236) <= 0; flappy_W(6, 237) <= 0; flappy_W(6, 238) <= 0; flappy_W(6, 239) <= 0; flappy_W(6, 240) <= 0; flappy_W(6, 241) <= 0; flappy_W(6, 242) <= 0; flappy_W(6, 243) <= 0; flappy_W(6, 244) <= 0; flappy_W(6, 245) <= 0; flappy_W(6, 246) <= 1; flappy_W(6, 247) <= 1; flappy_W(6, 248) <= 1; flappy_W(6, 249) <= 1; flappy_W(6, 250) <= 1; flappy_W(6, 251) <= 1; flappy_W(6, 252) <= 1; flappy_W(6, 253) <= 1; flappy_W(6, 254) <= 1; flappy_W(6, 255) <= 1; flappy_W(6, 256) <= 1; flappy_W(6, 257) <= 1; flappy_W(6, 258) <= 0; flappy_W(6, 259) <= 0; flappy_W(6, 260) <= 0; flappy_W(6, 261) <= 0; flappy_W(6, 262) <= 0; flappy_W(6, 263) <= 0; flappy_W(6, 264) <= 0; flappy_W(6, 265) <= 0; flappy_W(6, 266) <= 0; flappy_W(6, 267) <= 0; flappy_W(6, 268) <= 0; flappy_W(6, 269) <= 0; flappy_W(6, 270) <= 1; flappy_W(6, 271) <= 1; flappy_W(6, 272) <= 1; flappy_W(6, 273) <= 1; flappy_W(6, 274) <= 1; flappy_W(6, 275) <= 1; flappy_W(6, 276) <= 1; flappy_W(6, 277) <= 1; flappy_W(6, 278) <= 1; flappy_W(6, 279) <= 1; flappy_W(6, 280) <= 1; flappy_W(6, 281) <= 1; flappy_W(6, 282) <= 0; flappy_W(6, 283) <= 0; flappy_W(6, 284) <= 0; flappy_W(6, 285) <= 0; flappy_W(6, 286) <= 0; flappy_W(6, 287) <= 0; flappy_W(6, 288) <= 0; flappy_W(6, 289) <= 0; flappy_W(6, 290) <= 0; flappy_W(6, 291) <= 0; flappy_W(6, 292) <= 0; flappy_W(6, 293) <= 0; flappy_W(6, 294) <= 0; flappy_W(6, 295) <= 0; flappy_W(6, 296) <= 0; flappy_W(6, 297) <= 0; flappy_W(6, 298) <= 0; flappy_W(6, 299) <= 0; flappy_W(6, 300) <= 0; flappy_W(6, 301) <= 0; flappy_W(6, 302) <= 0; flappy_W(6, 303) <= 0; flappy_W(6, 304) <= 0; flappy_W(6, 305) <= 0; flappy_W(6, 306) <= 1; flappy_W(6, 307) <= 1; flappy_W(6, 308) <= 1; flappy_W(6, 309) <= 1; flappy_W(6, 310) <= 1; flappy_W(6, 311) <= 1; flappy_W(6, 312) <= 1; flappy_W(6, 313) <= 1; flappy_W(6, 314) <= 1; flappy_W(6, 315) <= 1; flappy_W(6, 316) <= 1; flappy_W(6, 317) <= 1; flappy_W(6, 318) <= 0; flappy_W(6, 319) <= 0; flappy_W(6, 320) <= 0; flappy_W(6, 321) <= 0; flappy_W(6, 322) <= 0; flappy_W(6, 323) <= 0; flappy_W(6, 324) <= 0; flappy_W(6, 325) <= 0; flappy_W(6, 326) <= 0; flappy_W(6, 327) <= 0; flappy_W(6, 328) <= 0; flappy_W(6, 329) <= 0; flappy_W(6, 330) <= 0; flappy_W(6, 331) <= 0; flappy_W(6, 332) <= 0; flappy_W(6, 333) <= 0; flappy_W(6, 334) <= 0; flappy_W(6, 335) <= 0; flappy_W(6, 336) <= 0; flappy_W(6, 337) <= 0; flappy_W(6, 338) <= 0; flappy_W(6, 339) <= 0; flappy_W(6, 340) <= 0; flappy_W(6, 341) <= 0; flappy_W(6, 342) <= 0; flappy_W(6, 343) <= 0; flappy_W(6, 344) <= 0; flappy_W(6, 345) <= 0; flappy_W(6, 346) <= 0; flappy_W(6, 347) <= 0; flappy_W(6, 348) <= 0; flappy_W(6, 349) <= 0; flappy_W(6, 350) <= 0; flappy_W(6, 351) <= 0; flappy_W(6, 352) <= 0; flappy_W(6, 353) <= 0; flappy_W(6, 354) <= 0; flappy_W(6, 355) <= 0; flappy_W(6, 356) <= 0; flappy_W(6, 357) <= 0; flappy_W(6, 358) <= 0; flappy_W(6, 359) <= 0; flappy_W(6, 360) <= 0; flappy_W(6, 361) <= 0; flappy_W(6, 362) <= 0; flappy_W(6, 363) <= 0; flappy_W(6, 364) <= 0; flappy_W(6, 365) <= 0; flappy_W(6, 366) <= 0; flappy_W(6, 367) <= 0; flappy_W(6, 368) <= 0; flappy_W(6, 369) <= 0; flappy_W(6, 370) <= 0; flappy_W(6, 371) <= 0; flappy_W(6, 372) <= 0; flappy_W(6, 373) <= 0; flappy_W(6, 374) <= 0; flappy_W(6, 375) <= 0; flappy_W(6, 376) <= 0; flappy_W(6, 377) <= 0; flappy_W(6, 378) <= 0; flappy_W(6, 379) <= 0; flappy_W(6, 380) <= 0; flappy_W(6, 381) <= 0; flappy_W(6, 382) <= 0; flappy_W(6, 383) <= 0; flappy_W(6, 384) <= 0; flappy_W(6, 385) <= 0; flappy_W(6, 386) <= 0; flappy_W(6, 387) <= 0; flappy_W(6, 388) <= 0; flappy_W(6, 389) <= 0; flappy_W(6, 390) <= 0; flappy_W(6, 391) <= 0; flappy_W(6, 392) <= 0; flappy_W(6, 393) <= 0; flappy_W(6, 394) <= 0; flappy_W(6, 395) <= 0; flappy_W(6, 396) <= 0; flappy_W(6, 397) <= 0; flappy_W(6, 398) <= 0; flappy_W(6, 399) <= 0; flappy_W(6, 400) <= 0; flappy_W(6, 401) <= 0; flappy_W(6, 402) <= 1; flappy_W(6, 403) <= 1; flappy_W(6, 404) <= 1; flappy_W(6, 405) <= 1; flappy_W(6, 406) <= 1; flappy_W(6, 407) <= 1; flappy_W(6, 408) <= 1; flappy_W(6, 409) <= 1; flappy_W(6, 410) <= 1; flappy_W(6, 411) <= 1; flappy_W(6, 412) <= 1; flappy_W(6, 413) <= 1; flappy_W(6, 414) <= 0; flappy_W(6, 415) <= 0; flappy_W(6, 416) <= 0; flappy_W(6, 417) <= 0; flappy_W(6, 418) <= 0; flappy_W(6, 419) <= 0; flappy_W(6, 420) <= 0; flappy_W(6, 421) <= 0; flappy_W(6, 422) <= 0; flappy_W(6, 423) <= 0; flappy_W(6, 424) <= 0; flappy_W(6, 425) <= 0; flappy_W(6, 426) <= 1; flappy_W(6, 427) <= 1; flappy_W(6, 428) <= 1; flappy_W(6, 429) <= 1; flappy_W(6, 430) <= 1; flappy_W(6, 431) <= 1; flappy_W(6, 432) <= 1; flappy_W(6, 433) <= 1; flappy_W(6, 434) <= 1; flappy_W(6, 435) <= 1; flappy_W(6, 436) <= 1; flappy_W(6, 437) <= 1; flappy_W(6, 438) <= 0; flappy_W(6, 439) <= 0; flappy_W(6, 440) <= 0; flappy_W(6, 441) <= 0; flappy_W(6, 442) <= 0; flappy_W(6, 443) <= 0; flappy_W(6, 444) <= 0; flappy_W(6, 445) <= 0; flappy_W(6, 446) <= 0; flappy_W(6, 447) <= 0; flappy_W(6, 448) <= 0; flappy_W(6, 449) <= 0; flappy_W(6, 450) <= 0; flappy_W(6, 451) <= 0; flappy_W(6, 452) <= 0; flappy_W(6, 453) <= 0; flappy_W(6, 454) <= 0; flappy_W(6, 455) <= 0; flappy_W(6, 456) <= 0; flappy_W(6, 457) <= 0; flappy_W(6, 458) <= 0; flappy_W(6, 459) <= 0; flappy_W(6, 460) <= 0; flappy_W(6, 461) <= 0; flappy_W(6, 462) <= 0; flappy_W(6, 463) <= 0; flappy_W(6, 464) <= 0; flappy_W(6, 465) <= 0; flappy_W(6, 466) <= 0; flappy_W(6, 467) <= 0; flappy_W(6, 468) <= 1; flappy_W(6, 469) <= 1; flappy_W(6, 470) <= 1; flappy_W(6, 471) <= 1; flappy_W(6, 472) <= 1; flappy_W(6, 473) <= 1; flappy_W(6, 474) <= 1; flappy_W(6, 475) <= 1; flappy_W(6, 476) <= 1; flappy_W(6, 477) <= 1; flappy_W(6, 478) <= 1; flappy_W(6, 479) <= 1; flappy_W(6, 480) <= 0; flappy_W(6, 481) <= 0; flappy_W(6, 482) <= 0; flappy_W(6, 483) <= 0; flappy_W(6, 484) <= 0; flappy_W(6, 485) <= 0; flappy_W(6, 486) <= 0; flappy_W(6, 487) <= 0; flappy_W(6, 488) <= 0; flappy_W(6, 489) <= 0; flappy_W(6, 490) <= 0; flappy_W(6, 491) <= 0; flappy_W(6, 492) <= 0; flappy_W(6, 493) <= 0; flappy_W(6, 494) <= 0; flappy_W(6, 495) <= 0; flappy_W(6, 496) <= 0; flappy_W(6, 497) <= 0; flappy_W(6, 498) <= 0; flappy_W(6, 499) <= 0; flappy_W(6, 500) <= 0; flappy_W(6, 501) <= 0; flappy_W(6, 502) <= 0; flappy_W(6, 503) <= 0; flappy_W(6, 504) <= 0; flappy_W(6, 505) <= 0; flappy_W(6, 506) <= 0; flappy_W(6, 507) <= 0; flappy_W(6, 508) <= 0; flappy_W(6, 509) <= 0; flappy_W(6, 510) <= 1; flappy_W(6, 511) <= 1; flappy_W(6, 512) <= 1; flappy_W(6, 513) <= 1; flappy_W(6, 514) <= 1; flappy_W(6, 515) <= 1; flappy_W(6, 516) <= 1; flappy_W(6, 517) <= 1; flappy_W(6, 518) <= 1; flappy_W(6, 519) <= 1; flappy_W(6, 520) <= 1; flappy_W(6, 521) <= 1; flappy_W(6, 522) <= 0; flappy_W(6, 523) <= 0; flappy_W(6, 524) <= 0; flappy_W(6, 525) <= 0; flappy_W(6, 526) <= 0; flappy_W(6, 527) <= 0; flappy_W(6, 528) <= 0; flappy_W(6, 529) <= 0; flappy_W(6, 530) <= 0; flappy_W(6, 531) <= 0; flappy_W(6, 532) <= 0; flappy_W(6, 533) <= 0; flappy_W(6, 534) <= 1; flappy_W(6, 535) <= 1; flappy_W(6, 536) <= 1; flappy_W(6, 537) <= 1; flappy_W(6, 538) <= 1; flappy_W(6, 539) <= 1; flappy_W(6, 540) <= 1; flappy_W(6, 541) <= 1; flappy_W(6, 542) <= 1; flappy_W(6, 543) <= 1; flappy_W(6, 544) <= 1; flappy_W(6, 545) <= 1; flappy_W(6, 546) <= 0; flappy_W(6, 547) <= 0; flappy_W(6, 548) <= 0; flappy_W(6, 549) <= 0; flappy_W(6, 550) <= 0; flappy_W(6, 551) <= 0; flappy_W(6, 552) <= 0; flappy_W(6, 553) <= 0; flappy_W(6, 554) <= 0; flappy_W(6, 555) <= 0; flappy_W(6, 556) <= 0; flappy_W(6, 557) <= 0; flappy_W(6, 558) <= 0; flappy_W(6, 559) <= 0; flappy_W(6, 560) <= 0; flappy_W(6, 561) <= 0; flappy_W(6, 562) <= 0; flappy_W(6, 563) <= 0; flappy_W(6, 564) <= 1; flappy_W(6, 565) <= 1; flappy_W(6, 566) <= 1; flappy_W(6, 567) <= 1; flappy_W(6, 568) <= 1; flappy_W(6, 569) <= 1; flappy_W(6, 570) <= 1; flappy_W(6, 571) <= 1; flappy_W(6, 572) <= 1; flappy_W(6, 573) <= 1; flappy_W(6, 574) <= 1; flappy_W(6, 575) <= 1; flappy_W(6, 576) <= 0; flappy_W(6, 577) <= 0; flappy_W(6, 578) <= 0; flappy_W(6, 579) <= 0; flappy_W(6, 580) <= 0; flappy_W(6, 581) <= 0; flappy_W(6, 582) <= 1; flappy_W(6, 583) <= 1; flappy_W(6, 584) <= 1; flappy_W(6, 585) <= 1; flappy_W(6, 586) <= 1; flappy_W(6, 587) <= 1; flappy_W(6, 588) <= 1; flappy_W(6, 589) <= 1; flappy_W(6, 590) <= 1; flappy_W(6, 591) <= 1; flappy_W(6, 592) <= 1; flappy_W(6, 593) <= 1; 
flappy_W(7, 0) <= 0; flappy_W(7, 1) <= 0; flappy_W(7, 2) <= 0; flappy_W(7, 3) <= 0; flappy_W(7, 4) <= 0; flappy_W(7, 5) <= 0; flappy_W(7, 6) <= 1; flappy_W(7, 7) <= 1; flappy_W(7, 8) <= 1; flappy_W(7, 9) <= 1; flappy_W(7, 10) <= 1; flappy_W(7, 11) <= 1; flappy_W(7, 12) <= 1; flappy_W(7, 13) <= 1; flappy_W(7, 14) <= 1; flappy_W(7, 15) <= 1; flappy_W(7, 16) <= 1; flappy_W(7, 17) <= 1; flappy_W(7, 18) <= 0; flappy_W(7, 19) <= 0; flappy_W(7, 20) <= 0; flappy_W(7, 21) <= 0; flappy_W(7, 22) <= 0; flappy_W(7, 23) <= 0; flappy_W(7, 24) <= 0; flappy_W(7, 25) <= 0; flappy_W(7, 26) <= 0; flappy_W(7, 27) <= 0; flappy_W(7, 28) <= 0; flappy_W(7, 29) <= 0; flappy_W(7, 30) <= 1; flappy_W(7, 31) <= 1; flappy_W(7, 32) <= 1; flappy_W(7, 33) <= 1; flappy_W(7, 34) <= 1; flappy_W(7, 35) <= 1; flappy_W(7, 36) <= 1; flappy_W(7, 37) <= 1; flappy_W(7, 38) <= 1; flappy_W(7, 39) <= 1; flappy_W(7, 40) <= 1; flappy_W(7, 41) <= 1; flappy_W(7, 42) <= 0; flappy_W(7, 43) <= 0; flappy_W(7, 44) <= 0; flappy_W(7, 45) <= 0; flappy_W(7, 46) <= 0; flappy_W(7, 47) <= 0; flappy_W(7, 48) <= 0; flappy_W(7, 49) <= 0; flappy_W(7, 50) <= 0; flappy_W(7, 51) <= 0; flappy_W(7, 52) <= 0; flappy_W(7, 53) <= 0; flappy_W(7, 54) <= 0; flappy_W(7, 55) <= 0; flappy_W(7, 56) <= 0; flappy_W(7, 57) <= 0; flappy_W(7, 58) <= 0; flappy_W(7, 59) <= 0; flappy_W(7, 60) <= 1; flappy_W(7, 61) <= 1; flappy_W(7, 62) <= 1; flappy_W(7, 63) <= 1; flappy_W(7, 64) <= 1; flappy_W(7, 65) <= 1; flappy_W(7, 66) <= 1; flappy_W(7, 67) <= 1; flappy_W(7, 68) <= 1; flappy_W(7, 69) <= 1; flappy_W(7, 70) <= 1; flappy_W(7, 71) <= 1; flappy_W(7, 72) <= 0; flappy_W(7, 73) <= 0; flappy_W(7, 74) <= 0; flappy_W(7, 75) <= 0; flappy_W(7, 76) <= 0; flappy_W(7, 77) <= 0; flappy_W(7, 78) <= 0; flappy_W(7, 79) <= 0; flappy_W(7, 80) <= 0; flappy_W(7, 81) <= 0; flappy_W(7, 82) <= 0; flappy_W(7, 83) <= 0; flappy_W(7, 84) <= 0; flappy_W(7, 85) <= 0; flappy_W(7, 86) <= 0; flappy_W(7, 87) <= 0; flappy_W(7, 88) <= 0; flappy_W(7, 89) <= 0; flappy_W(7, 90) <= 0; flappy_W(7, 91) <= 0; flappy_W(7, 92) <= 0; flappy_W(7, 93) <= 0; flappy_W(7, 94) <= 0; flappy_W(7, 95) <= 0; flappy_W(7, 96) <= 0; flappy_W(7, 97) <= 0; flappy_W(7, 98) <= 0; flappy_W(7, 99) <= 0; flappy_W(7, 100) <= 0; flappy_W(7, 101) <= 0; flappy_W(7, 102) <= 0; flappy_W(7, 103) <= 0; flappy_W(7, 104) <= 0; flappy_W(7, 105) <= 0; flappy_W(7, 106) <= 0; flappy_W(7, 107) <= 0; flappy_W(7, 108) <= 0; flappy_W(7, 109) <= 0; flappy_W(7, 110) <= 0; flappy_W(7, 111) <= 0; flappy_W(7, 112) <= 0; flappy_W(7, 113) <= 0; flappy_W(7, 114) <= 0; flappy_W(7, 115) <= 0; flappy_W(7, 116) <= 0; flappy_W(7, 117) <= 0; flappy_W(7, 118) <= 0; flappy_W(7, 119) <= 0; flappy_W(7, 120) <= 1; flappy_W(7, 121) <= 1; flappy_W(7, 122) <= 1; flappy_W(7, 123) <= 1; flappy_W(7, 124) <= 1; flappy_W(7, 125) <= 1; flappy_W(7, 126) <= 1; flappy_W(7, 127) <= 1; flappy_W(7, 128) <= 1; flappy_W(7, 129) <= 1; flappy_W(7, 130) <= 1; flappy_W(7, 131) <= 1; flappy_W(7, 132) <= 1; flappy_W(7, 133) <= 1; flappy_W(7, 134) <= 1; flappy_W(7, 135) <= 1; flappy_W(7, 136) <= 1; flappy_W(7, 137) <= 1; flappy_W(7, 138) <= 0; flappy_W(7, 139) <= 0; flappy_W(7, 140) <= 0; flappy_W(7, 141) <= 0; flappy_W(7, 142) <= 0; flappy_W(7, 143) <= 0; flappy_W(7, 144) <= 0; flappy_W(7, 145) <= 0; flappy_W(7, 146) <= 0; flappy_W(7, 147) <= 0; flappy_W(7, 148) <= 0; flappy_W(7, 149) <= 0; flappy_W(7, 150) <= 0; flappy_W(7, 151) <= 0; flappy_W(7, 152) <= 0; flappy_W(7, 153) <= 0; flappy_W(7, 154) <= 0; flappy_W(7, 155) <= 0; flappy_W(7, 156) <= 0; flappy_W(7, 157) <= 0; flappy_W(7, 158) <= 0; flappy_W(7, 159) <= 0; flappy_W(7, 160) <= 0; flappy_W(7, 161) <= 0; flappy_W(7, 162) <= 0; flappy_W(7, 163) <= 0; flappy_W(7, 164) <= 0; flappy_W(7, 165) <= 0; flappy_W(7, 166) <= 0; flappy_W(7, 167) <= 0; flappy_W(7, 168) <= 1; flappy_W(7, 169) <= 1; flappy_W(7, 170) <= 1; flappy_W(7, 171) <= 1; flappy_W(7, 172) <= 1; flappy_W(7, 173) <= 1; flappy_W(7, 174) <= 1; flappy_W(7, 175) <= 1; flappy_W(7, 176) <= 1; flappy_W(7, 177) <= 1; flappy_W(7, 178) <= 1; flappy_W(7, 179) <= 1; flappy_W(7, 180) <= 0; flappy_W(7, 181) <= 0; flappy_W(7, 182) <= 0; flappy_W(7, 183) <= 0; flappy_W(7, 184) <= 0; flappy_W(7, 185) <= 0; flappy_W(7, 186) <= 0; flappy_W(7, 187) <= 0; flappy_W(7, 188) <= 0; flappy_W(7, 189) <= 0; flappy_W(7, 190) <= 0; flappy_W(7, 191) <= 0; flappy_W(7, 192) <= 1; flappy_W(7, 193) <= 1; flappy_W(7, 194) <= 1; flappy_W(7, 195) <= 1; flappy_W(7, 196) <= 1; flappy_W(7, 197) <= 1; flappy_W(7, 198) <= 1; flappy_W(7, 199) <= 1; flappy_W(7, 200) <= 1; flappy_W(7, 201) <= 1; flappy_W(7, 202) <= 1; flappy_W(7, 203) <= 1; flappy_W(7, 204) <= 0; flappy_W(7, 205) <= 0; flappy_W(7, 206) <= 0; flappy_W(7, 207) <= 0; flappy_W(7, 208) <= 0; flappy_W(7, 209) <= 0; flappy_W(7, 210) <= 0; flappy_W(7, 211) <= 0; flappy_W(7, 212) <= 0; flappy_W(7, 213) <= 0; flappy_W(7, 214) <= 0; flappy_W(7, 215) <= 0; flappy_W(7, 216) <= 0; flappy_W(7, 217) <= 0; flappy_W(7, 218) <= 0; flappy_W(7, 219) <= 0; flappy_W(7, 220) <= 0; flappy_W(7, 221) <= 0; flappy_W(7, 222) <= 1; flappy_W(7, 223) <= 1; flappy_W(7, 224) <= 1; flappy_W(7, 225) <= 1; flappy_W(7, 226) <= 1; flappy_W(7, 227) <= 1; flappy_W(7, 228) <= 1; flappy_W(7, 229) <= 1; flappy_W(7, 230) <= 1; flappy_W(7, 231) <= 1; flappy_W(7, 232) <= 1; flappy_W(7, 233) <= 1; flappy_W(7, 234) <= 0; flappy_W(7, 235) <= 0; flappy_W(7, 236) <= 0; flappy_W(7, 237) <= 0; flappy_W(7, 238) <= 0; flappy_W(7, 239) <= 0; flappy_W(7, 240) <= 0; flappy_W(7, 241) <= 0; flappy_W(7, 242) <= 0; flappy_W(7, 243) <= 0; flappy_W(7, 244) <= 0; flappy_W(7, 245) <= 0; flappy_W(7, 246) <= 1; flappy_W(7, 247) <= 1; flappy_W(7, 248) <= 1; flappy_W(7, 249) <= 1; flappy_W(7, 250) <= 1; flappy_W(7, 251) <= 1; flappy_W(7, 252) <= 1; flappy_W(7, 253) <= 1; flappy_W(7, 254) <= 1; flappy_W(7, 255) <= 1; flappy_W(7, 256) <= 1; flappy_W(7, 257) <= 1; flappy_W(7, 258) <= 0; flappy_W(7, 259) <= 0; flappy_W(7, 260) <= 0; flappy_W(7, 261) <= 0; flappy_W(7, 262) <= 0; flappy_W(7, 263) <= 0; flappy_W(7, 264) <= 0; flappy_W(7, 265) <= 0; flappy_W(7, 266) <= 0; flappy_W(7, 267) <= 0; flappy_W(7, 268) <= 0; flappy_W(7, 269) <= 0; flappy_W(7, 270) <= 1; flappy_W(7, 271) <= 1; flappy_W(7, 272) <= 1; flappy_W(7, 273) <= 1; flappy_W(7, 274) <= 1; flappy_W(7, 275) <= 1; flappy_W(7, 276) <= 1; flappy_W(7, 277) <= 1; flappy_W(7, 278) <= 1; flappy_W(7, 279) <= 1; flappy_W(7, 280) <= 1; flappy_W(7, 281) <= 1; flappy_W(7, 282) <= 0; flappy_W(7, 283) <= 0; flappy_W(7, 284) <= 0; flappy_W(7, 285) <= 0; flappy_W(7, 286) <= 0; flappy_W(7, 287) <= 0; flappy_W(7, 288) <= 0; flappy_W(7, 289) <= 0; flappy_W(7, 290) <= 0; flappy_W(7, 291) <= 0; flappy_W(7, 292) <= 0; flappy_W(7, 293) <= 0; flappy_W(7, 294) <= 0; flappy_W(7, 295) <= 0; flappy_W(7, 296) <= 0; flappy_W(7, 297) <= 0; flappy_W(7, 298) <= 0; flappy_W(7, 299) <= 0; flappy_W(7, 300) <= 0; flappy_W(7, 301) <= 0; flappy_W(7, 302) <= 0; flappy_W(7, 303) <= 0; flappy_W(7, 304) <= 0; flappy_W(7, 305) <= 0; flappy_W(7, 306) <= 1; flappy_W(7, 307) <= 1; flappy_W(7, 308) <= 1; flappy_W(7, 309) <= 1; flappy_W(7, 310) <= 1; flappy_W(7, 311) <= 1; flappy_W(7, 312) <= 1; flappy_W(7, 313) <= 1; flappy_W(7, 314) <= 1; flappy_W(7, 315) <= 1; flappy_W(7, 316) <= 1; flappy_W(7, 317) <= 1; flappy_W(7, 318) <= 0; flappy_W(7, 319) <= 0; flappy_W(7, 320) <= 0; flappy_W(7, 321) <= 0; flappy_W(7, 322) <= 0; flappy_W(7, 323) <= 0; flappy_W(7, 324) <= 0; flappy_W(7, 325) <= 0; flappy_W(7, 326) <= 0; flappy_W(7, 327) <= 0; flappy_W(7, 328) <= 0; flappy_W(7, 329) <= 0; flappy_W(7, 330) <= 0; flappy_W(7, 331) <= 0; flappy_W(7, 332) <= 0; flappy_W(7, 333) <= 0; flappy_W(7, 334) <= 0; flappy_W(7, 335) <= 0; flappy_W(7, 336) <= 0; flappy_W(7, 337) <= 0; flappy_W(7, 338) <= 0; flappy_W(7, 339) <= 0; flappy_W(7, 340) <= 0; flappy_W(7, 341) <= 0; flappy_W(7, 342) <= 0; flappy_W(7, 343) <= 0; flappy_W(7, 344) <= 0; flappy_W(7, 345) <= 0; flappy_W(7, 346) <= 0; flappy_W(7, 347) <= 0; flappy_W(7, 348) <= 0; flappy_W(7, 349) <= 0; flappy_W(7, 350) <= 0; flappy_W(7, 351) <= 0; flappy_W(7, 352) <= 0; flappy_W(7, 353) <= 0; flappy_W(7, 354) <= 0; flappy_W(7, 355) <= 0; flappy_W(7, 356) <= 0; flappy_W(7, 357) <= 0; flappy_W(7, 358) <= 0; flappy_W(7, 359) <= 0; flappy_W(7, 360) <= 0; flappy_W(7, 361) <= 0; flappy_W(7, 362) <= 0; flappy_W(7, 363) <= 0; flappy_W(7, 364) <= 0; flappy_W(7, 365) <= 0; flappy_W(7, 366) <= 0; flappy_W(7, 367) <= 0; flappy_W(7, 368) <= 0; flappy_W(7, 369) <= 0; flappy_W(7, 370) <= 0; flappy_W(7, 371) <= 0; flappy_W(7, 372) <= 0; flappy_W(7, 373) <= 0; flappy_W(7, 374) <= 0; flappy_W(7, 375) <= 0; flappy_W(7, 376) <= 0; flappy_W(7, 377) <= 0; flappy_W(7, 378) <= 0; flappy_W(7, 379) <= 0; flappy_W(7, 380) <= 0; flappy_W(7, 381) <= 0; flappy_W(7, 382) <= 0; flappy_W(7, 383) <= 0; flappy_W(7, 384) <= 0; flappy_W(7, 385) <= 0; flappy_W(7, 386) <= 0; flappy_W(7, 387) <= 0; flappy_W(7, 388) <= 0; flappy_W(7, 389) <= 0; flappy_W(7, 390) <= 0; flappy_W(7, 391) <= 0; flappy_W(7, 392) <= 0; flappy_W(7, 393) <= 0; flappy_W(7, 394) <= 0; flappy_W(7, 395) <= 0; flappy_W(7, 396) <= 0; flappy_W(7, 397) <= 0; flappy_W(7, 398) <= 0; flappy_W(7, 399) <= 0; flappy_W(7, 400) <= 0; flappy_W(7, 401) <= 0; flappy_W(7, 402) <= 1; flappy_W(7, 403) <= 1; flappy_W(7, 404) <= 1; flappy_W(7, 405) <= 1; flappy_W(7, 406) <= 1; flappy_W(7, 407) <= 1; flappy_W(7, 408) <= 1; flappy_W(7, 409) <= 1; flappy_W(7, 410) <= 1; flappy_W(7, 411) <= 1; flappy_W(7, 412) <= 1; flappy_W(7, 413) <= 1; flappy_W(7, 414) <= 0; flappy_W(7, 415) <= 0; flappy_W(7, 416) <= 0; flappy_W(7, 417) <= 0; flappy_W(7, 418) <= 0; flappy_W(7, 419) <= 0; flappy_W(7, 420) <= 0; flappy_W(7, 421) <= 0; flappy_W(7, 422) <= 0; flappy_W(7, 423) <= 0; flappy_W(7, 424) <= 0; flappy_W(7, 425) <= 0; flappy_W(7, 426) <= 1; flappy_W(7, 427) <= 1; flappy_W(7, 428) <= 1; flappy_W(7, 429) <= 1; flappy_W(7, 430) <= 1; flappy_W(7, 431) <= 1; flappy_W(7, 432) <= 1; flappy_W(7, 433) <= 1; flappy_W(7, 434) <= 1; flappy_W(7, 435) <= 1; flappy_W(7, 436) <= 1; flappy_W(7, 437) <= 1; flappy_W(7, 438) <= 0; flappy_W(7, 439) <= 0; flappy_W(7, 440) <= 0; flappy_W(7, 441) <= 0; flappy_W(7, 442) <= 0; flappy_W(7, 443) <= 0; flappy_W(7, 444) <= 0; flappy_W(7, 445) <= 0; flappy_W(7, 446) <= 0; flappy_W(7, 447) <= 0; flappy_W(7, 448) <= 0; flappy_W(7, 449) <= 0; flappy_W(7, 450) <= 0; flappy_W(7, 451) <= 0; flappy_W(7, 452) <= 0; flappy_W(7, 453) <= 0; flappy_W(7, 454) <= 0; flappy_W(7, 455) <= 0; flappy_W(7, 456) <= 0; flappy_W(7, 457) <= 0; flappy_W(7, 458) <= 0; flappy_W(7, 459) <= 0; flappy_W(7, 460) <= 0; flappy_W(7, 461) <= 0; flappy_W(7, 462) <= 0; flappy_W(7, 463) <= 0; flappy_W(7, 464) <= 0; flappy_W(7, 465) <= 0; flappy_W(7, 466) <= 0; flappy_W(7, 467) <= 0; flappy_W(7, 468) <= 1; flappy_W(7, 469) <= 1; flappy_W(7, 470) <= 1; flappy_W(7, 471) <= 1; flappy_W(7, 472) <= 1; flappy_W(7, 473) <= 1; flappy_W(7, 474) <= 1; flappy_W(7, 475) <= 1; flappy_W(7, 476) <= 1; flappy_W(7, 477) <= 1; flappy_W(7, 478) <= 1; flappy_W(7, 479) <= 1; flappy_W(7, 480) <= 0; flappy_W(7, 481) <= 0; flappy_W(7, 482) <= 0; flappy_W(7, 483) <= 0; flappy_W(7, 484) <= 0; flappy_W(7, 485) <= 0; flappy_W(7, 486) <= 0; flappy_W(7, 487) <= 0; flappy_W(7, 488) <= 0; flappy_W(7, 489) <= 0; flappy_W(7, 490) <= 0; flappy_W(7, 491) <= 0; flappy_W(7, 492) <= 0; flappy_W(7, 493) <= 0; flappy_W(7, 494) <= 0; flappy_W(7, 495) <= 0; flappy_W(7, 496) <= 0; flappy_W(7, 497) <= 0; flappy_W(7, 498) <= 0; flappy_W(7, 499) <= 0; flappy_W(7, 500) <= 0; flappy_W(7, 501) <= 0; flappy_W(7, 502) <= 0; flappy_W(7, 503) <= 0; flappy_W(7, 504) <= 0; flappy_W(7, 505) <= 0; flappy_W(7, 506) <= 0; flappy_W(7, 507) <= 0; flappy_W(7, 508) <= 0; flappy_W(7, 509) <= 0; flappy_W(7, 510) <= 1; flappy_W(7, 511) <= 1; flappy_W(7, 512) <= 1; flappy_W(7, 513) <= 1; flappy_W(7, 514) <= 1; flappy_W(7, 515) <= 1; flappy_W(7, 516) <= 1; flappy_W(7, 517) <= 1; flappy_W(7, 518) <= 1; flappy_W(7, 519) <= 1; flappy_W(7, 520) <= 1; flappy_W(7, 521) <= 1; flappy_W(7, 522) <= 0; flappy_W(7, 523) <= 0; flappy_W(7, 524) <= 0; flappy_W(7, 525) <= 0; flappy_W(7, 526) <= 0; flappy_W(7, 527) <= 0; flappy_W(7, 528) <= 0; flappy_W(7, 529) <= 0; flappy_W(7, 530) <= 0; flappy_W(7, 531) <= 0; flappy_W(7, 532) <= 0; flappy_W(7, 533) <= 0; flappy_W(7, 534) <= 1; flappy_W(7, 535) <= 1; flappy_W(7, 536) <= 1; flappy_W(7, 537) <= 1; flappy_W(7, 538) <= 1; flappy_W(7, 539) <= 1; flappy_W(7, 540) <= 1; flappy_W(7, 541) <= 1; flappy_W(7, 542) <= 1; flappy_W(7, 543) <= 1; flappy_W(7, 544) <= 1; flappy_W(7, 545) <= 1; flappy_W(7, 546) <= 0; flappy_W(7, 547) <= 0; flappy_W(7, 548) <= 0; flappy_W(7, 549) <= 0; flappy_W(7, 550) <= 0; flappy_W(7, 551) <= 0; flappy_W(7, 552) <= 0; flappy_W(7, 553) <= 0; flappy_W(7, 554) <= 0; flappy_W(7, 555) <= 0; flappy_W(7, 556) <= 0; flappy_W(7, 557) <= 0; flappy_W(7, 558) <= 0; flappy_W(7, 559) <= 0; flappy_W(7, 560) <= 0; flappy_W(7, 561) <= 0; flappy_W(7, 562) <= 0; flappy_W(7, 563) <= 0; flappy_W(7, 564) <= 1; flappy_W(7, 565) <= 1; flappy_W(7, 566) <= 1; flappy_W(7, 567) <= 1; flappy_W(7, 568) <= 1; flappy_W(7, 569) <= 1; flappy_W(7, 570) <= 1; flappy_W(7, 571) <= 1; flappy_W(7, 572) <= 1; flappy_W(7, 573) <= 1; flappy_W(7, 574) <= 1; flappy_W(7, 575) <= 1; flappy_W(7, 576) <= 0; flappy_W(7, 577) <= 0; flappy_W(7, 578) <= 0; flappy_W(7, 579) <= 0; flappy_W(7, 580) <= 0; flappy_W(7, 581) <= 0; flappy_W(7, 582) <= 1; flappy_W(7, 583) <= 1; flappy_W(7, 584) <= 1; flappy_W(7, 585) <= 1; flappy_W(7, 586) <= 1; flappy_W(7, 587) <= 1; flappy_W(7, 588) <= 1; flappy_W(7, 589) <= 1; flappy_W(7, 590) <= 1; flappy_W(7, 591) <= 1; flappy_W(7, 592) <= 1; flappy_W(7, 593) <= 1; 
flappy_W(8, 0) <= 0; flappy_W(8, 1) <= 0; flappy_W(8, 2) <= 0; flappy_W(8, 3) <= 0; flappy_W(8, 4) <= 0; flappy_W(8, 5) <= 0; flappy_W(8, 6) <= 1; flappy_W(8, 7) <= 1; flappy_W(8, 8) <= 1; flappy_W(8, 9) <= 1; flappy_W(8, 10) <= 1; flappy_W(8, 11) <= 1; flappy_W(8, 12) <= 1; flappy_W(8, 13) <= 1; flappy_W(8, 14) <= 1; flappy_W(8, 15) <= 1; flappy_W(8, 16) <= 1; flappy_W(8, 17) <= 1; flappy_W(8, 18) <= 0; flappy_W(8, 19) <= 0; flappy_W(8, 20) <= 0; flappy_W(8, 21) <= 0; flappy_W(8, 22) <= 0; flappy_W(8, 23) <= 0; flappy_W(8, 24) <= 0; flappy_W(8, 25) <= 0; flappy_W(8, 26) <= 0; flappy_W(8, 27) <= 0; flappy_W(8, 28) <= 0; flappy_W(8, 29) <= 0; flappy_W(8, 30) <= 1; flappy_W(8, 31) <= 1; flappy_W(8, 32) <= 1; flappy_W(8, 33) <= 1; flappy_W(8, 34) <= 1; flappy_W(8, 35) <= 1; flappy_W(8, 36) <= 1; flappy_W(8, 37) <= 1; flappy_W(8, 38) <= 1; flappy_W(8, 39) <= 1; flappy_W(8, 40) <= 1; flappy_W(8, 41) <= 1; flappy_W(8, 42) <= 0; flappy_W(8, 43) <= 0; flappy_W(8, 44) <= 0; flappy_W(8, 45) <= 0; flappy_W(8, 46) <= 0; flappy_W(8, 47) <= 0; flappy_W(8, 48) <= 0; flappy_W(8, 49) <= 0; flappy_W(8, 50) <= 0; flappy_W(8, 51) <= 0; flappy_W(8, 52) <= 0; flappy_W(8, 53) <= 0; flappy_W(8, 54) <= 0; flappy_W(8, 55) <= 0; flappy_W(8, 56) <= 0; flappy_W(8, 57) <= 0; flappy_W(8, 58) <= 0; flappy_W(8, 59) <= 0; flappy_W(8, 60) <= 1; flappy_W(8, 61) <= 1; flappy_W(8, 62) <= 1; flappy_W(8, 63) <= 1; flappy_W(8, 64) <= 1; flappy_W(8, 65) <= 1; flappy_W(8, 66) <= 1; flappy_W(8, 67) <= 1; flappy_W(8, 68) <= 1; flappy_W(8, 69) <= 1; flappy_W(8, 70) <= 1; flappy_W(8, 71) <= 1; flappy_W(8, 72) <= 0; flappy_W(8, 73) <= 0; flappy_W(8, 74) <= 0; flappy_W(8, 75) <= 0; flappy_W(8, 76) <= 0; flappy_W(8, 77) <= 0; flappy_W(8, 78) <= 0; flappy_W(8, 79) <= 0; flappy_W(8, 80) <= 0; flappy_W(8, 81) <= 0; flappy_W(8, 82) <= 0; flappy_W(8, 83) <= 0; flappy_W(8, 84) <= 0; flappy_W(8, 85) <= 0; flappy_W(8, 86) <= 0; flappy_W(8, 87) <= 0; flappy_W(8, 88) <= 0; flappy_W(8, 89) <= 0; flappy_W(8, 90) <= 0; flappy_W(8, 91) <= 0; flappy_W(8, 92) <= 0; flappy_W(8, 93) <= 0; flappy_W(8, 94) <= 0; flappy_W(8, 95) <= 0; flappy_W(8, 96) <= 0; flappy_W(8, 97) <= 0; flappy_W(8, 98) <= 0; flappy_W(8, 99) <= 0; flappy_W(8, 100) <= 0; flappy_W(8, 101) <= 0; flappy_W(8, 102) <= 0; flappy_W(8, 103) <= 0; flappy_W(8, 104) <= 0; flappy_W(8, 105) <= 0; flappy_W(8, 106) <= 0; flappy_W(8, 107) <= 0; flappy_W(8, 108) <= 0; flappy_W(8, 109) <= 0; flappy_W(8, 110) <= 0; flappy_W(8, 111) <= 0; flappy_W(8, 112) <= 0; flappy_W(8, 113) <= 0; flappy_W(8, 114) <= 0; flappy_W(8, 115) <= 0; flappy_W(8, 116) <= 0; flappy_W(8, 117) <= 0; flappy_W(8, 118) <= 0; flappy_W(8, 119) <= 0; flappy_W(8, 120) <= 1; flappy_W(8, 121) <= 1; flappy_W(8, 122) <= 1; flappy_W(8, 123) <= 1; flappy_W(8, 124) <= 1; flappy_W(8, 125) <= 1; flappy_W(8, 126) <= 1; flappy_W(8, 127) <= 1; flappy_W(8, 128) <= 1; flappy_W(8, 129) <= 1; flappy_W(8, 130) <= 1; flappy_W(8, 131) <= 1; flappy_W(8, 132) <= 1; flappy_W(8, 133) <= 1; flappy_W(8, 134) <= 1; flappy_W(8, 135) <= 1; flappy_W(8, 136) <= 1; flappy_W(8, 137) <= 1; flappy_W(8, 138) <= 0; flappy_W(8, 139) <= 0; flappy_W(8, 140) <= 0; flappy_W(8, 141) <= 0; flappy_W(8, 142) <= 0; flappy_W(8, 143) <= 0; flappy_W(8, 144) <= 0; flappy_W(8, 145) <= 0; flappy_W(8, 146) <= 0; flappy_W(8, 147) <= 0; flappy_W(8, 148) <= 0; flappy_W(8, 149) <= 0; flappy_W(8, 150) <= 0; flappy_W(8, 151) <= 0; flappy_W(8, 152) <= 0; flappy_W(8, 153) <= 0; flappy_W(8, 154) <= 0; flappy_W(8, 155) <= 0; flappy_W(8, 156) <= 0; flappy_W(8, 157) <= 0; flappy_W(8, 158) <= 0; flappy_W(8, 159) <= 0; flappy_W(8, 160) <= 0; flappy_W(8, 161) <= 0; flappy_W(8, 162) <= 0; flappy_W(8, 163) <= 0; flappy_W(8, 164) <= 0; flappy_W(8, 165) <= 0; flappy_W(8, 166) <= 0; flappy_W(8, 167) <= 0; flappy_W(8, 168) <= 1; flappy_W(8, 169) <= 1; flappy_W(8, 170) <= 1; flappy_W(8, 171) <= 1; flappy_W(8, 172) <= 1; flappy_W(8, 173) <= 1; flappy_W(8, 174) <= 1; flappy_W(8, 175) <= 1; flappy_W(8, 176) <= 1; flappy_W(8, 177) <= 1; flappy_W(8, 178) <= 1; flappy_W(8, 179) <= 1; flappy_W(8, 180) <= 0; flappy_W(8, 181) <= 0; flappy_W(8, 182) <= 0; flappy_W(8, 183) <= 0; flappy_W(8, 184) <= 0; flappy_W(8, 185) <= 0; flappy_W(8, 186) <= 0; flappy_W(8, 187) <= 0; flappy_W(8, 188) <= 0; flappy_W(8, 189) <= 0; flappy_W(8, 190) <= 0; flappy_W(8, 191) <= 0; flappy_W(8, 192) <= 1; flappy_W(8, 193) <= 1; flappy_W(8, 194) <= 1; flappy_W(8, 195) <= 1; flappy_W(8, 196) <= 1; flappy_W(8, 197) <= 1; flappy_W(8, 198) <= 1; flappy_W(8, 199) <= 1; flappy_W(8, 200) <= 1; flappy_W(8, 201) <= 1; flappy_W(8, 202) <= 1; flappy_W(8, 203) <= 1; flappy_W(8, 204) <= 0; flappy_W(8, 205) <= 0; flappy_W(8, 206) <= 0; flappy_W(8, 207) <= 0; flappy_W(8, 208) <= 0; flappy_W(8, 209) <= 0; flappy_W(8, 210) <= 0; flappy_W(8, 211) <= 0; flappy_W(8, 212) <= 0; flappy_W(8, 213) <= 0; flappy_W(8, 214) <= 0; flappy_W(8, 215) <= 0; flappy_W(8, 216) <= 0; flappy_W(8, 217) <= 0; flappy_W(8, 218) <= 0; flappy_W(8, 219) <= 0; flappy_W(8, 220) <= 0; flappy_W(8, 221) <= 0; flappy_W(8, 222) <= 1; flappy_W(8, 223) <= 1; flappy_W(8, 224) <= 1; flappy_W(8, 225) <= 1; flappy_W(8, 226) <= 1; flappy_W(8, 227) <= 1; flappy_W(8, 228) <= 1; flappy_W(8, 229) <= 1; flappy_W(8, 230) <= 1; flappy_W(8, 231) <= 1; flappy_W(8, 232) <= 1; flappy_W(8, 233) <= 1; flappy_W(8, 234) <= 0; flappy_W(8, 235) <= 0; flappy_W(8, 236) <= 0; flappy_W(8, 237) <= 0; flappy_W(8, 238) <= 0; flappy_W(8, 239) <= 0; flappy_W(8, 240) <= 0; flappy_W(8, 241) <= 0; flappy_W(8, 242) <= 0; flappy_W(8, 243) <= 0; flappy_W(8, 244) <= 0; flappy_W(8, 245) <= 0; flappy_W(8, 246) <= 1; flappy_W(8, 247) <= 1; flappy_W(8, 248) <= 1; flappy_W(8, 249) <= 1; flappy_W(8, 250) <= 1; flappy_W(8, 251) <= 1; flappy_W(8, 252) <= 1; flappy_W(8, 253) <= 1; flappy_W(8, 254) <= 1; flappy_W(8, 255) <= 1; flappy_W(8, 256) <= 1; flappy_W(8, 257) <= 1; flappy_W(8, 258) <= 0; flappy_W(8, 259) <= 0; flappy_W(8, 260) <= 0; flappy_W(8, 261) <= 0; flappy_W(8, 262) <= 0; flappy_W(8, 263) <= 0; flappy_W(8, 264) <= 0; flappy_W(8, 265) <= 0; flappy_W(8, 266) <= 0; flappy_W(8, 267) <= 0; flappy_W(8, 268) <= 0; flappy_W(8, 269) <= 0; flappy_W(8, 270) <= 1; flappy_W(8, 271) <= 1; flappy_W(8, 272) <= 1; flappy_W(8, 273) <= 1; flappy_W(8, 274) <= 1; flappy_W(8, 275) <= 1; flappy_W(8, 276) <= 1; flappy_W(8, 277) <= 1; flappy_W(8, 278) <= 1; flappy_W(8, 279) <= 1; flappy_W(8, 280) <= 1; flappy_W(8, 281) <= 1; flappy_W(8, 282) <= 0; flappy_W(8, 283) <= 0; flappy_W(8, 284) <= 0; flappy_W(8, 285) <= 0; flappy_W(8, 286) <= 0; flappy_W(8, 287) <= 0; flappy_W(8, 288) <= 0; flappy_W(8, 289) <= 0; flappy_W(8, 290) <= 0; flappy_W(8, 291) <= 0; flappy_W(8, 292) <= 0; flappy_W(8, 293) <= 0; flappy_W(8, 294) <= 0; flappy_W(8, 295) <= 0; flappy_W(8, 296) <= 0; flappy_W(8, 297) <= 0; flappy_W(8, 298) <= 0; flappy_W(8, 299) <= 0; flappy_W(8, 300) <= 0; flappy_W(8, 301) <= 0; flappy_W(8, 302) <= 0; flappy_W(8, 303) <= 0; flappy_W(8, 304) <= 0; flappy_W(8, 305) <= 0; flappy_W(8, 306) <= 1; flappy_W(8, 307) <= 1; flappy_W(8, 308) <= 1; flappy_W(8, 309) <= 1; flappy_W(8, 310) <= 1; flappy_W(8, 311) <= 1; flappy_W(8, 312) <= 1; flappy_W(8, 313) <= 1; flappy_W(8, 314) <= 1; flappy_W(8, 315) <= 1; flappy_W(8, 316) <= 1; flappy_W(8, 317) <= 1; flappy_W(8, 318) <= 0; flappy_W(8, 319) <= 0; flappy_W(8, 320) <= 0; flappy_W(8, 321) <= 0; flappy_W(8, 322) <= 0; flappy_W(8, 323) <= 0; flappy_W(8, 324) <= 0; flappy_W(8, 325) <= 0; flappy_W(8, 326) <= 0; flappy_W(8, 327) <= 0; flappy_W(8, 328) <= 0; flappy_W(8, 329) <= 0; flappy_W(8, 330) <= 0; flappy_W(8, 331) <= 0; flappy_W(8, 332) <= 0; flappy_W(8, 333) <= 0; flappy_W(8, 334) <= 0; flappy_W(8, 335) <= 0; flappy_W(8, 336) <= 0; flappy_W(8, 337) <= 0; flappy_W(8, 338) <= 0; flappy_W(8, 339) <= 0; flappy_W(8, 340) <= 0; flappy_W(8, 341) <= 0; flappy_W(8, 342) <= 0; flappy_W(8, 343) <= 0; flappy_W(8, 344) <= 0; flappy_W(8, 345) <= 0; flappy_W(8, 346) <= 0; flappy_W(8, 347) <= 0; flappy_W(8, 348) <= 0; flappy_W(8, 349) <= 0; flappy_W(8, 350) <= 0; flappy_W(8, 351) <= 0; flappy_W(8, 352) <= 0; flappy_W(8, 353) <= 0; flappy_W(8, 354) <= 0; flappy_W(8, 355) <= 0; flappy_W(8, 356) <= 0; flappy_W(8, 357) <= 0; flappy_W(8, 358) <= 0; flappy_W(8, 359) <= 0; flappy_W(8, 360) <= 0; flappy_W(8, 361) <= 0; flappy_W(8, 362) <= 0; flappy_W(8, 363) <= 0; flappy_W(8, 364) <= 0; flappy_W(8, 365) <= 0; flappy_W(8, 366) <= 0; flappy_W(8, 367) <= 0; flappy_W(8, 368) <= 0; flappy_W(8, 369) <= 0; flappy_W(8, 370) <= 0; flappy_W(8, 371) <= 0; flappy_W(8, 372) <= 0; flappy_W(8, 373) <= 0; flappy_W(8, 374) <= 0; flappy_W(8, 375) <= 0; flappy_W(8, 376) <= 0; flappy_W(8, 377) <= 0; flappy_W(8, 378) <= 0; flappy_W(8, 379) <= 0; flappy_W(8, 380) <= 0; flappy_W(8, 381) <= 0; flappy_W(8, 382) <= 0; flappy_W(8, 383) <= 0; flappy_W(8, 384) <= 0; flappy_W(8, 385) <= 0; flappy_W(8, 386) <= 0; flappy_W(8, 387) <= 0; flappy_W(8, 388) <= 0; flappy_W(8, 389) <= 0; flappy_W(8, 390) <= 0; flappy_W(8, 391) <= 0; flappy_W(8, 392) <= 0; flappy_W(8, 393) <= 0; flappy_W(8, 394) <= 0; flappy_W(8, 395) <= 0; flappy_W(8, 396) <= 0; flappy_W(8, 397) <= 0; flappy_W(8, 398) <= 0; flappy_W(8, 399) <= 0; flappy_W(8, 400) <= 0; flappy_W(8, 401) <= 0; flappy_W(8, 402) <= 1; flappy_W(8, 403) <= 1; flappy_W(8, 404) <= 1; flappy_W(8, 405) <= 1; flappy_W(8, 406) <= 1; flappy_W(8, 407) <= 1; flappy_W(8, 408) <= 1; flappy_W(8, 409) <= 1; flappy_W(8, 410) <= 1; flappy_W(8, 411) <= 1; flappy_W(8, 412) <= 1; flappy_W(8, 413) <= 1; flappy_W(8, 414) <= 0; flappy_W(8, 415) <= 0; flappy_W(8, 416) <= 0; flappy_W(8, 417) <= 0; flappy_W(8, 418) <= 0; flappy_W(8, 419) <= 0; flappy_W(8, 420) <= 0; flappy_W(8, 421) <= 0; flappy_W(8, 422) <= 0; flappy_W(8, 423) <= 0; flappy_W(8, 424) <= 0; flappy_W(8, 425) <= 0; flappy_W(8, 426) <= 1; flappy_W(8, 427) <= 1; flappy_W(8, 428) <= 1; flappy_W(8, 429) <= 1; flappy_W(8, 430) <= 1; flappy_W(8, 431) <= 1; flappy_W(8, 432) <= 1; flappy_W(8, 433) <= 1; flappy_W(8, 434) <= 1; flappy_W(8, 435) <= 1; flappy_W(8, 436) <= 1; flappy_W(8, 437) <= 1; flappy_W(8, 438) <= 0; flappy_W(8, 439) <= 0; flappy_W(8, 440) <= 0; flappy_W(8, 441) <= 0; flappy_W(8, 442) <= 0; flappy_W(8, 443) <= 0; flappy_W(8, 444) <= 0; flappy_W(8, 445) <= 0; flappy_W(8, 446) <= 0; flappy_W(8, 447) <= 0; flappy_W(8, 448) <= 0; flappy_W(8, 449) <= 0; flappy_W(8, 450) <= 0; flappy_W(8, 451) <= 0; flappy_W(8, 452) <= 0; flappy_W(8, 453) <= 0; flappy_W(8, 454) <= 0; flappy_W(8, 455) <= 0; flappy_W(8, 456) <= 0; flappy_W(8, 457) <= 0; flappy_W(8, 458) <= 0; flappy_W(8, 459) <= 0; flappy_W(8, 460) <= 0; flappy_W(8, 461) <= 0; flappy_W(8, 462) <= 0; flappy_W(8, 463) <= 0; flappy_W(8, 464) <= 0; flappy_W(8, 465) <= 0; flappy_W(8, 466) <= 0; flappy_W(8, 467) <= 0; flappy_W(8, 468) <= 1; flappy_W(8, 469) <= 1; flappy_W(8, 470) <= 1; flappy_W(8, 471) <= 1; flappy_W(8, 472) <= 1; flappy_W(8, 473) <= 1; flappy_W(8, 474) <= 1; flappy_W(8, 475) <= 1; flappy_W(8, 476) <= 1; flappy_W(8, 477) <= 1; flappy_W(8, 478) <= 1; flappy_W(8, 479) <= 1; flappy_W(8, 480) <= 0; flappy_W(8, 481) <= 0; flappy_W(8, 482) <= 0; flappy_W(8, 483) <= 0; flappy_W(8, 484) <= 0; flappy_W(8, 485) <= 0; flappy_W(8, 486) <= 0; flappy_W(8, 487) <= 0; flappy_W(8, 488) <= 0; flappy_W(8, 489) <= 0; flappy_W(8, 490) <= 0; flappy_W(8, 491) <= 0; flappy_W(8, 492) <= 0; flappy_W(8, 493) <= 0; flappy_W(8, 494) <= 0; flappy_W(8, 495) <= 0; flappy_W(8, 496) <= 0; flappy_W(8, 497) <= 0; flappy_W(8, 498) <= 0; flappy_W(8, 499) <= 0; flappy_W(8, 500) <= 0; flappy_W(8, 501) <= 0; flappy_W(8, 502) <= 0; flappy_W(8, 503) <= 0; flappy_W(8, 504) <= 0; flappy_W(8, 505) <= 0; flappy_W(8, 506) <= 0; flappy_W(8, 507) <= 0; flappy_W(8, 508) <= 0; flappy_W(8, 509) <= 0; flappy_W(8, 510) <= 1; flappy_W(8, 511) <= 1; flappy_W(8, 512) <= 1; flappy_W(8, 513) <= 1; flappy_W(8, 514) <= 1; flappy_W(8, 515) <= 1; flappy_W(8, 516) <= 1; flappy_W(8, 517) <= 1; flappy_W(8, 518) <= 1; flappy_W(8, 519) <= 1; flappy_W(8, 520) <= 1; flappy_W(8, 521) <= 1; flappy_W(8, 522) <= 0; flappy_W(8, 523) <= 0; flappy_W(8, 524) <= 0; flappy_W(8, 525) <= 0; flappy_W(8, 526) <= 0; flappy_W(8, 527) <= 0; flappy_W(8, 528) <= 0; flappy_W(8, 529) <= 0; flappy_W(8, 530) <= 0; flappy_W(8, 531) <= 0; flappy_W(8, 532) <= 0; flappy_W(8, 533) <= 0; flappy_W(8, 534) <= 1; flappy_W(8, 535) <= 1; flappy_W(8, 536) <= 1; flappy_W(8, 537) <= 1; flappy_W(8, 538) <= 1; flappy_W(8, 539) <= 1; flappy_W(8, 540) <= 1; flappy_W(8, 541) <= 1; flappy_W(8, 542) <= 1; flappy_W(8, 543) <= 1; flappy_W(8, 544) <= 1; flappy_W(8, 545) <= 1; flappy_W(8, 546) <= 0; flappy_W(8, 547) <= 0; flappy_W(8, 548) <= 0; flappy_W(8, 549) <= 0; flappy_W(8, 550) <= 0; flappy_W(8, 551) <= 0; flappy_W(8, 552) <= 0; flappy_W(8, 553) <= 0; flappy_W(8, 554) <= 0; flappy_W(8, 555) <= 0; flappy_W(8, 556) <= 0; flappy_W(8, 557) <= 0; flappy_W(8, 558) <= 0; flappy_W(8, 559) <= 0; flappy_W(8, 560) <= 0; flappy_W(8, 561) <= 0; flappy_W(8, 562) <= 0; flappy_W(8, 563) <= 0; flappy_W(8, 564) <= 1; flappy_W(8, 565) <= 1; flappy_W(8, 566) <= 1; flappy_W(8, 567) <= 1; flappy_W(8, 568) <= 1; flappy_W(8, 569) <= 1; flappy_W(8, 570) <= 1; flappy_W(8, 571) <= 1; flappy_W(8, 572) <= 1; flappy_W(8, 573) <= 1; flappy_W(8, 574) <= 1; flappy_W(8, 575) <= 1; flappy_W(8, 576) <= 0; flappy_W(8, 577) <= 0; flappy_W(8, 578) <= 0; flappy_W(8, 579) <= 0; flappy_W(8, 580) <= 0; flappy_W(8, 581) <= 0; flappy_W(8, 582) <= 1; flappy_W(8, 583) <= 1; flappy_W(8, 584) <= 1; flappy_W(8, 585) <= 1; flappy_W(8, 586) <= 1; flappy_W(8, 587) <= 1; flappy_W(8, 588) <= 1; flappy_W(8, 589) <= 1; flappy_W(8, 590) <= 1; flappy_W(8, 591) <= 1; flappy_W(8, 592) <= 1; flappy_W(8, 593) <= 1; 
flappy_W(9, 0) <= 0; flappy_W(9, 1) <= 0; flappy_W(9, 2) <= 0; flappy_W(9, 3) <= 0; flappy_W(9, 4) <= 0; flappy_W(9, 5) <= 0; flappy_W(9, 6) <= 1; flappy_W(9, 7) <= 1; flappy_W(9, 8) <= 1; flappy_W(9, 9) <= 1; flappy_W(9, 10) <= 1; flappy_W(9, 11) <= 1; flappy_W(9, 12) <= 1; flappy_W(9, 13) <= 1; flappy_W(9, 14) <= 1; flappy_W(9, 15) <= 1; flappy_W(9, 16) <= 1; flappy_W(9, 17) <= 1; flappy_W(9, 18) <= 0; flappy_W(9, 19) <= 0; flappy_W(9, 20) <= 0; flappy_W(9, 21) <= 0; flappy_W(9, 22) <= 0; flappy_W(9, 23) <= 0; flappy_W(9, 24) <= 0; flappy_W(9, 25) <= 0; flappy_W(9, 26) <= 0; flappy_W(9, 27) <= 0; flappy_W(9, 28) <= 0; flappy_W(9, 29) <= 0; flappy_W(9, 30) <= 1; flappy_W(9, 31) <= 1; flappy_W(9, 32) <= 1; flappy_W(9, 33) <= 1; flappy_W(9, 34) <= 1; flappy_W(9, 35) <= 1; flappy_W(9, 36) <= 1; flappy_W(9, 37) <= 1; flappy_W(9, 38) <= 1; flappy_W(9, 39) <= 1; flappy_W(9, 40) <= 1; flappy_W(9, 41) <= 1; flappy_W(9, 42) <= 0; flappy_W(9, 43) <= 0; flappy_W(9, 44) <= 0; flappy_W(9, 45) <= 0; flappy_W(9, 46) <= 0; flappy_W(9, 47) <= 0; flappy_W(9, 48) <= 0; flappy_W(9, 49) <= 0; flappy_W(9, 50) <= 0; flappy_W(9, 51) <= 0; flappy_W(9, 52) <= 0; flappy_W(9, 53) <= 0; flappy_W(9, 54) <= 0; flappy_W(9, 55) <= 0; flappy_W(9, 56) <= 0; flappy_W(9, 57) <= 0; flappy_W(9, 58) <= 0; flappy_W(9, 59) <= 0; flappy_W(9, 60) <= 1; flappy_W(9, 61) <= 1; flappy_W(9, 62) <= 1; flappy_W(9, 63) <= 1; flappy_W(9, 64) <= 1; flappy_W(9, 65) <= 1; flappy_W(9, 66) <= 1; flappy_W(9, 67) <= 1; flappy_W(9, 68) <= 1; flappy_W(9, 69) <= 1; flappy_W(9, 70) <= 1; flappy_W(9, 71) <= 1; flappy_W(9, 72) <= 0; flappy_W(9, 73) <= 0; flappy_W(9, 74) <= 0; flappy_W(9, 75) <= 0; flappy_W(9, 76) <= 0; flappy_W(9, 77) <= 0; flappy_W(9, 78) <= 0; flappy_W(9, 79) <= 0; flappy_W(9, 80) <= 0; flappy_W(9, 81) <= 0; flappy_W(9, 82) <= 0; flappy_W(9, 83) <= 0; flappy_W(9, 84) <= 0; flappy_W(9, 85) <= 0; flappy_W(9, 86) <= 0; flappy_W(9, 87) <= 0; flappy_W(9, 88) <= 0; flappy_W(9, 89) <= 0; flappy_W(9, 90) <= 0; flappy_W(9, 91) <= 0; flappy_W(9, 92) <= 0; flappy_W(9, 93) <= 0; flappy_W(9, 94) <= 0; flappy_W(9, 95) <= 0; flappy_W(9, 96) <= 0; flappy_W(9, 97) <= 0; flappy_W(9, 98) <= 0; flappy_W(9, 99) <= 0; flappy_W(9, 100) <= 0; flappy_W(9, 101) <= 0; flappy_W(9, 102) <= 0; flappy_W(9, 103) <= 0; flappy_W(9, 104) <= 0; flappy_W(9, 105) <= 0; flappy_W(9, 106) <= 0; flappy_W(9, 107) <= 0; flappy_W(9, 108) <= 0; flappy_W(9, 109) <= 0; flappy_W(9, 110) <= 0; flappy_W(9, 111) <= 0; flappy_W(9, 112) <= 0; flappy_W(9, 113) <= 0; flappy_W(9, 114) <= 0; flappy_W(9, 115) <= 0; flappy_W(9, 116) <= 0; flappy_W(9, 117) <= 0; flappy_W(9, 118) <= 0; flappy_W(9, 119) <= 0; flappy_W(9, 120) <= 1; flappy_W(9, 121) <= 1; flappy_W(9, 122) <= 1; flappy_W(9, 123) <= 1; flappy_W(9, 124) <= 1; flappy_W(9, 125) <= 1; flappy_W(9, 126) <= 1; flappy_W(9, 127) <= 1; flappy_W(9, 128) <= 1; flappy_W(9, 129) <= 1; flappy_W(9, 130) <= 1; flappy_W(9, 131) <= 1; flappy_W(9, 132) <= 1; flappy_W(9, 133) <= 1; flappy_W(9, 134) <= 1; flappy_W(9, 135) <= 1; flappy_W(9, 136) <= 1; flappy_W(9, 137) <= 1; flappy_W(9, 138) <= 0; flappy_W(9, 139) <= 0; flappy_W(9, 140) <= 0; flappy_W(9, 141) <= 0; flappy_W(9, 142) <= 0; flappy_W(9, 143) <= 0; flappy_W(9, 144) <= 0; flappy_W(9, 145) <= 0; flappy_W(9, 146) <= 0; flappy_W(9, 147) <= 0; flappy_W(9, 148) <= 0; flappy_W(9, 149) <= 0; flappy_W(9, 150) <= 0; flappy_W(9, 151) <= 0; flappy_W(9, 152) <= 0; flappy_W(9, 153) <= 0; flappy_W(9, 154) <= 0; flappy_W(9, 155) <= 0; flappy_W(9, 156) <= 0; flappy_W(9, 157) <= 0; flappy_W(9, 158) <= 0; flappy_W(9, 159) <= 0; flappy_W(9, 160) <= 0; flappy_W(9, 161) <= 0; flappy_W(9, 162) <= 0; flappy_W(9, 163) <= 0; flappy_W(9, 164) <= 0; flappy_W(9, 165) <= 0; flappy_W(9, 166) <= 0; flappy_W(9, 167) <= 0; flappy_W(9, 168) <= 1; flappy_W(9, 169) <= 1; flappy_W(9, 170) <= 1; flappy_W(9, 171) <= 1; flappy_W(9, 172) <= 1; flappy_W(9, 173) <= 1; flappy_W(9, 174) <= 1; flappy_W(9, 175) <= 1; flappy_W(9, 176) <= 1; flappy_W(9, 177) <= 1; flappy_W(9, 178) <= 1; flappy_W(9, 179) <= 1; flappy_W(9, 180) <= 0; flappy_W(9, 181) <= 0; flappy_W(9, 182) <= 0; flappy_W(9, 183) <= 0; flappy_W(9, 184) <= 0; flappy_W(9, 185) <= 0; flappy_W(9, 186) <= 0; flappy_W(9, 187) <= 0; flappy_W(9, 188) <= 0; flappy_W(9, 189) <= 0; flappy_W(9, 190) <= 0; flappy_W(9, 191) <= 0; flappy_W(9, 192) <= 1; flappy_W(9, 193) <= 1; flappy_W(9, 194) <= 1; flappy_W(9, 195) <= 1; flappy_W(9, 196) <= 1; flappy_W(9, 197) <= 1; flappy_W(9, 198) <= 1; flappy_W(9, 199) <= 1; flappy_W(9, 200) <= 1; flappy_W(9, 201) <= 1; flappy_W(9, 202) <= 1; flappy_W(9, 203) <= 1; flappy_W(9, 204) <= 0; flappy_W(9, 205) <= 0; flappy_W(9, 206) <= 0; flappy_W(9, 207) <= 0; flappy_W(9, 208) <= 0; flappy_W(9, 209) <= 0; flappy_W(9, 210) <= 0; flappy_W(9, 211) <= 0; flappy_W(9, 212) <= 0; flappy_W(9, 213) <= 0; flappy_W(9, 214) <= 0; flappy_W(9, 215) <= 0; flappy_W(9, 216) <= 0; flappy_W(9, 217) <= 0; flappy_W(9, 218) <= 0; flappy_W(9, 219) <= 0; flappy_W(9, 220) <= 0; flappy_W(9, 221) <= 0; flappy_W(9, 222) <= 1; flappy_W(9, 223) <= 1; flappy_W(9, 224) <= 1; flappy_W(9, 225) <= 1; flappy_W(9, 226) <= 1; flappy_W(9, 227) <= 1; flappy_W(9, 228) <= 1; flappy_W(9, 229) <= 1; flappy_W(9, 230) <= 1; flappy_W(9, 231) <= 1; flappy_W(9, 232) <= 1; flappy_W(9, 233) <= 1; flappy_W(9, 234) <= 0; flappy_W(9, 235) <= 0; flappy_W(9, 236) <= 0; flappy_W(9, 237) <= 0; flappy_W(9, 238) <= 0; flappy_W(9, 239) <= 0; flappy_W(9, 240) <= 0; flappy_W(9, 241) <= 0; flappy_W(9, 242) <= 0; flappy_W(9, 243) <= 0; flappy_W(9, 244) <= 0; flappy_W(9, 245) <= 0; flappy_W(9, 246) <= 1; flappy_W(9, 247) <= 1; flappy_W(9, 248) <= 1; flappy_W(9, 249) <= 1; flappy_W(9, 250) <= 1; flappy_W(9, 251) <= 1; flappy_W(9, 252) <= 1; flappy_W(9, 253) <= 1; flappy_W(9, 254) <= 1; flappy_W(9, 255) <= 1; flappy_W(9, 256) <= 1; flappy_W(9, 257) <= 1; flappy_W(9, 258) <= 0; flappy_W(9, 259) <= 0; flappy_W(9, 260) <= 0; flappy_W(9, 261) <= 0; flappy_W(9, 262) <= 0; flappy_W(9, 263) <= 0; flappy_W(9, 264) <= 0; flappy_W(9, 265) <= 0; flappy_W(9, 266) <= 0; flappy_W(9, 267) <= 0; flappy_W(9, 268) <= 0; flappy_W(9, 269) <= 0; flappy_W(9, 270) <= 1; flappy_W(9, 271) <= 1; flappy_W(9, 272) <= 1; flappy_W(9, 273) <= 1; flappy_W(9, 274) <= 1; flappy_W(9, 275) <= 1; flappy_W(9, 276) <= 1; flappy_W(9, 277) <= 1; flappy_W(9, 278) <= 1; flappy_W(9, 279) <= 1; flappy_W(9, 280) <= 1; flappy_W(9, 281) <= 1; flappy_W(9, 282) <= 0; flappy_W(9, 283) <= 0; flappy_W(9, 284) <= 0; flappy_W(9, 285) <= 0; flappy_W(9, 286) <= 0; flappy_W(9, 287) <= 0; flappy_W(9, 288) <= 0; flappy_W(9, 289) <= 0; flappy_W(9, 290) <= 0; flappy_W(9, 291) <= 0; flappy_W(9, 292) <= 0; flappy_W(9, 293) <= 0; flappy_W(9, 294) <= 0; flappy_W(9, 295) <= 0; flappy_W(9, 296) <= 0; flappy_W(9, 297) <= 0; flappy_W(9, 298) <= 0; flappy_W(9, 299) <= 0; flappy_W(9, 300) <= 0; flappy_W(9, 301) <= 0; flappy_W(9, 302) <= 0; flappy_W(9, 303) <= 0; flappy_W(9, 304) <= 0; flappy_W(9, 305) <= 0; flappy_W(9, 306) <= 1; flappy_W(9, 307) <= 1; flappy_W(9, 308) <= 1; flappy_W(9, 309) <= 1; flappy_W(9, 310) <= 1; flappy_W(9, 311) <= 1; flappy_W(9, 312) <= 1; flappy_W(9, 313) <= 1; flappy_W(9, 314) <= 1; flappy_W(9, 315) <= 1; flappy_W(9, 316) <= 1; flappy_W(9, 317) <= 1; flappy_W(9, 318) <= 0; flappy_W(9, 319) <= 0; flappy_W(9, 320) <= 0; flappy_W(9, 321) <= 0; flappy_W(9, 322) <= 0; flappy_W(9, 323) <= 0; flappy_W(9, 324) <= 0; flappy_W(9, 325) <= 0; flappy_W(9, 326) <= 0; flappy_W(9, 327) <= 0; flappy_W(9, 328) <= 0; flappy_W(9, 329) <= 0; flappy_W(9, 330) <= 0; flappy_W(9, 331) <= 0; flappy_W(9, 332) <= 0; flappy_W(9, 333) <= 0; flappy_W(9, 334) <= 0; flappy_W(9, 335) <= 0; flappy_W(9, 336) <= 0; flappy_W(9, 337) <= 0; flappy_W(9, 338) <= 0; flappy_W(9, 339) <= 0; flappy_W(9, 340) <= 0; flappy_W(9, 341) <= 0; flappy_W(9, 342) <= 0; flappy_W(9, 343) <= 0; flappy_W(9, 344) <= 0; flappy_W(9, 345) <= 0; flappy_W(9, 346) <= 0; flappy_W(9, 347) <= 0; flappy_W(9, 348) <= 0; flappy_W(9, 349) <= 0; flappy_W(9, 350) <= 0; flappy_W(9, 351) <= 0; flappy_W(9, 352) <= 0; flappy_W(9, 353) <= 0; flappy_W(9, 354) <= 0; flappy_W(9, 355) <= 0; flappy_W(9, 356) <= 0; flappy_W(9, 357) <= 0; flappy_W(9, 358) <= 0; flappy_W(9, 359) <= 0; flappy_W(9, 360) <= 0; flappy_W(9, 361) <= 0; flappy_W(9, 362) <= 0; flappy_W(9, 363) <= 0; flappy_W(9, 364) <= 0; flappy_W(9, 365) <= 0; flappy_W(9, 366) <= 0; flappy_W(9, 367) <= 0; flappy_W(9, 368) <= 0; flappy_W(9, 369) <= 0; flappy_W(9, 370) <= 0; flappy_W(9, 371) <= 0; flappy_W(9, 372) <= 0; flappy_W(9, 373) <= 0; flappy_W(9, 374) <= 0; flappy_W(9, 375) <= 0; flappy_W(9, 376) <= 0; flappy_W(9, 377) <= 0; flappy_W(9, 378) <= 0; flappy_W(9, 379) <= 0; flappy_W(9, 380) <= 0; flappy_W(9, 381) <= 0; flappy_W(9, 382) <= 0; flappy_W(9, 383) <= 0; flappy_W(9, 384) <= 0; flappy_W(9, 385) <= 0; flappy_W(9, 386) <= 0; flappy_W(9, 387) <= 0; flappy_W(9, 388) <= 0; flappy_W(9, 389) <= 0; flappy_W(9, 390) <= 0; flappy_W(9, 391) <= 0; flappy_W(9, 392) <= 0; flappy_W(9, 393) <= 0; flappy_W(9, 394) <= 0; flappy_W(9, 395) <= 0; flappy_W(9, 396) <= 0; flappy_W(9, 397) <= 0; flappy_W(9, 398) <= 0; flappy_W(9, 399) <= 0; flappy_W(9, 400) <= 0; flappy_W(9, 401) <= 0; flappy_W(9, 402) <= 1; flappy_W(9, 403) <= 1; flappy_W(9, 404) <= 1; flappy_W(9, 405) <= 1; flappy_W(9, 406) <= 1; flappy_W(9, 407) <= 1; flappy_W(9, 408) <= 1; flappy_W(9, 409) <= 1; flappy_W(9, 410) <= 1; flappy_W(9, 411) <= 1; flappy_W(9, 412) <= 1; flappy_W(9, 413) <= 1; flappy_W(9, 414) <= 0; flappy_W(9, 415) <= 0; flappy_W(9, 416) <= 0; flappy_W(9, 417) <= 0; flappy_W(9, 418) <= 0; flappy_W(9, 419) <= 0; flappy_W(9, 420) <= 0; flappy_W(9, 421) <= 0; flappy_W(9, 422) <= 0; flappy_W(9, 423) <= 0; flappy_W(9, 424) <= 0; flappy_W(9, 425) <= 0; flappy_W(9, 426) <= 1; flappy_W(9, 427) <= 1; flappy_W(9, 428) <= 1; flappy_W(9, 429) <= 1; flappy_W(9, 430) <= 1; flappy_W(9, 431) <= 1; flappy_W(9, 432) <= 1; flappy_W(9, 433) <= 1; flappy_W(9, 434) <= 1; flappy_W(9, 435) <= 1; flappy_W(9, 436) <= 1; flappy_W(9, 437) <= 1; flappy_W(9, 438) <= 0; flappy_W(9, 439) <= 0; flappy_W(9, 440) <= 0; flappy_W(9, 441) <= 0; flappy_W(9, 442) <= 0; flappy_W(9, 443) <= 0; flappy_W(9, 444) <= 0; flappy_W(9, 445) <= 0; flappy_W(9, 446) <= 0; flappy_W(9, 447) <= 0; flappy_W(9, 448) <= 0; flappy_W(9, 449) <= 0; flappy_W(9, 450) <= 0; flappy_W(9, 451) <= 0; flappy_W(9, 452) <= 0; flappy_W(9, 453) <= 0; flappy_W(9, 454) <= 0; flappy_W(9, 455) <= 0; flappy_W(9, 456) <= 0; flappy_W(9, 457) <= 0; flappy_W(9, 458) <= 0; flappy_W(9, 459) <= 0; flappy_W(9, 460) <= 0; flappy_W(9, 461) <= 0; flappy_W(9, 462) <= 0; flappy_W(9, 463) <= 0; flappy_W(9, 464) <= 0; flappy_W(9, 465) <= 0; flappy_W(9, 466) <= 0; flappy_W(9, 467) <= 0; flappy_W(9, 468) <= 1; flappy_W(9, 469) <= 1; flappy_W(9, 470) <= 1; flappy_W(9, 471) <= 1; flappy_W(9, 472) <= 1; flappy_W(9, 473) <= 1; flappy_W(9, 474) <= 1; flappy_W(9, 475) <= 1; flappy_W(9, 476) <= 1; flappy_W(9, 477) <= 1; flappy_W(9, 478) <= 1; flappy_W(9, 479) <= 1; flappy_W(9, 480) <= 0; flappy_W(9, 481) <= 0; flappy_W(9, 482) <= 0; flappy_W(9, 483) <= 0; flappy_W(9, 484) <= 0; flappy_W(9, 485) <= 0; flappy_W(9, 486) <= 0; flappy_W(9, 487) <= 0; flappy_W(9, 488) <= 0; flappy_W(9, 489) <= 0; flappy_W(9, 490) <= 0; flappy_W(9, 491) <= 0; flappy_W(9, 492) <= 0; flappy_W(9, 493) <= 0; flappy_W(9, 494) <= 0; flappy_W(9, 495) <= 0; flappy_W(9, 496) <= 0; flappy_W(9, 497) <= 0; flappy_W(9, 498) <= 0; flappy_W(9, 499) <= 0; flappy_W(9, 500) <= 0; flappy_W(9, 501) <= 0; flappy_W(9, 502) <= 0; flappy_W(9, 503) <= 0; flappy_W(9, 504) <= 0; flappy_W(9, 505) <= 0; flappy_W(9, 506) <= 0; flappy_W(9, 507) <= 0; flappy_W(9, 508) <= 0; flappy_W(9, 509) <= 0; flappy_W(9, 510) <= 1; flappy_W(9, 511) <= 1; flappy_W(9, 512) <= 1; flappy_W(9, 513) <= 1; flappy_W(9, 514) <= 1; flappy_W(9, 515) <= 1; flappy_W(9, 516) <= 1; flappy_W(9, 517) <= 1; flappy_W(9, 518) <= 1; flappy_W(9, 519) <= 1; flappy_W(9, 520) <= 1; flappy_W(9, 521) <= 1; flappy_W(9, 522) <= 0; flappy_W(9, 523) <= 0; flappy_W(9, 524) <= 0; flappy_W(9, 525) <= 0; flappy_W(9, 526) <= 0; flappy_W(9, 527) <= 0; flappy_W(9, 528) <= 0; flappy_W(9, 529) <= 0; flappy_W(9, 530) <= 0; flappy_W(9, 531) <= 0; flappy_W(9, 532) <= 0; flappy_W(9, 533) <= 0; flappy_W(9, 534) <= 1; flappy_W(9, 535) <= 1; flappy_W(9, 536) <= 1; flappy_W(9, 537) <= 1; flappy_W(9, 538) <= 1; flappy_W(9, 539) <= 1; flappy_W(9, 540) <= 1; flappy_W(9, 541) <= 1; flappy_W(9, 542) <= 1; flappy_W(9, 543) <= 1; flappy_W(9, 544) <= 1; flappy_W(9, 545) <= 1; flappy_W(9, 546) <= 0; flappy_W(9, 547) <= 0; flappy_W(9, 548) <= 0; flappy_W(9, 549) <= 0; flappy_W(9, 550) <= 0; flappy_W(9, 551) <= 0; flappy_W(9, 552) <= 0; flappy_W(9, 553) <= 0; flappy_W(9, 554) <= 0; flappy_W(9, 555) <= 0; flappy_W(9, 556) <= 0; flappy_W(9, 557) <= 0; flappy_W(9, 558) <= 0; flappy_W(9, 559) <= 0; flappy_W(9, 560) <= 0; flappy_W(9, 561) <= 0; flappy_W(9, 562) <= 0; flappy_W(9, 563) <= 0; flappy_W(9, 564) <= 1; flappy_W(9, 565) <= 1; flappy_W(9, 566) <= 1; flappy_W(9, 567) <= 1; flappy_W(9, 568) <= 1; flappy_W(9, 569) <= 1; flappy_W(9, 570) <= 1; flappy_W(9, 571) <= 1; flappy_W(9, 572) <= 1; flappy_W(9, 573) <= 1; flappy_W(9, 574) <= 1; flappy_W(9, 575) <= 1; flappy_W(9, 576) <= 0; flappy_W(9, 577) <= 0; flappy_W(9, 578) <= 0; flappy_W(9, 579) <= 0; flappy_W(9, 580) <= 0; flappy_W(9, 581) <= 0; flappy_W(9, 582) <= 1; flappy_W(9, 583) <= 1; flappy_W(9, 584) <= 1; flappy_W(9, 585) <= 1; flappy_W(9, 586) <= 1; flappy_W(9, 587) <= 1; flappy_W(9, 588) <= 1; flappy_W(9, 589) <= 1; flappy_W(9, 590) <= 1; flappy_W(9, 591) <= 1; flappy_W(9, 592) <= 1; flappy_W(9, 593) <= 1; 
flappy_W(10, 0) <= 0; flappy_W(10, 1) <= 0; flappy_W(10, 2) <= 0; flappy_W(10, 3) <= 0; flappy_W(10, 4) <= 0; flappy_W(10, 5) <= 0; flappy_W(10, 6) <= 1; flappy_W(10, 7) <= 1; flappy_W(10, 8) <= 1; flappy_W(10, 9) <= 1; flappy_W(10, 10) <= 1; flappy_W(10, 11) <= 1; flappy_W(10, 12) <= 1; flappy_W(10, 13) <= 1; flappy_W(10, 14) <= 1; flappy_W(10, 15) <= 1; flappy_W(10, 16) <= 1; flappy_W(10, 17) <= 1; flappy_W(10, 18) <= 0; flappy_W(10, 19) <= 0; flappy_W(10, 20) <= 0; flappy_W(10, 21) <= 0; flappy_W(10, 22) <= 0; flappy_W(10, 23) <= 0; flappy_W(10, 24) <= 0; flappy_W(10, 25) <= 0; flappy_W(10, 26) <= 0; flappy_W(10, 27) <= 0; flappy_W(10, 28) <= 0; flappy_W(10, 29) <= 0; flappy_W(10, 30) <= 1; flappy_W(10, 31) <= 1; flappy_W(10, 32) <= 1; flappy_W(10, 33) <= 1; flappy_W(10, 34) <= 1; flappy_W(10, 35) <= 1; flappy_W(10, 36) <= 1; flappy_W(10, 37) <= 1; flappy_W(10, 38) <= 1; flappy_W(10, 39) <= 1; flappy_W(10, 40) <= 1; flappy_W(10, 41) <= 1; flappy_W(10, 42) <= 0; flappy_W(10, 43) <= 0; flappy_W(10, 44) <= 0; flappy_W(10, 45) <= 0; flappy_W(10, 46) <= 0; flappy_W(10, 47) <= 0; flappy_W(10, 48) <= 0; flappy_W(10, 49) <= 0; flappy_W(10, 50) <= 0; flappy_W(10, 51) <= 0; flappy_W(10, 52) <= 0; flappy_W(10, 53) <= 0; flappy_W(10, 54) <= 0; flappy_W(10, 55) <= 0; flappy_W(10, 56) <= 0; flappy_W(10, 57) <= 0; flappy_W(10, 58) <= 0; flappy_W(10, 59) <= 0; flappy_W(10, 60) <= 1; flappy_W(10, 61) <= 1; flappy_W(10, 62) <= 1; flappy_W(10, 63) <= 1; flappy_W(10, 64) <= 1; flappy_W(10, 65) <= 1; flappy_W(10, 66) <= 1; flappy_W(10, 67) <= 1; flappy_W(10, 68) <= 1; flappy_W(10, 69) <= 1; flappy_W(10, 70) <= 1; flappy_W(10, 71) <= 1; flappy_W(10, 72) <= 0; flappy_W(10, 73) <= 0; flappy_W(10, 74) <= 0; flappy_W(10, 75) <= 0; flappy_W(10, 76) <= 0; flappy_W(10, 77) <= 0; flappy_W(10, 78) <= 0; flappy_W(10, 79) <= 0; flappy_W(10, 80) <= 0; flappy_W(10, 81) <= 0; flappy_W(10, 82) <= 0; flappy_W(10, 83) <= 0; flappy_W(10, 84) <= 0; flappy_W(10, 85) <= 0; flappy_W(10, 86) <= 0; flappy_W(10, 87) <= 0; flappy_W(10, 88) <= 0; flappy_W(10, 89) <= 0; flappy_W(10, 90) <= 0; flappy_W(10, 91) <= 0; flappy_W(10, 92) <= 0; flappy_W(10, 93) <= 0; flappy_W(10, 94) <= 0; flappy_W(10, 95) <= 0; flappy_W(10, 96) <= 0; flappy_W(10, 97) <= 0; flappy_W(10, 98) <= 0; flappy_W(10, 99) <= 0; flappy_W(10, 100) <= 0; flappy_W(10, 101) <= 0; flappy_W(10, 102) <= 0; flappy_W(10, 103) <= 0; flappy_W(10, 104) <= 0; flappy_W(10, 105) <= 0; flappy_W(10, 106) <= 0; flappy_W(10, 107) <= 0; flappy_W(10, 108) <= 0; flappy_W(10, 109) <= 0; flappy_W(10, 110) <= 0; flappy_W(10, 111) <= 0; flappy_W(10, 112) <= 0; flappy_W(10, 113) <= 0; flappy_W(10, 114) <= 0; flappy_W(10, 115) <= 0; flappy_W(10, 116) <= 0; flappy_W(10, 117) <= 0; flappy_W(10, 118) <= 0; flappy_W(10, 119) <= 0; flappy_W(10, 120) <= 1; flappy_W(10, 121) <= 1; flappy_W(10, 122) <= 1; flappy_W(10, 123) <= 1; flappy_W(10, 124) <= 1; flappy_W(10, 125) <= 1; flappy_W(10, 126) <= 1; flappy_W(10, 127) <= 1; flappy_W(10, 128) <= 1; flappy_W(10, 129) <= 1; flappy_W(10, 130) <= 1; flappy_W(10, 131) <= 1; flappy_W(10, 132) <= 1; flappy_W(10, 133) <= 1; flappy_W(10, 134) <= 1; flappy_W(10, 135) <= 1; flappy_W(10, 136) <= 1; flappy_W(10, 137) <= 1; flappy_W(10, 138) <= 0; flappy_W(10, 139) <= 0; flappy_W(10, 140) <= 0; flappy_W(10, 141) <= 0; flappy_W(10, 142) <= 0; flappy_W(10, 143) <= 0; flappy_W(10, 144) <= 0; flappy_W(10, 145) <= 0; flappy_W(10, 146) <= 0; flappy_W(10, 147) <= 0; flappy_W(10, 148) <= 0; flappy_W(10, 149) <= 0; flappy_W(10, 150) <= 0; flappy_W(10, 151) <= 0; flappy_W(10, 152) <= 0; flappy_W(10, 153) <= 0; flappy_W(10, 154) <= 0; flappy_W(10, 155) <= 0; flappy_W(10, 156) <= 0; flappy_W(10, 157) <= 0; flappy_W(10, 158) <= 0; flappy_W(10, 159) <= 0; flappy_W(10, 160) <= 0; flappy_W(10, 161) <= 0; flappy_W(10, 162) <= 0; flappy_W(10, 163) <= 0; flappy_W(10, 164) <= 0; flappy_W(10, 165) <= 0; flappy_W(10, 166) <= 0; flappy_W(10, 167) <= 0; flappy_W(10, 168) <= 1; flappy_W(10, 169) <= 1; flappy_W(10, 170) <= 1; flappy_W(10, 171) <= 1; flappy_W(10, 172) <= 1; flappy_W(10, 173) <= 1; flappy_W(10, 174) <= 1; flappy_W(10, 175) <= 1; flappy_W(10, 176) <= 1; flappy_W(10, 177) <= 1; flappy_W(10, 178) <= 1; flappy_W(10, 179) <= 1; flappy_W(10, 180) <= 0; flappy_W(10, 181) <= 0; flappy_W(10, 182) <= 0; flappy_W(10, 183) <= 0; flappy_W(10, 184) <= 0; flappy_W(10, 185) <= 0; flappy_W(10, 186) <= 0; flappy_W(10, 187) <= 0; flappy_W(10, 188) <= 0; flappy_W(10, 189) <= 0; flappy_W(10, 190) <= 0; flappy_W(10, 191) <= 0; flappy_W(10, 192) <= 1; flappy_W(10, 193) <= 1; flappy_W(10, 194) <= 1; flappy_W(10, 195) <= 1; flappy_W(10, 196) <= 1; flappy_W(10, 197) <= 1; flappy_W(10, 198) <= 1; flappy_W(10, 199) <= 1; flappy_W(10, 200) <= 1; flappy_W(10, 201) <= 1; flappy_W(10, 202) <= 1; flappy_W(10, 203) <= 1; flappy_W(10, 204) <= 0; flappy_W(10, 205) <= 0; flappy_W(10, 206) <= 0; flappy_W(10, 207) <= 0; flappy_W(10, 208) <= 0; flappy_W(10, 209) <= 0; flappy_W(10, 210) <= 0; flappy_W(10, 211) <= 0; flappy_W(10, 212) <= 0; flappy_W(10, 213) <= 0; flappy_W(10, 214) <= 0; flappy_W(10, 215) <= 0; flappy_W(10, 216) <= 0; flappy_W(10, 217) <= 0; flappy_W(10, 218) <= 0; flappy_W(10, 219) <= 0; flappy_W(10, 220) <= 0; flappy_W(10, 221) <= 0; flappy_W(10, 222) <= 1; flappy_W(10, 223) <= 1; flappy_W(10, 224) <= 1; flappy_W(10, 225) <= 1; flappy_W(10, 226) <= 1; flappy_W(10, 227) <= 1; flappy_W(10, 228) <= 1; flappy_W(10, 229) <= 1; flappy_W(10, 230) <= 1; flappy_W(10, 231) <= 1; flappy_W(10, 232) <= 1; flappy_W(10, 233) <= 1; flappy_W(10, 234) <= 0; flappy_W(10, 235) <= 0; flappy_W(10, 236) <= 0; flappy_W(10, 237) <= 0; flappy_W(10, 238) <= 0; flappy_W(10, 239) <= 0; flappy_W(10, 240) <= 0; flappy_W(10, 241) <= 0; flappy_W(10, 242) <= 0; flappy_W(10, 243) <= 0; flappy_W(10, 244) <= 0; flappy_W(10, 245) <= 0; flappy_W(10, 246) <= 1; flappy_W(10, 247) <= 1; flappy_W(10, 248) <= 1; flappy_W(10, 249) <= 1; flappy_W(10, 250) <= 1; flappy_W(10, 251) <= 1; flappy_W(10, 252) <= 1; flappy_W(10, 253) <= 1; flappy_W(10, 254) <= 1; flappy_W(10, 255) <= 1; flappy_W(10, 256) <= 1; flappy_W(10, 257) <= 1; flappy_W(10, 258) <= 0; flappy_W(10, 259) <= 0; flappy_W(10, 260) <= 0; flappy_W(10, 261) <= 0; flappy_W(10, 262) <= 0; flappy_W(10, 263) <= 0; flappy_W(10, 264) <= 0; flappy_W(10, 265) <= 0; flappy_W(10, 266) <= 0; flappy_W(10, 267) <= 0; flappy_W(10, 268) <= 0; flappy_W(10, 269) <= 0; flappy_W(10, 270) <= 1; flappy_W(10, 271) <= 1; flappy_W(10, 272) <= 1; flappy_W(10, 273) <= 1; flappy_W(10, 274) <= 1; flappy_W(10, 275) <= 1; flappy_W(10, 276) <= 1; flappy_W(10, 277) <= 1; flappy_W(10, 278) <= 1; flappy_W(10, 279) <= 1; flappy_W(10, 280) <= 1; flappy_W(10, 281) <= 1; flappy_W(10, 282) <= 0; flappy_W(10, 283) <= 0; flappy_W(10, 284) <= 0; flappy_W(10, 285) <= 0; flappy_W(10, 286) <= 0; flappy_W(10, 287) <= 0; flappy_W(10, 288) <= 0; flappy_W(10, 289) <= 0; flappy_W(10, 290) <= 0; flappy_W(10, 291) <= 0; flappy_W(10, 292) <= 0; flappy_W(10, 293) <= 0; flappy_W(10, 294) <= 0; flappy_W(10, 295) <= 0; flappy_W(10, 296) <= 0; flappy_W(10, 297) <= 0; flappy_W(10, 298) <= 0; flappy_W(10, 299) <= 0; flappy_W(10, 300) <= 0; flappy_W(10, 301) <= 0; flappy_W(10, 302) <= 0; flappy_W(10, 303) <= 0; flappy_W(10, 304) <= 0; flappy_W(10, 305) <= 0; flappy_W(10, 306) <= 1; flappy_W(10, 307) <= 1; flappy_W(10, 308) <= 1; flappy_W(10, 309) <= 1; flappy_W(10, 310) <= 1; flappy_W(10, 311) <= 1; flappy_W(10, 312) <= 1; flappy_W(10, 313) <= 1; flappy_W(10, 314) <= 1; flappy_W(10, 315) <= 1; flappy_W(10, 316) <= 1; flappy_W(10, 317) <= 1; flappy_W(10, 318) <= 0; flappy_W(10, 319) <= 0; flappy_W(10, 320) <= 0; flappy_W(10, 321) <= 0; flappy_W(10, 322) <= 0; flappy_W(10, 323) <= 0; flappy_W(10, 324) <= 0; flappy_W(10, 325) <= 0; flappy_W(10, 326) <= 0; flappy_W(10, 327) <= 0; flappy_W(10, 328) <= 0; flappy_W(10, 329) <= 0; flappy_W(10, 330) <= 0; flappy_W(10, 331) <= 0; flappy_W(10, 332) <= 0; flappy_W(10, 333) <= 0; flappy_W(10, 334) <= 0; flappy_W(10, 335) <= 0; flappy_W(10, 336) <= 0; flappy_W(10, 337) <= 0; flappy_W(10, 338) <= 0; flappy_W(10, 339) <= 0; flappy_W(10, 340) <= 0; flappy_W(10, 341) <= 0; flappy_W(10, 342) <= 0; flappy_W(10, 343) <= 0; flappy_W(10, 344) <= 0; flappy_W(10, 345) <= 0; flappy_W(10, 346) <= 0; flappy_W(10, 347) <= 0; flappy_W(10, 348) <= 0; flappy_W(10, 349) <= 0; flappy_W(10, 350) <= 0; flappy_W(10, 351) <= 0; flappy_W(10, 352) <= 0; flappy_W(10, 353) <= 0; flappy_W(10, 354) <= 0; flappy_W(10, 355) <= 0; flappy_W(10, 356) <= 0; flappy_W(10, 357) <= 0; flappy_W(10, 358) <= 0; flappy_W(10, 359) <= 0; flappy_W(10, 360) <= 0; flappy_W(10, 361) <= 0; flappy_W(10, 362) <= 0; flappy_W(10, 363) <= 0; flappy_W(10, 364) <= 0; flappy_W(10, 365) <= 0; flappy_W(10, 366) <= 0; flappy_W(10, 367) <= 0; flappy_W(10, 368) <= 0; flappy_W(10, 369) <= 0; flappy_W(10, 370) <= 0; flappy_W(10, 371) <= 0; flappy_W(10, 372) <= 0; flappy_W(10, 373) <= 0; flappy_W(10, 374) <= 0; flappy_W(10, 375) <= 0; flappy_W(10, 376) <= 0; flappy_W(10, 377) <= 0; flappy_W(10, 378) <= 0; flappy_W(10, 379) <= 0; flappy_W(10, 380) <= 0; flappy_W(10, 381) <= 0; flappy_W(10, 382) <= 0; flappy_W(10, 383) <= 0; flappy_W(10, 384) <= 0; flappy_W(10, 385) <= 0; flappy_W(10, 386) <= 0; flappy_W(10, 387) <= 0; flappy_W(10, 388) <= 0; flappy_W(10, 389) <= 0; flappy_W(10, 390) <= 0; flappy_W(10, 391) <= 0; flappy_W(10, 392) <= 0; flappy_W(10, 393) <= 0; flappy_W(10, 394) <= 0; flappy_W(10, 395) <= 0; flappy_W(10, 396) <= 0; flappy_W(10, 397) <= 0; flappy_W(10, 398) <= 0; flappy_W(10, 399) <= 0; flappy_W(10, 400) <= 0; flappy_W(10, 401) <= 0; flappy_W(10, 402) <= 1; flappy_W(10, 403) <= 1; flappy_W(10, 404) <= 1; flappy_W(10, 405) <= 1; flappy_W(10, 406) <= 1; flappy_W(10, 407) <= 1; flappy_W(10, 408) <= 1; flappy_W(10, 409) <= 1; flappy_W(10, 410) <= 1; flappy_W(10, 411) <= 1; flappy_W(10, 412) <= 1; flappy_W(10, 413) <= 1; flappy_W(10, 414) <= 0; flappy_W(10, 415) <= 0; flappy_W(10, 416) <= 0; flappy_W(10, 417) <= 0; flappy_W(10, 418) <= 0; flappy_W(10, 419) <= 0; flappy_W(10, 420) <= 0; flappy_W(10, 421) <= 0; flappy_W(10, 422) <= 0; flappy_W(10, 423) <= 0; flappy_W(10, 424) <= 0; flappy_W(10, 425) <= 0; flappy_W(10, 426) <= 1; flappy_W(10, 427) <= 1; flappy_W(10, 428) <= 1; flappy_W(10, 429) <= 1; flappy_W(10, 430) <= 1; flappy_W(10, 431) <= 1; flappy_W(10, 432) <= 1; flappy_W(10, 433) <= 1; flappy_W(10, 434) <= 1; flappy_W(10, 435) <= 1; flappy_W(10, 436) <= 1; flappy_W(10, 437) <= 1; flappy_W(10, 438) <= 0; flappy_W(10, 439) <= 0; flappy_W(10, 440) <= 0; flappy_W(10, 441) <= 0; flappy_W(10, 442) <= 0; flappy_W(10, 443) <= 0; flappy_W(10, 444) <= 0; flappy_W(10, 445) <= 0; flappy_W(10, 446) <= 0; flappy_W(10, 447) <= 0; flappy_W(10, 448) <= 0; flappy_W(10, 449) <= 0; flappy_W(10, 450) <= 0; flappy_W(10, 451) <= 0; flappy_W(10, 452) <= 0; flappy_W(10, 453) <= 0; flappy_W(10, 454) <= 0; flappy_W(10, 455) <= 0; flappy_W(10, 456) <= 0; flappy_W(10, 457) <= 0; flappy_W(10, 458) <= 0; flappy_W(10, 459) <= 0; flappy_W(10, 460) <= 0; flappy_W(10, 461) <= 0; flappy_W(10, 462) <= 0; flappy_W(10, 463) <= 0; flappy_W(10, 464) <= 0; flappy_W(10, 465) <= 0; flappy_W(10, 466) <= 0; flappy_W(10, 467) <= 0; flappy_W(10, 468) <= 1; flappy_W(10, 469) <= 1; flappy_W(10, 470) <= 1; flappy_W(10, 471) <= 1; flappy_W(10, 472) <= 1; flappy_W(10, 473) <= 1; flappy_W(10, 474) <= 1; flappy_W(10, 475) <= 1; flappy_W(10, 476) <= 1; flappy_W(10, 477) <= 1; flappy_W(10, 478) <= 1; flappy_W(10, 479) <= 1; flappy_W(10, 480) <= 0; flappy_W(10, 481) <= 0; flappy_W(10, 482) <= 0; flappy_W(10, 483) <= 0; flappy_W(10, 484) <= 0; flappy_W(10, 485) <= 0; flappy_W(10, 486) <= 0; flappy_W(10, 487) <= 0; flappy_W(10, 488) <= 0; flappy_W(10, 489) <= 0; flappy_W(10, 490) <= 0; flappy_W(10, 491) <= 0; flappy_W(10, 492) <= 0; flappy_W(10, 493) <= 0; flappy_W(10, 494) <= 0; flappy_W(10, 495) <= 0; flappy_W(10, 496) <= 0; flappy_W(10, 497) <= 0; flappy_W(10, 498) <= 0; flappy_W(10, 499) <= 0; flappy_W(10, 500) <= 0; flappy_W(10, 501) <= 0; flappy_W(10, 502) <= 0; flappy_W(10, 503) <= 0; flappy_W(10, 504) <= 0; flappy_W(10, 505) <= 0; flappy_W(10, 506) <= 0; flappy_W(10, 507) <= 0; flappy_W(10, 508) <= 0; flappy_W(10, 509) <= 0; flappy_W(10, 510) <= 1; flappy_W(10, 511) <= 1; flappy_W(10, 512) <= 1; flappy_W(10, 513) <= 1; flappy_W(10, 514) <= 1; flappy_W(10, 515) <= 1; flappy_W(10, 516) <= 1; flappy_W(10, 517) <= 1; flappy_W(10, 518) <= 1; flappy_W(10, 519) <= 1; flappy_W(10, 520) <= 1; flappy_W(10, 521) <= 1; flappy_W(10, 522) <= 0; flappy_W(10, 523) <= 0; flappy_W(10, 524) <= 0; flappy_W(10, 525) <= 0; flappy_W(10, 526) <= 0; flappy_W(10, 527) <= 0; flappy_W(10, 528) <= 0; flappy_W(10, 529) <= 0; flappy_W(10, 530) <= 0; flappy_W(10, 531) <= 0; flappy_W(10, 532) <= 0; flappy_W(10, 533) <= 0; flappy_W(10, 534) <= 1; flappy_W(10, 535) <= 1; flappy_W(10, 536) <= 1; flappy_W(10, 537) <= 1; flappy_W(10, 538) <= 1; flappy_W(10, 539) <= 1; flappy_W(10, 540) <= 1; flappy_W(10, 541) <= 1; flappy_W(10, 542) <= 1; flappy_W(10, 543) <= 1; flappy_W(10, 544) <= 1; flappy_W(10, 545) <= 1; flappy_W(10, 546) <= 0; flappy_W(10, 547) <= 0; flappy_W(10, 548) <= 0; flappy_W(10, 549) <= 0; flappy_W(10, 550) <= 0; flappy_W(10, 551) <= 0; flappy_W(10, 552) <= 0; flappy_W(10, 553) <= 0; flappy_W(10, 554) <= 0; flappy_W(10, 555) <= 0; flappy_W(10, 556) <= 0; flappy_W(10, 557) <= 0; flappy_W(10, 558) <= 0; flappy_W(10, 559) <= 0; flappy_W(10, 560) <= 0; flappy_W(10, 561) <= 0; flappy_W(10, 562) <= 0; flappy_W(10, 563) <= 0; flappy_W(10, 564) <= 1; flappy_W(10, 565) <= 1; flappy_W(10, 566) <= 1; flappy_W(10, 567) <= 1; flappy_W(10, 568) <= 1; flappy_W(10, 569) <= 1; flappy_W(10, 570) <= 1; flappy_W(10, 571) <= 1; flappy_W(10, 572) <= 1; flappy_W(10, 573) <= 1; flappy_W(10, 574) <= 1; flappy_W(10, 575) <= 1; flappy_W(10, 576) <= 0; flappy_W(10, 577) <= 0; flappy_W(10, 578) <= 0; flappy_W(10, 579) <= 0; flappy_W(10, 580) <= 0; flappy_W(10, 581) <= 0; flappy_W(10, 582) <= 1; flappy_W(10, 583) <= 1; flappy_W(10, 584) <= 1; flappy_W(10, 585) <= 1; flappy_W(10, 586) <= 1; flappy_W(10, 587) <= 1; flappy_W(10, 588) <= 1; flappy_W(10, 589) <= 1; flappy_W(10, 590) <= 1; flappy_W(10, 591) <= 1; flappy_W(10, 592) <= 1; flappy_W(10, 593) <= 1; 
flappy_W(11, 0) <= 0; flappy_W(11, 1) <= 0; flappy_W(11, 2) <= 0; flappy_W(11, 3) <= 0; flappy_W(11, 4) <= 0; flappy_W(11, 5) <= 0; flappy_W(11, 6) <= 1; flappy_W(11, 7) <= 1; flappy_W(11, 8) <= 1; flappy_W(11, 9) <= 1; flappy_W(11, 10) <= 1; flappy_W(11, 11) <= 1; flappy_W(11, 12) <= 1; flappy_W(11, 13) <= 1; flappy_W(11, 14) <= 1; flappy_W(11, 15) <= 1; flappy_W(11, 16) <= 1; flappy_W(11, 17) <= 1; flappy_W(11, 18) <= 0; flappy_W(11, 19) <= 0; flappy_W(11, 20) <= 0; flappy_W(11, 21) <= 0; flappy_W(11, 22) <= 0; flappy_W(11, 23) <= 0; flappy_W(11, 24) <= 0; flappy_W(11, 25) <= 0; flappy_W(11, 26) <= 0; flappy_W(11, 27) <= 0; flappy_W(11, 28) <= 0; flappy_W(11, 29) <= 0; flappy_W(11, 30) <= 1; flappy_W(11, 31) <= 1; flappy_W(11, 32) <= 1; flappy_W(11, 33) <= 1; flappy_W(11, 34) <= 1; flappy_W(11, 35) <= 1; flappy_W(11, 36) <= 1; flappy_W(11, 37) <= 1; flappy_W(11, 38) <= 1; flappy_W(11, 39) <= 1; flappy_W(11, 40) <= 1; flappy_W(11, 41) <= 1; flappy_W(11, 42) <= 0; flappy_W(11, 43) <= 0; flappy_W(11, 44) <= 0; flappy_W(11, 45) <= 0; flappy_W(11, 46) <= 0; flappy_W(11, 47) <= 0; flappy_W(11, 48) <= 0; flappy_W(11, 49) <= 0; flappy_W(11, 50) <= 0; flappy_W(11, 51) <= 0; flappy_W(11, 52) <= 0; flappy_W(11, 53) <= 0; flappy_W(11, 54) <= 0; flappy_W(11, 55) <= 0; flappy_W(11, 56) <= 0; flappy_W(11, 57) <= 0; flappy_W(11, 58) <= 0; flappy_W(11, 59) <= 0; flappy_W(11, 60) <= 1; flappy_W(11, 61) <= 1; flappy_W(11, 62) <= 1; flappy_W(11, 63) <= 1; flappy_W(11, 64) <= 1; flappy_W(11, 65) <= 1; flappy_W(11, 66) <= 1; flappy_W(11, 67) <= 1; flappy_W(11, 68) <= 1; flappy_W(11, 69) <= 1; flappy_W(11, 70) <= 1; flappy_W(11, 71) <= 1; flappy_W(11, 72) <= 0; flappy_W(11, 73) <= 0; flappy_W(11, 74) <= 0; flappy_W(11, 75) <= 0; flappy_W(11, 76) <= 0; flappy_W(11, 77) <= 0; flappy_W(11, 78) <= 0; flappy_W(11, 79) <= 0; flappy_W(11, 80) <= 0; flappy_W(11, 81) <= 0; flappy_W(11, 82) <= 0; flappy_W(11, 83) <= 0; flappy_W(11, 84) <= 0; flappy_W(11, 85) <= 0; flappy_W(11, 86) <= 0; flappy_W(11, 87) <= 0; flappy_W(11, 88) <= 0; flappy_W(11, 89) <= 0; flappy_W(11, 90) <= 0; flappy_W(11, 91) <= 0; flappy_W(11, 92) <= 0; flappy_W(11, 93) <= 0; flappy_W(11, 94) <= 0; flappy_W(11, 95) <= 0; flappy_W(11, 96) <= 0; flappy_W(11, 97) <= 0; flappy_W(11, 98) <= 0; flappy_W(11, 99) <= 0; flappy_W(11, 100) <= 0; flappy_W(11, 101) <= 0; flappy_W(11, 102) <= 0; flappy_W(11, 103) <= 0; flappy_W(11, 104) <= 0; flappy_W(11, 105) <= 0; flappy_W(11, 106) <= 0; flappy_W(11, 107) <= 0; flappy_W(11, 108) <= 0; flappy_W(11, 109) <= 0; flappy_W(11, 110) <= 0; flappy_W(11, 111) <= 0; flappy_W(11, 112) <= 0; flappy_W(11, 113) <= 0; flappy_W(11, 114) <= 0; flappy_W(11, 115) <= 0; flappy_W(11, 116) <= 0; flappy_W(11, 117) <= 0; flappy_W(11, 118) <= 0; flappy_W(11, 119) <= 0; flappy_W(11, 120) <= 1; flappy_W(11, 121) <= 1; flappy_W(11, 122) <= 1; flappy_W(11, 123) <= 1; flappy_W(11, 124) <= 1; flappy_W(11, 125) <= 1; flappy_W(11, 126) <= 1; flappy_W(11, 127) <= 1; flappy_W(11, 128) <= 1; flappy_W(11, 129) <= 1; flappy_W(11, 130) <= 1; flappy_W(11, 131) <= 1; flappy_W(11, 132) <= 1; flappy_W(11, 133) <= 1; flappy_W(11, 134) <= 1; flappy_W(11, 135) <= 1; flappy_W(11, 136) <= 1; flappy_W(11, 137) <= 1; flappy_W(11, 138) <= 0; flappy_W(11, 139) <= 0; flappy_W(11, 140) <= 0; flappy_W(11, 141) <= 0; flappy_W(11, 142) <= 0; flappy_W(11, 143) <= 0; flappy_W(11, 144) <= 0; flappy_W(11, 145) <= 0; flappy_W(11, 146) <= 0; flappy_W(11, 147) <= 0; flappy_W(11, 148) <= 0; flappy_W(11, 149) <= 0; flappy_W(11, 150) <= 0; flappy_W(11, 151) <= 0; flappy_W(11, 152) <= 0; flappy_W(11, 153) <= 0; flappy_W(11, 154) <= 0; flappy_W(11, 155) <= 0; flappy_W(11, 156) <= 0; flappy_W(11, 157) <= 0; flappy_W(11, 158) <= 0; flappy_W(11, 159) <= 0; flappy_W(11, 160) <= 0; flappy_W(11, 161) <= 0; flappy_W(11, 162) <= 0; flappy_W(11, 163) <= 0; flappy_W(11, 164) <= 0; flappy_W(11, 165) <= 0; flappy_W(11, 166) <= 0; flappy_W(11, 167) <= 0; flappy_W(11, 168) <= 1; flappy_W(11, 169) <= 1; flappy_W(11, 170) <= 1; flappy_W(11, 171) <= 1; flappy_W(11, 172) <= 1; flappy_W(11, 173) <= 1; flappy_W(11, 174) <= 1; flappy_W(11, 175) <= 1; flappy_W(11, 176) <= 1; flappy_W(11, 177) <= 1; flappy_W(11, 178) <= 1; flappy_W(11, 179) <= 1; flappy_W(11, 180) <= 0; flappy_W(11, 181) <= 0; flappy_W(11, 182) <= 0; flappy_W(11, 183) <= 0; flappy_W(11, 184) <= 0; flappy_W(11, 185) <= 0; flappy_W(11, 186) <= 0; flappy_W(11, 187) <= 0; flappy_W(11, 188) <= 0; flappy_W(11, 189) <= 0; flappy_W(11, 190) <= 0; flappy_W(11, 191) <= 0; flappy_W(11, 192) <= 1; flappy_W(11, 193) <= 1; flappy_W(11, 194) <= 1; flappy_W(11, 195) <= 1; flappy_W(11, 196) <= 1; flappy_W(11, 197) <= 1; flappy_W(11, 198) <= 1; flappy_W(11, 199) <= 1; flappy_W(11, 200) <= 1; flappy_W(11, 201) <= 1; flappy_W(11, 202) <= 1; flappy_W(11, 203) <= 1; flappy_W(11, 204) <= 0; flappy_W(11, 205) <= 0; flappy_W(11, 206) <= 0; flappy_W(11, 207) <= 0; flappy_W(11, 208) <= 0; flappy_W(11, 209) <= 0; flappy_W(11, 210) <= 0; flappy_W(11, 211) <= 0; flappy_W(11, 212) <= 0; flappy_W(11, 213) <= 0; flappy_W(11, 214) <= 0; flappy_W(11, 215) <= 0; flappy_W(11, 216) <= 0; flappy_W(11, 217) <= 0; flappy_W(11, 218) <= 0; flappy_W(11, 219) <= 0; flappy_W(11, 220) <= 0; flappy_W(11, 221) <= 0; flappy_W(11, 222) <= 1; flappy_W(11, 223) <= 1; flappy_W(11, 224) <= 1; flappy_W(11, 225) <= 1; flappy_W(11, 226) <= 1; flappy_W(11, 227) <= 1; flappy_W(11, 228) <= 1; flappy_W(11, 229) <= 1; flappy_W(11, 230) <= 1; flappy_W(11, 231) <= 1; flappy_W(11, 232) <= 1; flappy_W(11, 233) <= 1; flappy_W(11, 234) <= 0; flappy_W(11, 235) <= 0; flappy_W(11, 236) <= 0; flappy_W(11, 237) <= 0; flappy_W(11, 238) <= 0; flappy_W(11, 239) <= 0; flappy_W(11, 240) <= 0; flappy_W(11, 241) <= 0; flappy_W(11, 242) <= 0; flappy_W(11, 243) <= 0; flappy_W(11, 244) <= 0; flappy_W(11, 245) <= 0; flappy_W(11, 246) <= 1; flappy_W(11, 247) <= 1; flappy_W(11, 248) <= 1; flappy_W(11, 249) <= 1; flappy_W(11, 250) <= 1; flappy_W(11, 251) <= 1; flappy_W(11, 252) <= 1; flappy_W(11, 253) <= 1; flappy_W(11, 254) <= 1; flappy_W(11, 255) <= 1; flappy_W(11, 256) <= 1; flappy_W(11, 257) <= 1; flappy_W(11, 258) <= 0; flappy_W(11, 259) <= 0; flappy_W(11, 260) <= 0; flappy_W(11, 261) <= 0; flappy_W(11, 262) <= 0; flappy_W(11, 263) <= 0; flappy_W(11, 264) <= 0; flappy_W(11, 265) <= 0; flappy_W(11, 266) <= 0; flappy_W(11, 267) <= 0; flappy_W(11, 268) <= 0; flappy_W(11, 269) <= 0; flappy_W(11, 270) <= 1; flappy_W(11, 271) <= 1; flappy_W(11, 272) <= 1; flappy_W(11, 273) <= 1; flappy_W(11, 274) <= 1; flappy_W(11, 275) <= 1; flappy_W(11, 276) <= 1; flappy_W(11, 277) <= 1; flappy_W(11, 278) <= 1; flappy_W(11, 279) <= 1; flappy_W(11, 280) <= 1; flappy_W(11, 281) <= 1; flappy_W(11, 282) <= 0; flappy_W(11, 283) <= 0; flappy_W(11, 284) <= 0; flappy_W(11, 285) <= 0; flappy_W(11, 286) <= 0; flappy_W(11, 287) <= 0; flappy_W(11, 288) <= 0; flappy_W(11, 289) <= 0; flappy_W(11, 290) <= 0; flappy_W(11, 291) <= 0; flappy_W(11, 292) <= 0; flappy_W(11, 293) <= 0; flappy_W(11, 294) <= 0; flappy_W(11, 295) <= 0; flappy_W(11, 296) <= 0; flappy_W(11, 297) <= 0; flappy_W(11, 298) <= 0; flappy_W(11, 299) <= 0; flappy_W(11, 300) <= 0; flappy_W(11, 301) <= 0; flappy_W(11, 302) <= 0; flappy_W(11, 303) <= 0; flappy_W(11, 304) <= 0; flappy_W(11, 305) <= 0; flappy_W(11, 306) <= 1; flappy_W(11, 307) <= 1; flappy_W(11, 308) <= 1; flappy_W(11, 309) <= 1; flappy_W(11, 310) <= 1; flappy_W(11, 311) <= 1; flappy_W(11, 312) <= 1; flappy_W(11, 313) <= 1; flappy_W(11, 314) <= 1; flappy_W(11, 315) <= 1; flappy_W(11, 316) <= 1; flappy_W(11, 317) <= 1; flappy_W(11, 318) <= 0; flappy_W(11, 319) <= 0; flappy_W(11, 320) <= 0; flappy_W(11, 321) <= 0; flappy_W(11, 322) <= 0; flappy_W(11, 323) <= 0; flappy_W(11, 324) <= 0; flappy_W(11, 325) <= 0; flappy_W(11, 326) <= 0; flappy_W(11, 327) <= 0; flappy_W(11, 328) <= 0; flappy_W(11, 329) <= 0; flappy_W(11, 330) <= 0; flappy_W(11, 331) <= 0; flappy_W(11, 332) <= 0; flappy_W(11, 333) <= 0; flappy_W(11, 334) <= 0; flappy_W(11, 335) <= 0; flappy_W(11, 336) <= 0; flappy_W(11, 337) <= 0; flappy_W(11, 338) <= 0; flappy_W(11, 339) <= 0; flappy_W(11, 340) <= 0; flappy_W(11, 341) <= 0; flappy_W(11, 342) <= 0; flappy_W(11, 343) <= 0; flappy_W(11, 344) <= 0; flappy_W(11, 345) <= 0; flappy_W(11, 346) <= 0; flappy_W(11, 347) <= 0; flappy_W(11, 348) <= 0; flappy_W(11, 349) <= 0; flappy_W(11, 350) <= 0; flappy_W(11, 351) <= 0; flappy_W(11, 352) <= 0; flappy_W(11, 353) <= 0; flappy_W(11, 354) <= 0; flappy_W(11, 355) <= 0; flappy_W(11, 356) <= 0; flappy_W(11, 357) <= 0; flappy_W(11, 358) <= 0; flappy_W(11, 359) <= 0; flappy_W(11, 360) <= 0; flappy_W(11, 361) <= 0; flappy_W(11, 362) <= 0; flappy_W(11, 363) <= 0; flappy_W(11, 364) <= 0; flappy_W(11, 365) <= 0; flappy_W(11, 366) <= 0; flappy_W(11, 367) <= 0; flappy_W(11, 368) <= 0; flappy_W(11, 369) <= 0; flappy_W(11, 370) <= 0; flappy_W(11, 371) <= 0; flappy_W(11, 372) <= 0; flappy_W(11, 373) <= 0; flappy_W(11, 374) <= 0; flappy_W(11, 375) <= 0; flappy_W(11, 376) <= 0; flappy_W(11, 377) <= 0; flappy_W(11, 378) <= 0; flappy_W(11, 379) <= 0; flappy_W(11, 380) <= 0; flappy_W(11, 381) <= 0; flappy_W(11, 382) <= 0; flappy_W(11, 383) <= 0; flappy_W(11, 384) <= 0; flappy_W(11, 385) <= 0; flappy_W(11, 386) <= 0; flappy_W(11, 387) <= 0; flappy_W(11, 388) <= 0; flappy_W(11, 389) <= 0; flappy_W(11, 390) <= 0; flappy_W(11, 391) <= 0; flappy_W(11, 392) <= 0; flappy_W(11, 393) <= 0; flappy_W(11, 394) <= 0; flappy_W(11, 395) <= 0; flappy_W(11, 396) <= 0; flappy_W(11, 397) <= 0; flappy_W(11, 398) <= 0; flappy_W(11, 399) <= 0; flappy_W(11, 400) <= 0; flappy_W(11, 401) <= 0; flappy_W(11, 402) <= 1; flappy_W(11, 403) <= 1; flappy_W(11, 404) <= 1; flappy_W(11, 405) <= 1; flappy_W(11, 406) <= 1; flappy_W(11, 407) <= 1; flappy_W(11, 408) <= 1; flappy_W(11, 409) <= 1; flappy_W(11, 410) <= 1; flappy_W(11, 411) <= 1; flappy_W(11, 412) <= 1; flappy_W(11, 413) <= 1; flappy_W(11, 414) <= 0; flappy_W(11, 415) <= 0; flappy_W(11, 416) <= 0; flappy_W(11, 417) <= 0; flappy_W(11, 418) <= 0; flappy_W(11, 419) <= 0; flappy_W(11, 420) <= 0; flappy_W(11, 421) <= 0; flappy_W(11, 422) <= 0; flappy_W(11, 423) <= 0; flappy_W(11, 424) <= 0; flappy_W(11, 425) <= 0; flappy_W(11, 426) <= 1; flappy_W(11, 427) <= 1; flappy_W(11, 428) <= 1; flappy_W(11, 429) <= 1; flappy_W(11, 430) <= 1; flappy_W(11, 431) <= 1; flappy_W(11, 432) <= 1; flappy_W(11, 433) <= 1; flappy_W(11, 434) <= 1; flappy_W(11, 435) <= 1; flappy_W(11, 436) <= 1; flappy_W(11, 437) <= 1; flappy_W(11, 438) <= 0; flappy_W(11, 439) <= 0; flappy_W(11, 440) <= 0; flappy_W(11, 441) <= 0; flappy_W(11, 442) <= 0; flappy_W(11, 443) <= 0; flappy_W(11, 444) <= 0; flappy_W(11, 445) <= 0; flappy_W(11, 446) <= 0; flappy_W(11, 447) <= 0; flappy_W(11, 448) <= 0; flappy_W(11, 449) <= 0; flappy_W(11, 450) <= 0; flappy_W(11, 451) <= 0; flappy_W(11, 452) <= 0; flappy_W(11, 453) <= 0; flappy_W(11, 454) <= 0; flappy_W(11, 455) <= 0; flappy_W(11, 456) <= 0; flappy_W(11, 457) <= 0; flappy_W(11, 458) <= 0; flappy_W(11, 459) <= 0; flappy_W(11, 460) <= 0; flappy_W(11, 461) <= 0; flappy_W(11, 462) <= 0; flappy_W(11, 463) <= 0; flappy_W(11, 464) <= 0; flappy_W(11, 465) <= 0; flappy_W(11, 466) <= 0; flappy_W(11, 467) <= 0; flappy_W(11, 468) <= 1; flappy_W(11, 469) <= 1; flappy_W(11, 470) <= 1; flappy_W(11, 471) <= 1; flappy_W(11, 472) <= 1; flappy_W(11, 473) <= 1; flappy_W(11, 474) <= 1; flappy_W(11, 475) <= 1; flappy_W(11, 476) <= 1; flappy_W(11, 477) <= 1; flappy_W(11, 478) <= 1; flappy_W(11, 479) <= 1; flappy_W(11, 480) <= 0; flappy_W(11, 481) <= 0; flappy_W(11, 482) <= 0; flappy_W(11, 483) <= 0; flappy_W(11, 484) <= 0; flappy_W(11, 485) <= 0; flappy_W(11, 486) <= 0; flappy_W(11, 487) <= 0; flappy_W(11, 488) <= 0; flappy_W(11, 489) <= 0; flappy_W(11, 490) <= 0; flappy_W(11, 491) <= 0; flappy_W(11, 492) <= 0; flappy_W(11, 493) <= 0; flappy_W(11, 494) <= 0; flappy_W(11, 495) <= 0; flappy_W(11, 496) <= 0; flappy_W(11, 497) <= 0; flappy_W(11, 498) <= 0; flappy_W(11, 499) <= 0; flappy_W(11, 500) <= 0; flappy_W(11, 501) <= 0; flappy_W(11, 502) <= 0; flappy_W(11, 503) <= 0; flappy_W(11, 504) <= 0; flappy_W(11, 505) <= 0; flappy_W(11, 506) <= 0; flappy_W(11, 507) <= 0; flappy_W(11, 508) <= 0; flappy_W(11, 509) <= 0; flappy_W(11, 510) <= 1; flappy_W(11, 511) <= 1; flappy_W(11, 512) <= 1; flappy_W(11, 513) <= 1; flappy_W(11, 514) <= 1; flappy_W(11, 515) <= 1; flappy_W(11, 516) <= 1; flappy_W(11, 517) <= 1; flappy_W(11, 518) <= 1; flappy_W(11, 519) <= 1; flappy_W(11, 520) <= 1; flappy_W(11, 521) <= 1; flappy_W(11, 522) <= 0; flappy_W(11, 523) <= 0; flappy_W(11, 524) <= 0; flappy_W(11, 525) <= 0; flappy_W(11, 526) <= 0; flappy_W(11, 527) <= 0; flappy_W(11, 528) <= 0; flappy_W(11, 529) <= 0; flappy_W(11, 530) <= 0; flappy_W(11, 531) <= 0; flappy_W(11, 532) <= 0; flappy_W(11, 533) <= 0; flappy_W(11, 534) <= 1; flappy_W(11, 535) <= 1; flappy_W(11, 536) <= 1; flappy_W(11, 537) <= 1; flappy_W(11, 538) <= 1; flappy_W(11, 539) <= 1; flappy_W(11, 540) <= 1; flappy_W(11, 541) <= 1; flappy_W(11, 542) <= 1; flappy_W(11, 543) <= 1; flappy_W(11, 544) <= 1; flappy_W(11, 545) <= 1; flappy_W(11, 546) <= 0; flappy_W(11, 547) <= 0; flappy_W(11, 548) <= 0; flappy_W(11, 549) <= 0; flappy_W(11, 550) <= 0; flappy_W(11, 551) <= 0; flappy_W(11, 552) <= 0; flappy_W(11, 553) <= 0; flappy_W(11, 554) <= 0; flappy_W(11, 555) <= 0; flappy_W(11, 556) <= 0; flappy_W(11, 557) <= 0; flappy_W(11, 558) <= 0; flappy_W(11, 559) <= 0; flappy_W(11, 560) <= 0; flappy_W(11, 561) <= 0; flappy_W(11, 562) <= 0; flappy_W(11, 563) <= 0; flappy_W(11, 564) <= 1; flappy_W(11, 565) <= 1; flappy_W(11, 566) <= 1; flappy_W(11, 567) <= 1; flappy_W(11, 568) <= 1; flappy_W(11, 569) <= 1; flappy_W(11, 570) <= 1; flappy_W(11, 571) <= 1; flappy_W(11, 572) <= 1; flappy_W(11, 573) <= 1; flappy_W(11, 574) <= 1; flappy_W(11, 575) <= 1; flappy_W(11, 576) <= 0; flappy_W(11, 577) <= 0; flappy_W(11, 578) <= 0; flappy_W(11, 579) <= 0; flappy_W(11, 580) <= 0; flappy_W(11, 581) <= 0; flappy_W(11, 582) <= 1; flappy_W(11, 583) <= 1; flappy_W(11, 584) <= 1; flappy_W(11, 585) <= 1; flappy_W(11, 586) <= 1; flappy_W(11, 587) <= 1; flappy_W(11, 588) <= 1; flappy_W(11, 589) <= 1; flappy_W(11, 590) <= 1; flappy_W(11, 591) <= 1; flappy_W(11, 592) <= 1; flappy_W(11, 593) <= 1; 
flappy_W(12, 0) <= 0; flappy_W(12, 1) <= 0; flappy_W(12, 2) <= 0; flappy_W(12, 3) <= 0; flappy_W(12, 4) <= 0; flappy_W(12, 5) <= 0; flappy_W(12, 6) <= 1; flappy_W(12, 7) <= 1; flappy_W(12, 8) <= 1; flappy_W(12, 9) <= 1; flappy_W(12, 10) <= 1; flappy_W(12, 11) <= 1; flappy_W(12, 12) <= 1; flappy_W(12, 13) <= 1; flappy_W(12, 14) <= 1; flappy_W(12, 15) <= 1; flappy_W(12, 16) <= 1; flappy_W(12, 17) <= 1; flappy_W(12, 18) <= 0; flappy_W(12, 19) <= 0; flappy_W(12, 20) <= 0; flappy_W(12, 21) <= 0; flappy_W(12, 22) <= 0; flappy_W(12, 23) <= 0; flappy_W(12, 24) <= 0; flappy_W(12, 25) <= 0; flappy_W(12, 26) <= 0; flappy_W(12, 27) <= 0; flappy_W(12, 28) <= 0; flappy_W(12, 29) <= 0; flappy_W(12, 30) <= 0; flappy_W(12, 31) <= 0; flappy_W(12, 32) <= 0; flappy_W(12, 33) <= 0; flappy_W(12, 34) <= 0; flappy_W(12, 35) <= 0; flappy_W(12, 36) <= 1; flappy_W(12, 37) <= 1; flappy_W(12, 38) <= 1; flappy_W(12, 39) <= 1; flappy_W(12, 40) <= 1; flappy_W(12, 41) <= 1; flappy_W(12, 42) <= 0; flappy_W(12, 43) <= 0; flappy_W(12, 44) <= 0; flappy_W(12, 45) <= 0; flappy_W(12, 46) <= 0; flappy_W(12, 47) <= 0; flappy_W(12, 48) <= 0; flappy_W(12, 49) <= 0; flappy_W(12, 50) <= 0; flappy_W(12, 51) <= 0; flappy_W(12, 52) <= 0; flappy_W(12, 53) <= 0; flappy_W(12, 54) <= 0; flappy_W(12, 55) <= 0; flappy_W(12, 56) <= 0; flappy_W(12, 57) <= 0; flappy_W(12, 58) <= 0; flappy_W(12, 59) <= 0; flappy_W(12, 60) <= 1; flappy_W(12, 61) <= 1; flappy_W(12, 62) <= 1; flappy_W(12, 63) <= 1; flappy_W(12, 64) <= 1; flappy_W(12, 65) <= 1; flappy_W(12, 66) <= 1; flappy_W(12, 67) <= 1; flappy_W(12, 68) <= 1; flappy_W(12, 69) <= 1; flappy_W(12, 70) <= 1; flappy_W(12, 71) <= 1; flappy_W(12, 72) <= 0; flappy_W(12, 73) <= 0; flappy_W(12, 74) <= 0; flappy_W(12, 75) <= 0; flappy_W(12, 76) <= 0; flappy_W(12, 77) <= 0; flappy_W(12, 78) <= 0; flappy_W(12, 79) <= 0; flappy_W(12, 80) <= 0; flappy_W(12, 81) <= 0; flappy_W(12, 82) <= 0; flappy_W(12, 83) <= 0; flappy_W(12, 84) <= 0; flappy_W(12, 85) <= 0; flappy_W(12, 86) <= 0; flappy_W(12, 87) <= 0; flappy_W(12, 88) <= 0; flappy_W(12, 89) <= 0; flappy_W(12, 90) <= 0; flappy_W(12, 91) <= 0; flappy_W(12, 92) <= 0; flappy_W(12, 93) <= 0; flappy_W(12, 94) <= 0; flappy_W(12, 95) <= 0; flappy_W(12, 96) <= 0; flappy_W(12, 97) <= 0; flappy_W(12, 98) <= 0; flappy_W(12, 99) <= 0; flappy_W(12, 100) <= 0; flappy_W(12, 101) <= 0; flappy_W(12, 102) <= 0; flappy_W(12, 103) <= 0; flappy_W(12, 104) <= 0; flappy_W(12, 105) <= 0; flappy_W(12, 106) <= 0; flappy_W(12, 107) <= 0; flappy_W(12, 108) <= 0; flappy_W(12, 109) <= 0; flappy_W(12, 110) <= 0; flappy_W(12, 111) <= 0; flappy_W(12, 112) <= 0; flappy_W(12, 113) <= 0; flappy_W(12, 114) <= 1; flappy_W(12, 115) <= 1; flappy_W(12, 116) <= 1; flappy_W(12, 117) <= 1; flappy_W(12, 118) <= 1; flappy_W(12, 119) <= 1; flappy_W(12, 120) <= 1; flappy_W(12, 121) <= 1; flappy_W(12, 122) <= 1; flappy_W(12, 123) <= 1; flappy_W(12, 124) <= 1; flappy_W(12, 125) <= 1; flappy_W(12, 126) <= 0; flappy_W(12, 127) <= 0; flappy_W(12, 128) <= 0; flappy_W(12, 129) <= 0; flappy_W(12, 130) <= 0; flappy_W(12, 131) <= 0; flappy_W(12, 132) <= 1; flappy_W(12, 133) <= 1; flappy_W(12, 134) <= 1; flappy_W(12, 135) <= 1; flappy_W(12, 136) <= 1; flappy_W(12, 137) <= 1; flappy_W(12, 138) <= 1; flappy_W(12, 139) <= 1; flappy_W(12, 140) <= 1; flappy_W(12, 141) <= 1; flappy_W(12, 142) <= 1; flappy_W(12, 143) <= 1; flappy_W(12, 144) <= 0; flappy_W(12, 145) <= 0; flappy_W(12, 146) <= 0; flappy_W(12, 147) <= 0; flappy_W(12, 148) <= 0; flappy_W(12, 149) <= 0; flappy_W(12, 150) <= 0; flappy_W(12, 151) <= 0; flappy_W(12, 152) <= 0; flappy_W(12, 153) <= 0; flappy_W(12, 154) <= 0; flappy_W(12, 155) <= 0; flappy_W(12, 156) <= 0; flappy_W(12, 157) <= 0; flappy_W(12, 158) <= 0; flappy_W(12, 159) <= 0; flappy_W(12, 160) <= 0; flappy_W(12, 161) <= 0; flappy_W(12, 162) <= 0; flappy_W(12, 163) <= 0; flappy_W(12, 164) <= 0; flappy_W(12, 165) <= 0; flappy_W(12, 166) <= 0; flappy_W(12, 167) <= 0; flappy_W(12, 168) <= 1; flappy_W(12, 169) <= 1; flappy_W(12, 170) <= 1; flappy_W(12, 171) <= 1; flappy_W(12, 172) <= 1; flappy_W(12, 173) <= 1; flappy_W(12, 174) <= 1; flappy_W(12, 175) <= 1; flappy_W(12, 176) <= 1; flappy_W(12, 177) <= 1; flappy_W(12, 178) <= 1; flappy_W(12, 179) <= 1; flappy_W(12, 180) <= 0; flappy_W(12, 181) <= 0; flappy_W(12, 182) <= 0; flappy_W(12, 183) <= 0; flappy_W(12, 184) <= 0; flappy_W(12, 185) <= 0; flappy_W(12, 186) <= 0; flappy_W(12, 187) <= 0; flappy_W(12, 188) <= 0; flappy_W(12, 189) <= 0; flappy_W(12, 190) <= 0; flappy_W(12, 191) <= 0; flappy_W(12, 192) <= 1; flappy_W(12, 193) <= 1; flappy_W(12, 194) <= 1; flappy_W(12, 195) <= 1; flappy_W(12, 196) <= 1; flappy_W(12, 197) <= 1; flappy_W(12, 198) <= 1; flappy_W(12, 199) <= 1; flappy_W(12, 200) <= 1; flappy_W(12, 201) <= 1; flappy_W(12, 202) <= 1; flappy_W(12, 203) <= 1; flappy_W(12, 204) <= 0; flappy_W(12, 205) <= 0; flappy_W(12, 206) <= 0; flappy_W(12, 207) <= 0; flappy_W(12, 208) <= 0; flappy_W(12, 209) <= 0; flappy_W(12, 210) <= 0; flappy_W(12, 211) <= 0; flappy_W(12, 212) <= 0; flappy_W(12, 213) <= 0; flappy_W(12, 214) <= 0; flappy_W(12, 215) <= 0; flappy_W(12, 216) <= 0; flappy_W(12, 217) <= 0; flappy_W(12, 218) <= 0; flappy_W(12, 219) <= 0; flappy_W(12, 220) <= 0; flappy_W(12, 221) <= 0; flappy_W(12, 222) <= 1; flappy_W(12, 223) <= 1; flappy_W(12, 224) <= 1; flappy_W(12, 225) <= 1; flappy_W(12, 226) <= 1; flappy_W(12, 227) <= 1; flappy_W(12, 228) <= 1; flappy_W(12, 229) <= 1; flappy_W(12, 230) <= 1; flappy_W(12, 231) <= 1; flappy_W(12, 232) <= 1; flappy_W(12, 233) <= 1; flappy_W(12, 234) <= 0; flappy_W(12, 235) <= 0; flappy_W(12, 236) <= 0; flappy_W(12, 237) <= 0; flappy_W(12, 238) <= 0; flappy_W(12, 239) <= 0; flappy_W(12, 240) <= 0; flappy_W(12, 241) <= 0; flappy_W(12, 242) <= 0; flappy_W(12, 243) <= 0; flappy_W(12, 244) <= 0; flappy_W(12, 245) <= 0; flappy_W(12, 246) <= 1; flappy_W(12, 247) <= 1; flappy_W(12, 248) <= 1; flappy_W(12, 249) <= 1; flappy_W(12, 250) <= 1; flappy_W(12, 251) <= 1; flappy_W(12, 252) <= 1; flappy_W(12, 253) <= 1; flappy_W(12, 254) <= 1; flappy_W(12, 255) <= 1; flappy_W(12, 256) <= 1; flappy_W(12, 257) <= 1; flappy_W(12, 258) <= 0; flappy_W(12, 259) <= 0; flappy_W(12, 260) <= 0; flappy_W(12, 261) <= 0; flappy_W(12, 262) <= 0; flappy_W(12, 263) <= 0; flappy_W(12, 264) <= 0; flappy_W(12, 265) <= 0; flappy_W(12, 266) <= 0; flappy_W(12, 267) <= 0; flappy_W(12, 268) <= 0; flappy_W(12, 269) <= 0; flappy_W(12, 270) <= 1; flappy_W(12, 271) <= 1; flappy_W(12, 272) <= 1; flappy_W(12, 273) <= 1; flappy_W(12, 274) <= 1; flappy_W(12, 275) <= 1; flappy_W(12, 276) <= 1; flappy_W(12, 277) <= 1; flappy_W(12, 278) <= 1; flappy_W(12, 279) <= 1; flappy_W(12, 280) <= 1; flappy_W(12, 281) <= 1; flappy_W(12, 282) <= 0; flappy_W(12, 283) <= 0; flappy_W(12, 284) <= 0; flappy_W(12, 285) <= 0; flappy_W(12, 286) <= 0; flappy_W(12, 287) <= 0; flappy_W(12, 288) <= 0; flappy_W(12, 289) <= 0; flappy_W(12, 290) <= 0; flappy_W(12, 291) <= 0; flappy_W(12, 292) <= 0; flappy_W(12, 293) <= 0; flappy_W(12, 294) <= 0; flappy_W(12, 295) <= 0; flappy_W(12, 296) <= 0; flappy_W(12, 297) <= 0; flappy_W(12, 298) <= 0; flappy_W(12, 299) <= 0; flappy_W(12, 300) <= 0; flappy_W(12, 301) <= 0; flappy_W(12, 302) <= 0; flappy_W(12, 303) <= 0; flappy_W(12, 304) <= 0; flappy_W(12, 305) <= 0; flappy_W(12, 306) <= 1; flappy_W(12, 307) <= 1; flappy_W(12, 308) <= 1; flappy_W(12, 309) <= 1; flappy_W(12, 310) <= 1; flappy_W(12, 311) <= 1; flappy_W(12, 312) <= 1; flappy_W(12, 313) <= 1; flappy_W(12, 314) <= 1; flappy_W(12, 315) <= 1; flappy_W(12, 316) <= 1; flappy_W(12, 317) <= 1; flappy_W(12, 318) <= 0; flappy_W(12, 319) <= 0; flappy_W(12, 320) <= 0; flappy_W(12, 321) <= 0; flappy_W(12, 322) <= 0; flappy_W(12, 323) <= 0; flappy_W(12, 324) <= 0; flappy_W(12, 325) <= 0; flappy_W(12, 326) <= 0; flappy_W(12, 327) <= 0; flappy_W(12, 328) <= 0; flappy_W(12, 329) <= 0; flappy_W(12, 330) <= 0; flappy_W(12, 331) <= 0; flappy_W(12, 332) <= 0; flappy_W(12, 333) <= 0; flappy_W(12, 334) <= 0; flappy_W(12, 335) <= 0; flappy_W(12, 336) <= 0; flappy_W(12, 337) <= 0; flappy_W(12, 338) <= 0; flappy_W(12, 339) <= 0; flappy_W(12, 340) <= 0; flappy_W(12, 341) <= 0; flappy_W(12, 342) <= 0; flappy_W(12, 343) <= 0; flappy_W(12, 344) <= 0; flappy_W(12, 345) <= 0; flappy_W(12, 346) <= 0; flappy_W(12, 347) <= 0; flappy_W(12, 348) <= 0; flappy_W(12, 349) <= 0; flappy_W(12, 350) <= 0; flappy_W(12, 351) <= 0; flappy_W(12, 352) <= 0; flappy_W(12, 353) <= 0; flappy_W(12, 354) <= 0; flappy_W(12, 355) <= 0; flappy_W(12, 356) <= 0; flappy_W(12, 357) <= 0; flappy_W(12, 358) <= 0; flappy_W(12, 359) <= 0; flappy_W(12, 360) <= 0; flappy_W(12, 361) <= 0; flappy_W(12, 362) <= 0; flappy_W(12, 363) <= 0; flappy_W(12, 364) <= 0; flappy_W(12, 365) <= 0; flappy_W(12, 366) <= 0; flappy_W(12, 367) <= 0; flappy_W(12, 368) <= 0; flappy_W(12, 369) <= 0; flappy_W(12, 370) <= 0; flappy_W(12, 371) <= 0; flappy_W(12, 372) <= 0; flappy_W(12, 373) <= 0; flappy_W(12, 374) <= 0; flappy_W(12, 375) <= 0; flappy_W(12, 376) <= 0; flappy_W(12, 377) <= 0; flappy_W(12, 378) <= 0; flappy_W(12, 379) <= 0; flappy_W(12, 380) <= 0; flappy_W(12, 381) <= 0; flappy_W(12, 382) <= 0; flappy_W(12, 383) <= 0; flappy_W(12, 384) <= 0; flappy_W(12, 385) <= 0; flappy_W(12, 386) <= 0; flappy_W(12, 387) <= 0; flappy_W(12, 388) <= 0; flappy_W(12, 389) <= 0; flappy_W(12, 390) <= 0; flappy_W(12, 391) <= 0; flappy_W(12, 392) <= 0; flappy_W(12, 393) <= 0; flappy_W(12, 394) <= 0; flappy_W(12, 395) <= 0; flappy_W(12, 396) <= 0; flappy_W(12, 397) <= 0; flappy_W(12, 398) <= 0; flappy_W(12, 399) <= 0; flappy_W(12, 400) <= 0; flappy_W(12, 401) <= 0; flappy_W(12, 402) <= 1; flappy_W(12, 403) <= 1; flappy_W(12, 404) <= 1; flappy_W(12, 405) <= 1; flappy_W(12, 406) <= 1; flappy_W(12, 407) <= 1; flappy_W(12, 408) <= 1; flappy_W(12, 409) <= 1; flappy_W(12, 410) <= 1; flappy_W(12, 411) <= 1; flappy_W(12, 412) <= 1; flappy_W(12, 413) <= 1; flappy_W(12, 414) <= 0; flappy_W(12, 415) <= 0; flappy_W(12, 416) <= 0; flappy_W(12, 417) <= 0; flappy_W(12, 418) <= 0; flappy_W(12, 419) <= 0; flappy_W(12, 420) <= 0; flappy_W(12, 421) <= 0; flappy_W(12, 422) <= 0; flappy_W(12, 423) <= 0; flappy_W(12, 424) <= 0; flappy_W(12, 425) <= 0; flappy_W(12, 426) <= 1; flappy_W(12, 427) <= 1; flappy_W(12, 428) <= 1; flappy_W(12, 429) <= 1; flappy_W(12, 430) <= 1; flappy_W(12, 431) <= 1; flappy_W(12, 432) <= 1; flappy_W(12, 433) <= 1; flappy_W(12, 434) <= 1; flappy_W(12, 435) <= 1; flappy_W(12, 436) <= 1; flappy_W(12, 437) <= 1; flappy_W(12, 438) <= 0; flappy_W(12, 439) <= 0; flappy_W(12, 440) <= 0; flappy_W(12, 441) <= 0; flappy_W(12, 442) <= 0; flappy_W(12, 443) <= 0; flappy_W(12, 444) <= 0; flappy_W(12, 445) <= 0; flappy_W(12, 446) <= 0; flappy_W(12, 447) <= 0; flappy_W(12, 448) <= 0; flappy_W(12, 449) <= 0; flappy_W(12, 450) <= 0; flappy_W(12, 451) <= 0; flappy_W(12, 452) <= 0; flappy_W(12, 453) <= 0; flappy_W(12, 454) <= 0; flappy_W(12, 455) <= 0; flappy_W(12, 456) <= 0; flappy_W(12, 457) <= 0; flappy_W(12, 458) <= 0; flappy_W(12, 459) <= 0; flappy_W(12, 460) <= 0; flappy_W(12, 461) <= 0; flappy_W(12, 462) <= 0; flappy_W(12, 463) <= 0; flappy_W(12, 464) <= 0; flappy_W(12, 465) <= 0; flappy_W(12, 466) <= 0; flappy_W(12, 467) <= 0; flappy_W(12, 468) <= 1; flappy_W(12, 469) <= 1; flappy_W(12, 470) <= 1; flappy_W(12, 471) <= 1; flappy_W(12, 472) <= 1; flappy_W(12, 473) <= 1; flappy_W(12, 474) <= 1; flappy_W(12, 475) <= 1; flappy_W(12, 476) <= 1; flappy_W(12, 477) <= 1; flappy_W(12, 478) <= 1; flappy_W(12, 479) <= 1; flappy_W(12, 480) <= 0; flappy_W(12, 481) <= 0; flappy_W(12, 482) <= 0; flappy_W(12, 483) <= 0; flappy_W(12, 484) <= 0; flappy_W(12, 485) <= 0; flappy_W(12, 486) <= 0; flappy_W(12, 487) <= 0; flappy_W(12, 488) <= 0; flappy_W(12, 489) <= 0; flappy_W(12, 490) <= 0; flappy_W(12, 491) <= 0; flappy_W(12, 492) <= 0; flappy_W(12, 493) <= 0; flappy_W(12, 494) <= 0; flappy_W(12, 495) <= 0; flappy_W(12, 496) <= 0; flappy_W(12, 497) <= 0; flappy_W(12, 498) <= 0; flappy_W(12, 499) <= 0; flappy_W(12, 500) <= 0; flappy_W(12, 501) <= 0; flappy_W(12, 502) <= 0; flappy_W(12, 503) <= 0; flappy_W(12, 504) <= 0; flappy_W(12, 505) <= 0; flappy_W(12, 506) <= 0; flappy_W(12, 507) <= 0; flappy_W(12, 508) <= 0; flappy_W(12, 509) <= 0; flappy_W(12, 510) <= 1; flappy_W(12, 511) <= 1; flappy_W(12, 512) <= 1; flappy_W(12, 513) <= 1; flappy_W(12, 514) <= 1; flappy_W(12, 515) <= 1; flappy_W(12, 516) <= 1; flappy_W(12, 517) <= 1; flappy_W(12, 518) <= 1; flappy_W(12, 519) <= 1; flappy_W(12, 520) <= 1; flappy_W(12, 521) <= 1; flappy_W(12, 522) <= 0; flappy_W(12, 523) <= 0; flappy_W(12, 524) <= 0; flappy_W(12, 525) <= 0; flappy_W(12, 526) <= 0; flappy_W(12, 527) <= 0; flappy_W(12, 528) <= 0; flappy_W(12, 529) <= 0; flappy_W(12, 530) <= 0; flappy_W(12, 531) <= 0; flappy_W(12, 532) <= 0; flappy_W(12, 533) <= 0; flappy_W(12, 534) <= 1; flappy_W(12, 535) <= 1; flappy_W(12, 536) <= 1; flappy_W(12, 537) <= 1; flappy_W(12, 538) <= 1; flappy_W(12, 539) <= 1; flappy_W(12, 540) <= 1; flappy_W(12, 541) <= 1; flappy_W(12, 542) <= 1; flappy_W(12, 543) <= 1; flappy_W(12, 544) <= 1; flappy_W(12, 545) <= 1; flappy_W(12, 546) <= 0; flappy_W(12, 547) <= 0; flappy_W(12, 548) <= 0; flappy_W(12, 549) <= 0; flappy_W(12, 550) <= 0; flappy_W(12, 551) <= 0; flappy_W(12, 552) <= 0; flappy_W(12, 553) <= 0; flappy_W(12, 554) <= 0; flappy_W(12, 555) <= 0; flappy_W(12, 556) <= 0; flappy_W(12, 557) <= 0; flappy_W(12, 558) <= 0; flappy_W(12, 559) <= 0; flappy_W(12, 560) <= 0; flappy_W(12, 561) <= 0; flappy_W(12, 562) <= 0; flappy_W(12, 563) <= 0; flappy_W(12, 564) <= 1; flappy_W(12, 565) <= 1; flappy_W(12, 566) <= 1; flappy_W(12, 567) <= 1; flappy_W(12, 568) <= 1; flappy_W(12, 569) <= 1; flappy_W(12, 570) <= 1; flappy_W(12, 571) <= 1; flappy_W(12, 572) <= 1; flappy_W(12, 573) <= 1; flappy_W(12, 574) <= 1; flappy_W(12, 575) <= 1; flappy_W(12, 576) <= 0; flappy_W(12, 577) <= 0; flappy_W(12, 578) <= 0; flappy_W(12, 579) <= 0; flappy_W(12, 580) <= 0; flappy_W(12, 581) <= 0; flappy_W(12, 582) <= 0; flappy_W(12, 583) <= 0; flappy_W(12, 584) <= 0; flappy_W(12, 585) <= 0; flappy_W(12, 586) <= 0; flappy_W(12, 587) <= 0; flappy_W(12, 588) <= 1; flappy_W(12, 589) <= 1; flappy_W(12, 590) <= 1; flappy_W(12, 591) <= 1; flappy_W(12, 592) <= 1; flappy_W(12, 593) <= 1; 
flappy_W(13, 0) <= 0; flappy_W(13, 1) <= 0; flappy_W(13, 2) <= 0; flappy_W(13, 3) <= 0; flappy_W(13, 4) <= 0; flappy_W(13, 5) <= 0; flappy_W(13, 6) <= 1; flappy_W(13, 7) <= 1; flappy_W(13, 8) <= 1; flappy_W(13, 9) <= 1; flappy_W(13, 10) <= 1; flappy_W(13, 11) <= 1; flappy_W(13, 12) <= 1; flappy_W(13, 13) <= 1; flappy_W(13, 14) <= 1; flappy_W(13, 15) <= 1; flappy_W(13, 16) <= 1; flappy_W(13, 17) <= 1; flappy_W(13, 18) <= 0; flappy_W(13, 19) <= 0; flappy_W(13, 20) <= 0; flappy_W(13, 21) <= 0; flappy_W(13, 22) <= 0; flappy_W(13, 23) <= 0; flappy_W(13, 24) <= 0; flappy_W(13, 25) <= 0; flappy_W(13, 26) <= 0; flappy_W(13, 27) <= 0; flappy_W(13, 28) <= 0; flappy_W(13, 29) <= 0; flappy_W(13, 30) <= 0; flappy_W(13, 31) <= 0; flappy_W(13, 32) <= 0; flappy_W(13, 33) <= 0; flappy_W(13, 34) <= 0; flappy_W(13, 35) <= 0; flappy_W(13, 36) <= 1; flappy_W(13, 37) <= 1; flappy_W(13, 38) <= 1; flappy_W(13, 39) <= 1; flappy_W(13, 40) <= 1; flappy_W(13, 41) <= 1; flappy_W(13, 42) <= 0; flappy_W(13, 43) <= 0; flappy_W(13, 44) <= 0; flappy_W(13, 45) <= 0; flappy_W(13, 46) <= 0; flappy_W(13, 47) <= 0; flappy_W(13, 48) <= 0; flappy_W(13, 49) <= 0; flappy_W(13, 50) <= 0; flappy_W(13, 51) <= 0; flappy_W(13, 52) <= 0; flappy_W(13, 53) <= 0; flappy_W(13, 54) <= 0; flappy_W(13, 55) <= 0; flappy_W(13, 56) <= 0; flappy_W(13, 57) <= 0; flappy_W(13, 58) <= 0; flappy_W(13, 59) <= 0; flappy_W(13, 60) <= 1; flappy_W(13, 61) <= 1; flappy_W(13, 62) <= 1; flappy_W(13, 63) <= 1; flappy_W(13, 64) <= 1; flappy_W(13, 65) <= 1; flappy_W(13, 66) <= 1; flappy_W(13, 67) <= 1; flappy_W(13, 68) <= 1; flappy_W(13, 69) <= 1; flappy_W(13, 70) <= 1; flappy_W(13, 71) <= 1; flappy_W(13, 72) <= 0; flappy_W(13, 73) <= 0; flappy_W(13, 74) <= 0; flappy_W(13, 75) <= 0; flappy_W(13, 76) <= 0; flappy_W(13, 77) <= 0; flappy_W(13, 78) <= 0; flappy_W(13, 79) <= 0; flappy_W(13, 80) <= 0; flappy_W(13, 81) <= 0; flappy_W(13, 82) <= 0; flappy_W(13, 83) <= 0; flappy_W(13, 84) <= 0; flappy_W(13, 85) <= 0; flappy_W(13, 86) <= 0; flappy_W(13, 87) <= 0; flappy_W(13, 88) <= 0; flappy_W(13, 89) <= 0; flappy_W(13, 90) <= 0; flappy_W(13, 91) <= 0; flappy_W(13, 92) <= 0; flappy_W(13, 93) <= 0; flappy_W(13, 94) <= 0; flappy_W(13, 95) <= 0; flappy_W(13, 96) <= 0; flappy_W(13, 97) <= 0; flappy_W(13, 98) <= 0; flappy_W(13, 99) <= 0; flappy_W(13, 100) <= 0; flappy_W(13, 101) <= 0; flappy_W(13, 102) <= 0; flappy_W(13, 103) <= 0; flappy_W(13, 104) <= 0; flappy_W(13, 105) <= 0; flappy_W(13, 106) <= 0; flappy_W(13, 107) <= 0; flappy_W(13, 108) <= 0; flappy_W(13, 109) <= 0; flappy_W(13, 110) <= 0; flappy_W(13, 111) <= 0; flappy_W(13, 112) <= 0; flappy_W(13, 113) <= 0; flappy_W(13, 114) <= 1; flappy_W(13, 115) <= 1; flappy_W(13, 116) <= 1; flappy_W(13, 117) <= 1; flappy_W(13, 118) <= 1; flappy_W(13, 119) <= 1; flappy_W(13, 120) <= 1; flappy_W(13, 121) <= 1; flappy_W(13, 122) <= 1; flappy_W(13, 123) <= 1; flappy_W(13, 124) <= 1; flappy_W(13, 125) <= 1; flappy_W(13, 126) <= 0; flappy_W(13, 127) <= 0; flappy_W(13, 128) <= 0; flappy_W(13, 129) <= 0; flappy_W(13, 130) <= 0; flappy_W(13, 131) <= 0; flappy_W(13, 132) <= 1; flappy_W(13, 133) <= 1; flappy_W(13, 134) <= 1; flappy_W(13, 135) <= 1; flappy_W(13, 136) <= 1; flappy_W(13, 137) <= 1; flappy_W(13, 138) <= 1; flappy_W(13, 139) <= 1; flappy_W(13, 140) <= 1; flappy_W(13, 141) <= 1; flappy_W(13, 142) <= 1; flappy_W(13, 143) <= 1; flappy_W(13, 144) <= 0; flappy_W(13, 145) <= 0; flappy_W(13, 146) <= 0; flappy_W(13, 147) <= 0; flappy_W(13, 148) <= 0; flappy_W(13, 149) <= 0; flappy_W(13, 150) <= 0; flappy_W(13, 151) <= 0; flappy_W(13, 152) <= 0; flappy_W(13, 153) <= 0; flappy_W(13, 154) <= 0; flappy_W(13, 155) <= 0; flappy_W(13, 156) <= 0; flappy_W(13, 157) <= 0; flappy_W(13, 158) <= 0; flappy_W(13, 159) <= 0; flappy_W(13, 160) <= 0; flappy_W(13, 161) <= 0; flappy_W(13, 162) <= 0; flappy_W(13, 163) <= 0; flappy_W(13, 164) <= 0; flappy_W(13, 165) <= 0; flappy_W(13, 166) <= 0; flappy_W(13, 167) <= 0; flappy_W(13, 168) <= 1; flappy_W(13, 169) <= 1; flappy_W(13, 170) <= 1; flappy_W(13, 171) <= 1; flappy_W(13, 172) <= 1; flappy_W(13, 173) <= 1; flappy_W(13, 174) <= 1; flappy_W(13, 175) <= 1; flappy_W(13, 176) <= 1; flappy_W(13, 177) <= 1; flappy_W(13, 178) <= 1; flappy_W(13, 179) <= 1; flappy_W(13, 180) <= 0; flappy_W(13, 181) <= 0; flappy_W(13, 182) <= 0; flappy_W(13, 183) <= 0; flappy_W(13, 184) <= 0; flappy_W(13, 185) <= 0; flappy_W(13, 186) <= 0; flappy_W(13, 187) <= 0; flappy_W(13, 188) <= 0; flappy_W(13, 189) <= 0; flappy_W(13, 190) <= 0; flappy_W(13, 191) <= 0; flappy_W(13, 192) <= 1; flappy_W(13, 193) <= 1; flappy_W(13, 194) <= 1; flappy_W(13, 195) <= 1; flappy_W(13, 196) <= 1; flappy_W(13, 197) <= 1; flappy_W(13, 198) <= 1; flappy_W(13, 199) <= 1; flappy_W(13, 200) <= 1; flappy_W(13, 201) <= 1; flappy_W(13, 202) <= 1; flappy_W(13, 203) <= 1; flappy_W(13, 204) <= 0; flappy_W(13, 205) <= 0; flappy_W(13, 206) <= 0; flappy_W(13, 207) <= 0; flappy_W(13, 208) <= 0; flappy_W(13, 209) <= 0; flappy_W(13, 210) <= 0; flappy_W(13, 211) <= 0; flappy_W(13, 212) <= 0; flappy_W(13, 213) <= 0; flappy_W(13, 214) <= 0; flappy_W(13, 215) <= 0; flappy_W(13, 216) <= 0; flappy_W(13, 217) <= 0; flappy_W(13, 218) <= 0; flappy_W(13, 219) <= 0; flappy_W(13, 220) <= 0; flappy_W(13, 221) <= 0; flappy_W(13, 222) <= 1; flappy_W(13, 223) <= 1; flappy_W(13, 224) <= 1; flappy_W(13, 225) <= 1; flappy_W(13, 226) <= 1; flappy_W(13, 227) <= 1; flappy_W(13, 228) <= 1; flappy_W(13, 229) <= 1; flappy_W(13, 230) <= 1; flappy_W(13, 231) <= 1; flappy_W(13, 232) <= 1; flappy_W(13, 233) <= 1; flappy_W(13, 234) <= 0; flappy_W(13, 235) <= 0; flappy_W(13, 236) <= 0; flappy_W(13, 237) <= 0; flappy_W(13, 238) <= 0; flappy_W(13, 239) <= 0; flappy_W(13, 240) <= 0; flappy_W(13, 241) <= 0; flappy_W(13, 242) <= 0; flappy_W(13, 243) <= 0; flappy_W(13, 244) <= 0; flappy_W(13, 245) <= 0; flappy_W(13, 246) <= 1; flappy_W(13, 247) <= 1; flappy_W(13, 248) <= 1; flappy_W(13, 249) <= 1; flappy_W(13, 250) <= 1; flappy_W(13, 251) <= 1; flappy_W(13, 252) <= 1; flappy_W(13, 253) <= 1; flappy_W(13, 254) <= 1; flappy_W(13, 255) <= 1; flappy_W(13, 256) <= 1; flappy_W(13, 257) <= 1; flappy_W(13, 258) <= 0; flappy_W(13, 259) <= 0; flappy_W(13, 260) <= 0; flappy_W(13, 261) <= 0; flappy_W(13, 262) <= 0; flappy_W(13, 263) <= 0; flappy_W(13, 264) <= 0; flappy_W(13, 265) <= 0; flappy_W(13, 266) <= 0; flappy_W(13, 267) <= 0; flappy_W(13, 268) <= 0; flappy_W(13, 269) <= 0; flappy_W(13, 270) <= 1; flappy_W(13, 271) <= 1; flappy_W(13, 272) <= 1; flappy_W(13, 273) <= 1; flappy_W(13, 274) <= 1; flappy_W(13, 275) <= 1; flappy_W(13, 276) <= 1; flappy_W(13, 277) <= 1; flappy_W(13, 278) <= 1; flappy_W(13, 279) <= 1; flappy_W(13, 280) <= 1; flappy_W(13, 281) <= 1; flappy_W(13, 282) <= 0; flappy_W(13, 283) <= 0; flappy_W(13, 284) <= 0; flappy_W(13, 285) <= 0; flappy_W(13, 286) <= 0; flappy_W(13, 287) <= 0; flappy_W(13, 288) <= 0; flappy_W(13, 289) <= 0; flappy_W(13, 290) <= 0; flappy_W(13, 291) <= 0; flappy_W(13, 292) <= 0; flappy_W(13, 293) <= 0; flappy_W(13, 294) <= 0; flappy_W(13, 295) <= 0; flappy_W(13, 296) <= 0; flappy_W(13, 297) <= 0; flappy_W(13, 298) <= 0; flappy_W(13, 299) <= 0; flappy_W(13, 300) <= 0; flappy_W(13, 301) <= 0; flappy_W(13, 302) <= 0; flappy_W(13, 303) <= 0; flappy_W(13, 304) <= 0; flappy_W(13, 305) <= 0; flappy_W(13, 306) <= 1; flappy_W(13, 307) <= 1; flappy_W(13, 308) <= 1; flappy_W(13, 309) <= 1; flappy_W(13, 310) <= 1; flappy_W(13, 311) <= 1; flappy_W(13, 312) <= 1; flappy_W(13, 313) <= 1; flappy_W(13, 314) <= 1; flappy_W(13, 315) <= 1; flappy_W(13, 316) <= 1; flappy_W(13, 317) <= 1; flappy_W(13, 318) <= 0; flappy_W(13, 319) <= 0; flappy_W(13, 320) <= 0; flappy_W(13, 321) <= 0; flappy_W(13, 322) <= 0; flappy_W(13, 323) <= 0; flappy_W(13, 324) <= 0; flappy_W(13, 325) <= 0; flappy_W(13, 326) <= 0; flappy_W(13, 327) <= 0; flappy_W(13, 328) <= 0; flappy_W(13, 329) <= 0; flappy_W(13, 330) <= 0; flappy_W(13, 331) <= 0; flappy_W(13, 332) <= 0; flappy_W(13, 333) <= 0; flappy_W(13, 334) <= 0; flappy_W(13, 335) <= 0; flappy_W(13, 336) <= 0; flappy_W(13, 337) <= 0; flappy_W(13, 338) <= 0; flappy_W(13, 339) <= 0; flappy_W(13, 340) <= 0; flappy_W(13, 341) <= 0; flappy_W(13, 342) <= 0; flappy_W(13, 343) <= 0; flappy_W(13, 344) <= 0; flappy_W(13, 345) <= 0; flappy_W(13, 346) <= 0; flappy_W(13, 347) <= 0; flappy_W(13, 348) <= 0; flappy_W(13, 349) <= 0; flappy_W(13, 350) <= 0; flappy_W(13, 351) <= 0; flappy_W(13, 352) <= 0; flappy_W(13, 353) <= 0; flappy_W(13, 354) <= 0; flappy_W(13, 355) <= 0; flappy_W(13, 356) <= 0; flappy_W(13, 357) <= 0; flappy_W(13, 358) <= 0; flappy_W(13, 359) <= 0; flappy_W(13, 360) <= 0; flappy_W(13, 361) <= 0; flappy_W(13, 362) <= 0; flappy_W(13, 363) <= 0; flappy_W(13, 364) <= 0; flappy_W(13, 365) <= 0; flappy_W(13, 366) <= 0; flappy_W(13, 367) <= 0; flappy_W(13, 368) <= 0; flappy_W(13, 369) <= 0; flappy_W(13, 370) <= 0; flappy_W(13, 371) <= 0; flappy_W(13, 372) <= 0; flappy_W(13, 373) <= 0; flappy_W(13, 374) <= 0; flappy_W(13, 375) <= 0; flappy_W(13, 376) <= 0; flappy_W(13, 377) <= 0; flappy_W(13, 378) <= 0; flappy_W(13, 379) <= 0; flappy_W(13, 380) <= 0; flappy_W(13, 381) <= 0; flappy_W(13, 382) <= 0; flappy_W(13, 383) <= 0; flappy_W(13, 384) <= 0; flappy_W(13, 385) <= 0; flappy_W(13, 386) <= 0; flappy_W(13, 387) <= 0; flappy_W(13, 388) <= 0; flappy_W(13, 389) <= 0; flappy_W(13, 390) <= 0; flappy_W(13, 391) <= 0; flappy_W(13, 392) <= 0; flappy_W(13, 393) <= 0; flappy_W(13, 394) <= 0; flappy_W(13, 395) <= 0; flappy_W(13, 396) <= 0; flappy_W(13, 397) <= 0; flappy_W(13, 398) <= 0; flappy_W(13, 399) <= 0; flappy_W(13, 400) <= 0; flappy_W(13, 401) <= 0; flappy_W(13, 402) <= 1; flappy_W(13, 403) <= 1; flappy_W(13, 404) <= 1; flappy_W(13, 405) <= 1; flappy_W(13, 406) <= 1; flappy_W(13, 407) <= 1; flappy_W(13, 408) <= 1; flappy_W(13, 409) <= 1; flappy_W(13, 410) <= 1; flappy_W(13, 411) <= 1; flappy_W(13, 412) <= 1; flappy_W(13, 413) <= 1; flappy_W(13, 414) <= 0; flappy_W(13, 415) <= 0; flappy_W(13, 416) <= 0; flappy_W(13, 417) <= 0; flappy_W(13, 418) <= 0; flappy_W(13, 419) <= 0; flappy_W(13, 420) <= 0; flappy_W(13, 421) <= 0; flappy_W(13, 422) <= 0; flappy_W(13, 423) <= 0; flappy_W(13, 424) <= 0; flappy_W(13, 425) <= 0; flappy_W(13, 426) <= 1; flappy_W(13, 427) <= 1; flappy_W(13, 428) <= 1; flappy_W(13, 429) <= 1; flappy_W(13, 430) <= 1; flappy_W(13, 431) <= 1; flappy_W(13, 432) <= 1; flappy_W(13, 433) <= 1; flappy_W(13, 434) <= 1; flappy_W(13, 435) <= 1; flappy_W(13, 436) <= 1; flappy_W(13, 437) <= 1; flappy_W(13, 438) <= 0; flappy_W(13, 439) <= 0; flappy_W(13, 440) <= 0; flappy_W(13, 441) <= 0; flappy_W(13, 442) <= 0; flappy_W(13, 443) <= 0; flappy_W(13, 444) <= 0; flappy_W(13, 445) <= 0; flappy_W(13, 446) <= 0; flappy_W(13, 447) <= 0; flappy_W(13, 448) <= 0; flappy_W(13, 449) <= 0; flappy_W(13, 450) <= 0; flappy_W(13, 451) <= 0; flappy_W(13, 452) <= 0; flappy_W(13, 453) <= 0; flappy_W(13, 454) <= 0; flappy_W(13, 455) <= 0; flappy_W(13, 456) <= 0; flappy_W(13, 457) <= 0; flappy_W(13, 458) <= 0; flappy_W(13, 459) <= 0; flappy_W(13, 460) <= 0; flappy_W(13, 461) <= 0; flappy_W(13, 462) <= 0; flappy_W(13, 463) <= 0; flappy_W(13, 464) <= 0; flappy_W(13, 465) <= 0; flappy_W(13, 466) <= 0; flappy_W(13, 467) <= 0; flappy_W(13, 468) <= 1; flappy_W(13, 469) <= 1; flappy_W(13, 470) <= 1; flappy_W(13, 471) <= 1; flappy_W(13, 472) <= 1; flappy_W(13, 473) <= 1; flappy_W(13, 474) <= 1; flappy_W(13, 475) <= 1; flappy_W(13, 476) <= 1; flappy_W(13, 477) <= 1; flappy_W(13, 478) <= 1; flappy_W(13, 479) <= 1; flappy_W(13, 480) <= 0; flappy_W(13, 481) <= 0; flappy_W(13, 482) <= 0; flappy_W(13, 483) <= 0; flappy_W(13, 484) <= 0; flappy_W(13, 485) <= 0; flappy_W(13, 486) <= 0; flappy_W(13, 487) <= 0; flappy_W(13, 488) <= 0; flappy_W(13, 489) <= 0; flappy_W(13, 490) <= 0; flappy_W(13, 491) <= 0; flappy_W(13, 492) <= 0; flappy_W(13, 493) <= 0; flappy_W(13, 494) <= 0; flappy_W(13, 495) <= 0; flappy_W(13, 496) <= 0; flappy_W(13, 497) <= 0; flappy_W(13, 498) <= 0; flappy_W(13, 499) <= 0; flappy_W(13, 500) <= 0; flappy_W(13, 501) <= 0; flappy_W(13, 502) <= 0; flappy_W(13, 503) <= 0; flappy_W(13, 504) <= 0; flappy_W(13, 505) <= 0; flappy_W(13, 506) <= 0; flappy_W(13, 507) <= 0; flappy_W(13, 508) <= 0; flappy_W(13, 509) <= 0; flappy_W(13, 510) <= 1; flappy_W(13, 511) <= 1; flappy_W(13, 512) <= 1; flappy_W(13, 513) <= 1; flappy_W(13, 514) <= 1; flappy_W(13, 515) <= 1; flappy_W(13, 516) <= 1; flappy_W(13, 517) <= 1; flappy_W(13, 518) <= 1; flappy_W(13, 519) <= 1; flappy_W(13, 520) <= 1; flappy_W(13, 521) <= 1; flappy_W(13, 522) <= 0; flappy_W(13, 523) <= 0; flappy_W(13, 524) <= 0; flappy_W(13, 525) <= 0; flappy_W(13, 526) <= 0; flappy_W(13, 527) <= 0; flappy_W(13, 528) <= 0; flappy_W(13, 529) <= 0; flappy_W(13, 530) <= 0; flappy_W(13, 531) <= 0; flappy_W(13, 532) <= 0; flappy_W(13, 533) <= 0; flappy_W(13, 534) <= 1; flappy_W(13, 535) <= 1; flappy_W(13, 536) <= 1; flappy_W(13, 537) <= 1; flappy_W(13, 538) <= 1; flappy_W(13, 539) <= 1; flappy_W(13, 540) <= 1; flappy_W(13, 541) <= 1; flappy_W(13, 542) <= 1; flappy_W(13, 543) <= 1; flappy_W(13, 544) <= 1; flappy_W(13, 545) <= 1; flappy_W(13, 546) <= 0; flappy_W(13, 547) <= 0; flappy_W(13, 548) <= 0; flappy_W(13, 549) <= 0; flappy_W(13, 550) <= 0; flappy_W(13, 551) <= 0; flappy_W(13, 552) <= 0; flappy_W(13, 553) <= 0; flappy_W(13, 554) <= 0; flappy_W(13, 555) <= 0; flappy_W(13, 556) <= 0; flappy_W(13, 557) <= 0; flappy_W(13, 558) <= 0; flappy_W(13, 559) <= 0; flappy_W(13, 560) <= 0; flappy_W(13, 561) <= 0; flappy_W(13, 562) <= 0; flappy_W(13, 563) <= 0; flappy_W(13, 564) <= 1; flappy_W(13, 565) <= 1; flappy_W(13, 566) <= 1; flappy_W(13, 567) <= 1; flappy_W(13, 568) <= 1; flappy_W(13, 569) <= 1; flappy_W(13, 570) <= 1; flappy_W(13, 571) <= 1; flappy_W(13, 572) <= 1; flappy_W(13, 573) <= 1; flappy_W(13, 574) <= 1; flappy_W(13, 575) <= 1; flappy_W(13, 576) <= 0; flappy_W(13, 577) <= 0; flappy_W(13, 578) <= 0; flappy_W(13, 579) <= 0; flappy_W(13, 580) <= 0; flappy_W(13, 581) <= 0; flappy_W(13, 582) <= 0; flappy_W(13, 583) <= 0; flappy_W(13, 584) <= 0; flappy_W(13, 585) <= 0; flappy_W(13, 586) <= 0; flappy_W(13, 587) <= 0; flappy_W(13, 588) <= 1; flappy_W(13, 589) <= 1; flappy_W(13, 590) <= 1; flappy_W(13, 591) <= 1; flappy_W(13, 592) <= 1; flappy_W(13, 593) <= 1; 
flappy_W(14, 0) <= 0; flappy_W(14, 1) <= 0; flappy_W(14, 2) <= 0; flappy_W(14, 3) <= 0; flappy_W(14, 4) <= 0; flappy_W(14, 5) <= 0; flappy_W(14, 6) <= 1; flappy_W(14, 7) <= 1; flappy_W(14, 8) <= 1; flappy_W(14, 9) <= 1; flappy_W(14, 10) <= 1; flappy_W(14, 11) <= 1; flappy_W(14, 12) <= 1; flappy_W(14, 13) <= 1; flappy_W(14, 14) <= 1; flappy_W(14, 15) <= 1; flappy_W(14, 16) <= 1; flappy_W(14, 17) <= 1; flappy_W(14, 18) <= 0; flappy_W(14, 19) <= 0; flappy_W(14, 20) <= 0; flappy_W(14, 21) <= 0; flappy_W(14, 22) <= 0; flappy_W(14, 23) <= 0; flappy_W(14, 24) <= 0; flappy_W(14, 25) <= 0; flappy_W(14, 26) <= 0; flappy_W(14, 27) <= 0; flappy_W(14, 28) <= 0; flappy_W(14, 29) <= 0; flappy_W(14, 30) <= 0; flappy_W(14, 31) <= 0; flappy_W(14, 32) <= 0; flappy_W(14, 33) <= 0; flappy_W(14, 34) <= 0; flappy_W(14, 35) <= 0; flappy_W(14, 36) <= 1; flappy_W(14, 37) <= 1; flappy_W(14, 38) <= 1; flappy_W(14, 39) <= 1; flappy_W(14, 40) <= 1; flappy_W(14, 41) <= 1; flappy_W(14, 42) <= 0; flappy_W(14, 43) <= 0; flappy_W(14, 44) <= 0; flappy_W(14, 45) <= 0; flappy_W(14, 46) <= 0; flappy_W(14, 47) <= 0; flappy_W(14, 48) <= 0; flappy_W(14, 49) <= 0; flappy_W(14, 50) <= 0; flappy_W(14, 51) <= 0; flappy_W(14, 52) <= 0; flappy_W(14, 53) <= 0; flappy_W(14, 54) <= 0; flappy_W(14, 55) <= 0; flappy_W(14, 56) <= 0; flappy_W(14, 57) <= 0; flappy_W(14, 58) <= 0; flappy_W(14, 59) <= 0; flappy_W(14, 60) <= 1; flappy_W(14, 61) <= 1; flappy_W(14, 62) <= 1; flappy_W(14, 63) <= 1; flappy_W(14, 64) <= 1; flappy_W(14, 65) <= 1; flappy_W(14, 66) <= 1; flappy_W(14, 67) <= 1; flappy_W(14, 68) <= 1; flappy_W(14, 69) <= 1; flappy_W(14, 70) <= 1; flappy_W(14, 71) <= 1; flappy_W(14, 72) <= 0; flappy_W(14, 73) <= 0; flappy_W(14, 74) <= 0; flappy_W(14, 75) <= 0; flappy_W(14, 76) <= 0; flappy_W(14, 77) <= 0; flappy_W(14, 78) <= 0; flappy_W(14, 79) <= 0; flappy_W(14, 80) <= 0; flappy_W(14, 81) <= 0; flappy_W(14, 82) <= 0; flappy_W(14, 83) <= 0; flappy_W(14, 84) <= 0; flappy_W(14, 85) <= 0; flappy_W(14, 86) <= 0; flappy_W(14, 87) <= 0; flappy_W(14, 88) <= 0; flappy_W(14, 89) <= 0; flappy_W(14, 90) <= 0; flappy_W(14, 91) <= 0; flappy_W(14, 92) <= 0; flappy_W(14, 93) <= 0; flappy_W(14, 94) <= 0; flappy_W(14, 95) <= 0; flappy_W(14, 96) <= 0; flappy_W(14, 97) <= 0; flappy_W(14, 98) <= 0; flappy_W(14, 99) <= 0; flappy_W(14, 100) <= 0; flappy_W(14, 101) <= 0; flappy_W(14, 102) <= 0; flappy_W(14, 103) <= 0; flappy_W(14, 104) <= 0; flappy_W(14, 105) <= 0; flappy_W(14, 106) <= 0; flappy_W(14, 107) <= 0; flappy_W(14, 108) <= 0; flappy_W(14, 109) <= 0; flappy_W(14, 110) <= 0; flappy_W(14, 111) <= 0; flappy_W(14, 112) <= 0; flappy_W(14, 113) <= 0; flappy_W(14, 114) <= 1; flappy_W(14, 115) <= 1; flappy_W(14, 116) <= 1; flappy_W(14, 117) <= 1; flappy_W(14, 118) <= 1; flappy_W(14, 119) <= 1; flappy_W(14, 120) <= 1; flappy_W(14, 121) <= 1; flappy_W(14, 122) <= 1; flappy_W(14, 123) <= 1; flappy_W(14, 124) <= 1; flappy_W(14, 125) <= 1; flappy_W(14, 126) <= 0; flappy_W(14, 127) <= 0; flappy_W(14, 128) <= 0; flappy_W(14, 129) <= 0; flappy_W(14, 130) <= 0; flappy_W(14, 131) <= 0; flappy_W(14, 132) <= 1; flappy_W(14, 133) <= 1; flappy_W(14, 134) <= 1; flappy_W(14, 135) <= 1; flappy_W(14, 136) <= 1; flappy_W(14, 137) <= 1; flappy_W(14, 138) <= 1; flappy_W(14, 139) <= 1; flappy_W(14, 140) <= 1; flappy_W(14, 141) <= 1; flappy_W(14, 142) <= 1; flappy_W(14, 143) <= 1; flappy_W(14, 144) <= 0; flappy_W(14, 145) <= 0; flappy_W(14, 146) <= 0; flappy_W(14, 147) <= 0; flappy_W(14, 148) <= 0; flappy_W(14, 149) <= 0; flappy_W(14, 150) <= 0; flappy_W(14, 151) <= 0; flappy_W(14, 152) <= 0; flappy_W(14, 153) <= 0; flappy_W(14, 154) <= 0; flappy_W(14, 155) <= 0; flappy_W(14, 156) <= 0; flappy_W(14, 157) <= 0; flappy_W(14, 158) <= 0; flappy_W(14, 159) <= 0; flappy_W(14, 160) <= 0; flappy_W(14, 161) <= 0; flappy_W(14, 162) <= 0; flappy_W(14, 163) <= 0; flappy_W(14, 164) <= 0; flappy_W(14, 165) <= 0; flappy_W(14, 166) <= 0; flappy_W(14, 167) <= 0; flappy_W(14, 168) <= 1; flappy_W(14, 169) <= 1; flappy_W(14, 170) <= 1; flappy_W(14, 171) <= 1; flappy_W(14, 172) <= 1; flappy_W(14, 173) <= 1; flappy_W(14, 174) <= 1; flappy_W(14, 175) <= 1; flappy_W(14, 176) <= 1; flappy_W(14, 177) <= 1; flappy_W(14, 178) <= 1; flappy_W(14, 179) <= 1; flappy_W(14, 180) <= 0; flappy_W(14, 181) <= 0; flappy_W(14, 182) <= 0; flappy_W(14, 183) <= 0; flappy_W(14, 184) <= 0; flappy_W(14, 185) <= 0; flappy_W(14, 186) <= 0; flappy_W(14, 187) <= 0; flappy_W(14, 188) <= 0; flappy_W(14, 189) <= 0; flappy_W(14, 190) <= 0; flappy_W(14, 191) <= 0; flappy_W(14, 192) <= 1; flappy_W(14, 193) <= 1; flappy_W(14, 194) <= 1; flappy_W(14, 195) <= 1; flappy_W(14, 196) <= 1; flappy_W(14, 197) <= 1; flappy_W(14, 198) <= 1; flappy_W(14, 199) <= 1; flappy_W(14, 200) <= 1; flappy_W(14, 201) <= 1; flappy_W(14, 202) <= 1; flappy_W(14, 203) <= 1; flappy_W(14, 204) <= 0; flappy_W(14, 205) <= 0; flappy_W(14, 206) <= 0; flappy_W(14, 207) <= 0; flappy_W(14, 208) <= 0; flappy_W(14, 209) <= 0; flappy_W(14, 210) <= 0; flappy_W(14, 211) <= 0; flappy_W(14, 212) <= 0; flappy_W(14, 213) <= 0; flappy_W(14, 214) <= 0; flappy_W(14, 215) <= 0; flappy_W(14, 216) <= 0; flappy_W(14, 217) <= 0; flappy_W(14, 218) <= 0; flappy_W(14, 219) <= 0; flappy_W(14, 220) <= 0; flappy_W(14, 221) <= 0; flappy_W(14, 222) <= 1; flappy_W(14, 223) <= 1; flappy_W(14, 224) <= 1; flappy_W(14, 225) <= 1; flappy_W(14, 226) <= 1; flappy_W(14, 227) <= 1; flappy_W(14, 228) <= 1; flappy_W(14, 229) <= 1; flappy_W(14, 230) <= 1; flappy_W(14, 231) <= 1; flappy_W(14, 232) <= 1; flappy_W(14, 233) <= 1; flappy_W(14, 234) <= 0; flappy_W(14, 235) <= 0; flappy_W(14, 236) <= 0; flappy_W(14, 237) <= 0; flappy_W(14, 238) <= 0; flappy_W(14, 239) <= 0; flappy_W(14, 240) <= 0; flappy_W(14, 241) <= 0; flappy_W(14, 242) <= 0; flappy_W(14, 243) <= 0; flappy_W(14, 244) <= 0; flappy_W(14, 245) <= 0; flappy_W(14, 246) <= 1; flappy_W(14, 247) <= 1; flappy_W(14, 248) <= 1; flappy_W(14, 249) <= 1; flappy_W(14, 250) <= 1; flappy_W(14, 251) <= 1; flappy_W(14, 252) <= 1; flappy_W(14, 253) <= 1; flappy_W(14, 254) <= 1; flappy_W(14, 255) <= 1; flappy_W(14, 256) <= 1; flappy_W(14, 257) <= 1; flappy_W(14, 258) <= 0; flappy_W(14, 259) <= 0; flappy_W(14, 260) <= 0; flappy_W(14, 261) <= 0; flappy_W(14, 262) <= 0; flappy_W(14, 263) <= 0; flappy_W(14, 264) <= 0; flappy_W(14, 265) <= 0; flappy_W(14, 266) <= 0; flappy_W(14, 267) <= 0; flappy_W(14, 268) <= 0; flappy_W(14, 269) <= 0; flappy_W(14, 270) <= 1; flappy_W(14, 271) <= 1; flappy_W(14, 272) <= 1; flappy_W(14, 273) <= 1; flappy_W(14, 274) <= 1; flappy_W(14, 275) <= 1; flappy_W(14, 276) <= 1; flappy_W(14, 277) <= 1; flappy_W(14, 278) <= 1; flappy_W(14, 279) <= 1; flappy_W(14, 280) <= 1; flappy_W(14, 281) <= 1; flappy_W(14, 282) <= 0; flappy_W(14, 283) <= 0; flappy_W(14, 284) <= 0; flappy_W(14, 285) <= 0; flappy_W(14, 286) <= 0; flappy_W(14, 287) <= 0; flappy_W(14, 288) <= 0; flappy_W(14, 289) <= 0; flappy_W(14, 290) <= 0; flappy_W(14, 291) <= 0; flappy_W(14, 292) <= 0; flappy_W(14, 293) <= 0; flappy_W(14, 294) <= 0; flappy_W(14, 295) <= 0; flappy_W(14, 296) <= 0; flappy_W(14, 297) <= 0; flappy_W(14, 298) <= 0; flappy_W(14, 299) <= 0; flappy_W(14, 300) <= 0; flappy_W(14, 301) <= 0; flappy_W(14, 302) <= 0; flappy_W(14, 303) <= 0; flappy_W(14, 304) <= 0; flappy_W(14, 305) <= 0; flappy_W(14, 306) <= 1; flappy_W(14, 307) <= 1; flappy_W(14, 308) <= 1; flappy_W(14, 309) <= 1; flappy_W(14, 310) <= 1; flappy_W(14, 311) <= 1; flappy_W(14, 312) <= 1; flappy_W(14, 313) <= 1; flappy_W(14, 314) <= 1; flappy_W(14, 315) <= 1; flappy_W(14, 316) <= 1; flappy_W(14, 317) <= 1; flappy_W(14, 318) <= 0; flappy_W(14, 319) <= 0; flappy_W(14, 320) <= 0; flappy_W(14, 321) <= 0; flappy_W(14, 322) <= 0; flappy_W(14, 323) <= 0; flappy_W(14, 324) <= 0; flappy_W(14, 325) <= 0; flappy_W(14, 326) <= 0; flappy_W(14, 327) <= 0; flappy_W(14, 328) <= 0; flappy_W(14, 329) <= 0; flappy_W(14, 330) <= 0; flappy_W(14, 331) <= 0; flappy_W(14, 332) <= 0; flappy_W(14, 333) <= 0; flappy_W(14, 334) <= 0; flappy_W(14, 335) <= 0; flappy_W(14, 336) <= 0; flappy_W(14, 337) <= 0; flappy_W(14, 338) <= 0; flappy_W(14, 339) <= 0; flappy_W(14, 340) <= 0; flappy_W(14, 341) <= 0; flappy_W(14, 342) <= 0; flappy_W(14, 343) <= 0; flappy_W(14, 344) <= 0; flappy_W(14, 345) <= 0; flappy_W(14, 346) <= 0; flappy_W(14, 347) <= 0; flappy_W(14, 348) <= 0; flappy_W(14, 349) <= 0; flappy_W(14, 350) <= 0; flappy_W(14, 351) <= 0; flappy_W(14, 352) <= 0; flappy_W(14, 353) <= 0; flappy_W(14, 354) <= 0; flappy_W(14, 355) <= 0; flappy_W(14, 356) <= 0; flappy_W(14, 357) <= 0; flappy_W(14, 358) <= 0; flappy_W(14, 359) <= 0; flappy_W(14, 360) <= 0; flappy_W(14, 361) <= 0; flappy_W(14, 362) <= 0; flappy_W(14, 363) <= 0; flappy_W(14, 364) <= 0; flappy_W(14, 365) <= 0; flappy_W(14, 366) <= 0; flappy_W(14, 367) <= 0; flappy_W(14, 368) <= 0; flappy_W(14, 369) <= 0; flappy_W(14, 370) <= 0; flappy_W(14, 371) <= 0; flappy_W(14, 372) <= 0; flappy_W(14, 373) <= 0; flappy_W(14, 374) <= 0; flappy_W(14, 375) <= 0; flappy_W(14, 376) <= 0; flappy_W(14, 377) <= 0; flappy_W(14, 378) <= 0; flappy_W(14, 379) <= 0; flappy_W(14, 380) <= 0; flappy_W(14, 381) <= 0; flappy_W(14, 382) <= 0; flappy_W(14, 383) <= 0; flappy_W(14, 384) <= 0; flappy_W(14, 385) <= 0; flappy_W(14, 386) <= 0; flappy_W(14, 387) <= 0; flappy_W(14, 388) <= 0; flappy_W(14, 389) <= 0; flappy_W(14, 390) <= 0; flappy_W(14, 391) <= 0; flappy_W(14, 392) <= 0; flappy_W(14, 393) <= 0; flappy_W(14, 394) <= 0; flappy_W(14, 395) <= 0; flappy_W(14, 396) <= 0; flappy_W(14, 397) <= 0; flappy_W(14, 398) <= 0; flappy_W(14, 399) <= 0; flappy_W(14, 400) <= 0; flappy_W(14, 401) <= 0; flappy_W(14, 402) <= 1; flappy_W(14, 403) <= 1; flappy_W(14, 404) <= 1; flappy_W(14, 405) <= 1; flappy_W(14, 406) <= 1; flappy_W(14, 407) <= 1; flappy_W(14, 408) <= 1; flappy_W(14, 409) <= 1; flappy_W(14, 410) <= 1; flappy_W(14, 411) <= 1; flappy_W(14, 412) <= 1; flappy_W(14, 413) <= 1; flappy_W(14, 414) <= 0; flappy_W(14, 415) <= 0; flappy_W(14, 416) <= 0; flappy_W(14, 417) <= 0; flappy_W(14, 418) <= 0; flappy_W(14, 419) <= 0; flappy_W(14, 420) <= 0; flappy_W(14, 421) <= 0; flappy_W(14, 422) <= 0; flappy_W(14, 423) <= 0; flappy_W(14, 424) <= 0; flappy_W(14, 425) <= 0; flappy_W(14, 426) <= 1; flappy_W(14, 427) <= 1; flappy_W(14, 428) <= 1; flappy_W(14, 429) <= 1; flappy_W(14, 430) <= 1; flappy_W(14, 431) <= 1; flappy_W(14, 432) <= 1; flappy_W(14, 433) <= 1; flappy_W(14, 434) <= 1; flappy_W(14, 435) <= 1; flappy_W(14, 436) <= 1; flappy_W(14, 437) <= 1; flappy_W(14, 438) <= 0; flappy_W(14, 439) <= 0; flappy_W(14, 440) <= 0; flappy_W(14, 441) <= 0; flappy_W(14, 442) <= 0; flappy_W(14, 443) <= 0; flappy_W(14, 444) <= 0; flappy_W(14, 445) <= 0; flappy_W(14, 446) <= 0; flappy_W(14, 447) <= 0; flappy_W(14, 448) <= 0; flappy_W(14, 449) <= 0; flappy_W(14, 450) <= 0; flappy_W(14, 451) <= 0; flappy_W(14, 452) <= 0; flappy_W(14, 453) <= 0; flappy_W(14, 454) <= 0; flappy_W(14, 455) <= 0; flappy_W(14, 456) <= 0; flappy_W(14, 457) <= 0; flappy_W(14, 458) <= 0; flappy_W(14, 459) <= 0; flappy_W(14, 460) <= 0; flappy_W(14, 461) <= 0; flappy_W(14, 462) <= 0; flappy_W(14, 463) <= 0; flappy_W(14, 464) <= 0; flappy_W(14, 465) <= 0; flappy_W(14, 466) <= 0; flappy_W(14, 467) <= 0; flappy_W(14, 468) <= 1; flappy_W(14, 469) <= 1; flappy_W(14, 470) <= 1; flappy_W(14, 471) <= 1; flappy_W(14, 472) <= 1; flappy_W(14, 473) <= 1; flappy_W(14, 474) <= 1; flappy_W(14, 475) <= 1; flappy_W(14, 476) <= 1; flappy_W(14, 477) <= 1; flappy_W(14, 478) <= 1; flappy_W(14, 479) <= 1; flappy_W(14, 480) <= 0; flappy_W(14, 481) <= 0; flappy_W(14, 482) <= 0; flappy_W(14, 483) <= 0; flappy_W(14, 484) <= 0; flappy_W(14, 485) <= 0; flappy_W(14, 486) <= 0; flappy_W(14, 487) <= 0; flappy_W(14, 488) <= 0; flappy_W(14, 489) <= 0; flappy_W(14, 490) <= 0; flappy_W(14, 491) <= 0; flappy_W(14, 492) <= 0; flappy_W(14, 493) <= 0; flappy_W(14, 494) <= 0; flappy_W(14, 495) <= 0; flappy_W(14, 496) <= 0; flappy_W(14, 497) <= 0; flappy_W(14, 498) <= 0; flappy_W(14, 499) <= 0; flappy_W(14, 500) <= 0; flappy_W(14, 501) <= 0; flappy_W(14, 502) <= 0; flappy_W(14, 503) <= 0; flappy_W(14, 504) <= 0; flappy_W(14, 505) <= 0; flappy_W(14, 506) <= 0; flappy_W(14, 507) <= 0; flappy_W(14, 508) <= 0; flappy_W(14, 509) <= 0; flappy_W(14, 510) <= 1; flappy_W(14, 511) <= 1; flappy_W(14, 512) <= 1; flappy_W(14, 513) <= 1; flappy_W(14, 514) <= 1; flappy_W(14, 515) <= 1; flappy_W(14, 516) <= 1; flappy_W(14, 517) <= 1; flappy_W(14, 518) <= 1; flappy_W(14, 519) <= 1; flappy_W(14, 520) <= 1; flappy_W(14, 521) <= 1; flappy_W(14, 522) <= 0; flappy_W(14, 523) <= 0; flappy_W(14, 524) <= 0; flappy_W(14, 525) <= 0; flappy_W(14, 526) <= 0; flappy_W(14, 527) <= 0; flappy_W(14, 528) <= 0; flappy_W(14, 529) <= 0; flappy_W(14, 530) <= 0; flappy_W(14, 531) <= 0; flappy_W(14, 532) <= 0; flappy_W(14, 533) <= 0; flappy_W(14, 534) <= 1; flappy_W(14, 535) <= 1; flappy_W(14, 536) <= 1; flappy_W(14, 537) <= 1; flappy_W(14, 538) <= 1; flappy_W(14, 539) <= 1; flappy_W(14, 540) <= 1; flappy_W(14, 541) <= 1; flappy_W(14, 542) <= 1; flappy_W(14, 543) <= 1; flappy_W(14, 544) <= 1; flappy_W(14, 545) <= 1; flappy_W(14, 546) <= 0; flappy_W(14, 547) <= 0; flappy_W(14, 548) <= 0; flappy_W(14, 549) <= 0; flappy_W(14, 550) <= 0; flappy_W(14, 551) <= 0; flappy_W(14, 552) <= 0; flappy_W(14, 553) <= 0; flappy_W(14, 554) <= 0; flappy_W(14, 555) <= 0; flappy_W(14, 556) <= 0; flappy_W(14, 557) <= 0; flappy_W(14, 558) <= 0; flappy_W(14, 559) <= 0; flappy_W(14, 560) <= 0; flappy_W(14, 561) <= 0; flappy_W(14, 562) <= 0; flappy_W(14, 563) <= 0; flappy_W(14, 564) <= 1; flappy_W(14, 565) <= 1; flappy_W(14, 566) <= 1; flappy_W(14, 567) <= 1; flappy_W(14, 568) <= 1; flappy_W(14, 569) <= 1; flappy_W(14, 570) <= 1; flappy_W(14, 571) <= 1; flappy_W(14, 572) <= 1; flappy_W(14, 573) <= 1; flappy_W(14, 574) <= 1; flappy_W(14, 575) <= 1; flappy_W(14, 576) <= 0; flappy_W(14, 577) <= 0; flappy_W(14, 578) <= 0; flappy_W(14, 579) <= 0; flappy_W(14, 580) <= 0; flappy_W(14, 581) <= 0; flappy_W(14, 582) <= 0; flappy_W(14, 583) <= 0; flappy_W(14, 584) <= 0; flappy_W(14, 585) <= 0; flappy_W(14, 586) <= 0; flappy_W(14, 587) <= 0; flappy_W(14, 588) <= 1; flappy_W(14, 589) <= 1; flappy_W(14, 590) <= 1; flappy_W(14, 591) <= 1; flappy_W(14, 592) <= 1; flappy_W(14, 593) <= 1; 
flappy_W(15, 0) <= 0; flappy_W(15, 1) <= 0; flappy_W(15, 2) <= 0; flappy_W(15, 3) <= 0; flappy_W(15, 4) <= 0; flappy_W(15, 5) <= 0; flappy_W(15, 6) <= 1; flappy_W(15, 7) <= 1; flappy_W(15, 8) <= 1; flappy_W(15, 9) <= 1; flappy_W(15, 10) <= 1; flappy_W(15, 11) <= 1; flappy_W(15, 12) <= 1; flappy_W(15, 13) <= 1; flappy_W(15, 14) <= 1; flappy_W(15, 15) <= 1; flappy_W(15, 16) <= 1; flappy_W(15, 17) <= 1; flappy_W(15, 18) <= 0; flappy_W(15, 19) <= 0; flappy_W(15, 20) <= 0; flappy_W(15, 21) <= 0; flappy_W(15, 22) <= 0; flappy_W(15, 23) <= 0; flappy_W(15, 24) <= 0; flappy_W(15, 25) <= 0; flappy_W(15, 26) <= 0; flappy_W(15, 27) <= 0; flappy_W(15, 28) <= 0; flappy_W(15, 29) <= 0; flappy_W(15, 30) <= 0; flappy_W(15, 31) <= 0; flappy_W(15, 32) <= 0; flappy_W(15, 33) <= 0; flappy_W(15, 34) <= 0; flappy_W(15, 35) <= 0; flappy_W(15, 36) <= 1; flappy_W(15, 37) <= 1; flappy_W(15, 38) <= 1; flappy_W(15, 39) <= 1; flappy_W(15, 40) <= 1; flappy_W(15, 41) <= 1; flappy_W(15, 42) <= 0; flappy_W(15, 43) <= 0; flappy_W(15, 44) <= 0; flappy_W(15, 45) <= 0; flappy_W(15, 46) <= 0; flappy_W(15, 47) <= 0; flappy_W(15, 48) <= 0; flappy_W(15, 49) <= 0; flappy_W(15, 50) <= 0; flappy_W(15, 51) <= 0; flappy_W(15, 52) <= 0; flappy_W(15, 53) <= 0; flappy_W(15, 54) <= 0; flappy_W(15, 55) <= 0; flappy_W(15, 56) <= 0; flappy_W(15, 57) <= 0; flappy_W(15, 58) <= 0; flappy_W(15, 59) <= 0; flappy_W(15, 60) <= 1; flappy_W(15, 61) <= 1; flappy_W(15, 62) <= 1; flappy_W(15, 63) <= 1; flappy_W(15, 64) <= 1; flappy_W(15, 65) <= 1; flappy_W(15, 66) <= 1; flappy_W(15, 67) <= 1; flappy_W(15, 68) <= 1; flappy_W(15, 69) <= 1; flappy_W(15, 70) <= 1; flappy_W(15, 71) <= 1; flappy_W(15, 72) <= 0; flappy_W(15, 73) <= 0; flappy_W(15, 74) <= 0; flappy_W(15, 75) <= 0; flappy_W(15, 76) <= 0; flappy_W(15, 77) <= 0; flappy_W(15, 78) <= 0; flappy_W(15, 79) <= 0; flappy_W(15, 80) <= 0; flappy_W(15, 81) <= 0; flappy_W(15, 82) <= 0; flappy_W(15, 83) <= 0; flappy_W(15, 84) <= 0; flappy_W(15, 85) <= 0; flappy_W(15, 86) <= 0; flappy_W(15, 87) <= 0; flappy_W(15, 88) <= 0; flappy_W(15, 89) <= 0; flappy_W(15, 90) <= 0; flappy_W(15, 91) <= 0; flappy_W(15, 92) <= 0; flappy_W(15, 93) <= 0; flappy_W(15, 94) <= 0; flappy_W(15, 95) <= 0; flappy_W(15, 96) <= 0; flappy_W(15, 97) <= 0; flappy_W(15, 98) <= 0; flappy_W(15, 99) <= 0; flappy_W(15, 100) <= 0; flappy_W(15, 101) <= 0; flappy_W(15, 102) <= 0; flappy_W(15, 103) <= 0; flappy_W(15, 104) <= 0; flappy_W(15, 105) <= 0; flappy_W(15, 106) <= 0; flappy_W(15, 107) <= 0; flappy_W(15, 108) <= 0; flappy_W(15, 109) <= 0; flappy_W(15, 110) <= 0; flappy_W(15, 111) <= 0; flappy_W(15, 112) <= 0; flappy_W(15, 113) <= 0; flappy_W(15, 114) <= 1; flappy_W(15, 115) <= 1; flappy_W(15, 116) <= 1; flappy_W(15, 117) <= 1; flappy_W(15, 118) <= 1; flappy_W(15, 119) <= 1; flappy_W(15, 120) <= 1; flappy_W(15, 121) <= 1; flappy_W(15, 122) <= 1; flappy_W(15, 123) <= 1; flappy_W(15, 124) <= 1; flappy_W(15, 125) <= 1; flappy_W(15, 126) <= 0; flappy_W(15, 127) <= 0; flappy_W(15, 128) <= 0; flappy_W(15, 129) <= 0; flappy_W(15, 130) <= 0; flappy_W(15, 131) <= 0; flappy_W(15, 132) <= 1; flappy_W(15, 133) <= 1; flappy_W(15, 134) <= 1; flappy_W(15, 135) <= 1; flappy_W(15, 136) <= 1; flappy_W(15, 137) <= 1; flappy_W(15, 138) <= 1; flappy_W(15, 139) <= 1; flappy_W(15, 140) <= 1; flappy_W(15, 141) <= 1; flappy_W(15, 142) <= 1; flappy_W(15, 143) <= 1; flappy_W(15, 144) <= 0; flappy_W(15, 145) <= 0; flappy_W(15, 146) <= 0; flappy_W(15, 147) <= 0; flappy_W(15, 148) <= 0; flappy_W(15, 149) <= 0; flappy_W(15, 150) <= 0; flappy_W(15, 151) <= 0; flappy_W(15, 152) <= 0; flappy_W(15, 153) <= 0; flappy_W(15, 154) <= 0; flappy_W(15, 155) <= 0; flappy_W(15, 156) <= 0; flappy_W(15, 157) <= 0; flappy_W(15, 158) <= 0; flappy_W(15, 159) <= 0; flappy_W(15, 160) <= 0; flappy_W(15, 161) <= 0; flappy_W(15, 162) <= 0; flappy_W(15, 163) <= 0; flappy_W(15, 164) <= 0; flappy_W(15, 165) <= 0; flappy_W(15, 166) <= 0; flappy_W(15, 167) <= 0; flappy_W(15, 168) <= 1; flappy_W(15, 169) <= 1; flappy_W(15, 170) <= 1; flappy_W(15, 171) <= 1; flappy_W(15, 172) <= 1; flappy_W(15, 173) <= 1; flappy_W(15, 174) <= 1; flappy_W(15, 175) <= 1; flappy_W(15, 176) <= 1; flappy_W(15, 177) <= 1; flappy_W(15, 178) <= 1; flappy_W(15, 179) <= 1; flappy_W(15, 180) <= 0; flappy_W(15, 181) <= 0; flappy_W(15, 182) <= 0; flappy_W(15, 183) <= 0; flappy_W(15, 184) <= 0; flappy_W(15, 185) <= 0; flappy_W(15, 186) <= 0; flappy_W(15, 187) <= 0; flappy_W(15, 188) <= 0; flappy_W(15, 189) <= 0; flappy_W(15, 190) <= 0; flappy_W(15, 191) <= 0; flappy_W(15, 192) <= 1; flappy_W(15, 193) <= 1; flappy_W(15, 194) <= 1; flappy_W(15, 195) <= 1; flappy_W(15, 196) <= 1; flappy_W(15, 197) <= 1; flappy_W(15, 198) <= 1; flappy_W(15, 199) <= 1; flappy_W(15, 200) <= 1; flappy_W(15, 201) <= 1; flappy_W(15, 202) <= 1; flappy_W(15, 203) <= 1; flappy_W(15, 204) <= 0; flappy_W(15, 205) <= 0; flappy_W(15, 206) <= 0; flappy_W(15, 207) <= 0; flappy_W(15, 208) <= 0; flappy_W(15, 209) <= 0; flappy_W(15, 210) <= 0; flappy_W(15, 211) <= 0; flappy_W(15, 212) <= 0; flappy_W(15, 213) <= 0; flappy_W(15, 214) <= 0; flappy_W(15, 215) <= 0; flappy_W(15, 216) <= 0; flappy_W(15, 217) <= 0; flappy_W(15, 218) <= 0; flappy_W(15, 219) <= 0; flappy_W(15, 220) <= 0; flappy_W(15, 221) <= 0; flappy_W(15, 222) <= 1; flappy_W(15, 223) <= 1; flappy_W(15, 224) <= 1; flappy_W(15, 225) <= 1; flappy_W(15, 226) <= 1; flappy_W(15, 227) <= 1; flappy_W(15, 228) <= 1; flappy_W(15, 229) <= 1; flappy_W(15, 230) <= 1; flappy_W(15, 231) <= 1; flappy_W(15, 232) <= 1; flappy_W(15, 233) <= 1; flappy_W(15, 234) <= 0; flappy_W(15, 235) <= 0; flappy_W(15, 236) <= 0; flappy_W(15, 237) <= 0; flappy_W(15, 238) <= 0; flappy_W(15, 239) <= 0; flappy_W(15, 240) <= 0; flappy_W(15, 241) <= 0; flappy_W(15, 242) <= 0; flappy_W(15, 243) <= 0; flappy_W(15, 244) <= 0; flappy_W(15, 245) <= 0; flappy_W(15, 246) <= 1; flappy_W(15, 247) <= 1; flappy_W(15, 248) <= 1; flappy_W(15, 249) <= 1; flappy_W(15, 250) <= 1; flappy_W(15, 251) <= 1; flappy_W(15, 252) <= 1; flappy_W(15, 253) <= 1; flappy_W(15, 254) <= 1; flappy_W(15, 255) <= 1; flappy_W(15, 256) <= 1; flappy_W(15, 257) <= 1; flappy_W(15, 258) <= 0; flappy_W(15, 259) <= 0; flappy_W(15, 260) <= 0; flappy_W(15, 261) <= 0; flappy_W(15, 262) <= 0; flappy_W(15, 263) <= 0; flappy_W(15, 264) <= 0; flappy_W(15, 265) <= 0; flappy_W(15, 266) <= 0; flappy_W(15, 267) <= 0; flappy_W(15, 268) <= 0; flappy_W(15, 269) <= 0; flappy_W(15, 270) <= 1; flappy_W(15, 271) <= 1; flappy_W(15, 272) <= 1; flappy_W(15, 273) <= 1; flappy_W(15, 274) <= 1; flappy_W(15, 275) <= 1; flappy_W(15, 276) <= 1; flappy_W(15, 277) <= 1; flappy_W(15, 278) <= 1; flappy_W(15, 279) <= 1; flappy_W(15, 280) <= 1; flappy_W(15, 281) <= 1; flappy_W(15, 282) <= 0; flappy_W(15, 283) <= 0; flappy_W(15, 284) <= 0; flappy_W(15, 285) <= 0; flappy_W(15, 286) <= 0; flappy_W(15, 287) <= 0; flappy_W(15, 288) <= 0; flappy_W(15, 289) <= 0; flappy_W(15, 290) <= 0; flappy_W(15, 291) <= 0; flappy_W(15, 292) <= 0; flappy_W(15, 293) <= 0; flappy_W(15, 294) <= 0; flappy_W(15, 295) <= 0; flappy_W(15, 296) <= 0; flappy_W(15, 297) <= 0; flappy_W(15, 298) <= 0; flappy_W(15, 299) <= 0; flappy_W(15, 300) <= 0; flappy_W(15, 301) <= 0; flappy_W(15, 302) <= 0; flappy_W(15, 303) <= 0; flappy_W(15, 304) <= 0; flappy_W(15, 305) <= 0; flappy_W(15, 306) <= 1; flappy_W(15, 307) <= 1; flappy_W(15, 308) <= 1; flappy_W(15, 309) <= 1; flappy_W(15, 310) <= 1; flappy_W(15, 311) <= 1; flappy_W(15, 312) <= 1; flappy_W(15, 313) <= 1; flappy_W(15, 314) <= 1; flappy_W(15, 315) <= 1; flappy_W(15, 316) <= 1; flappy_W(15, 317) <= 1; flappy_W(15, 318) <= 0; flappy_W(15, 319) <= 0; flappy_W(15, 320) <= 0; flappy_W(15, 321) <= 0; flappy_W(15, 322) <= 0; flappy_W(15, 323) <= 0; flappy_W(15, 324) <= 0; flappy_W(15, 325) <= 0; flappy_W(15, 326) <= 0; flappy_W(15, 327) <= 0; flappy_W(15, 328) <= 0; flappy_W(15, 329) <= 0; flappy_W(15, 330) <= 0; flappy_W(15, 331) <= 0; flappy_W(15, 332) <= 0; flappy_W(15, 333) <= 0; flappy_W(15, 334) <= 0; flappy_W(15, 335) <= 0; flappy_W(15, 336) <= 0; flappy_W(15, 337) <= 0; flappy_W(15, 338) <= 0; flappy_W(15, 339) <= 0; flappy_W(15, 340) <= 0; flappy_W(15, 341) <= 0; flappy_W(15, 342) <= 0; flappy_W(15, 343) <= 0; flappy_W(15, 344) <= 0; flappy_W(15, 345) <= 0; flappy_W(15, 346) <= 0; flappy_W(15, 347) <= 0; flappy_W(15, 348) <= 0; flappy_W(15, 349) <= 0; flappy_W(15, 350) <= 0; flappy_W(15, 351) <= 0; flappy_W(15, 352) <= 0; flappy_W(15, 353) <= 0; flappy_W(15, 354) <= 0; flappy_W(15, 355) <= 0; flappy_W(15, 356) <= 0; flappy_W(15, 357) <= 0; flappy_W(15, 358) <= 0; flappy_W(15, 359) <= 0; flappy_W(15, 360) <= 0; flappy_W(15, 361) <= 0; flappy_W(15, 362) <= 0; flappy_W(15, 363) <= 0; flappy_W(15, 364) <= 0; flappy_W(15, 365) <= 0; flappy_W(15, 366) <= 0; flappy_W(15, 367) <= 0; flappy_W(15, 368) <= 0; flappy_W(15, 369) <= 0; flappy_W(15, 370) <= 0; flappy_W(15, 371) <= 0; flappy_W(15, 372) <= 0; flappy_W(15, 373) <= 0; flappy_W(15, 374) <= 0; flappy_W(15, 375) <= 0; flappy_W(15, 376) <= 0; flappy_W(15, 377) <= 0; flappy_W(15, 378) <= 0; flappy_W(15, 379) <= 0; flappy_W(15, 380) <= 0; flappy_W(15, 381) <= 0; flappy_W(15, 382) <= 0; flappy_W(15, 383) <= 0; flappy_W(15, 384) <= 0; flappy_W(15, 385) <= 0; flappy_W(15, 386) <= 0; flappy_W(15, 387) <= 0; flappy_W(15, 388) <= 0; flappy_W(15, 389) <= 0; flappy_W(15, 390) <= 0; flappy_W(15, 391) <= 0; flappy_W(15, 392) <= 0; flappy_W(15, 393) <= 0; flappy_W(15, 394) <= 0; flappy_W(15, 395) <= 0; flappy_W(15, 396) <= 0; flappy_W(15, 397) <= 0; flappy_W(15, 398) <= 0; flappy_W(15, 399) <= 0; flappy_W(15, 400) <= 0; flappy_W(15, 401) <= 0; flappy_W(15, 402) <= 1; flappy_W(15, 403) <= 1; flappy_W(15, 404) <= 1; flappy_W(15, 405) <= 1; flappy_W(15, 406) <= 1; flappy_W(15, 407) <= 1; flappy_W(15, 408) <= 1; flappy_W(15, 409) <= 1; flappy_W(15, 410) <= 1; flappy_W(15, 411) <= 1; flappy_W(15, 412) <= 1; flappy_W(15, 413) <= 1; flappy_W(15, 414) <= 0; flappy_W(15, 415) <= 0; flappy_W(15, 416) <= 0; flappy_W(15, 417) <= 0; flappy_W(15, 418) <= 0; flappy_W(15, 419) <= 0; flappy_W(15, 420) <= 0; flappy_W(15, 421) <= 0; flappy_W(15, 422) <= 0; flappy_W(15, 423) <= 0; flappy_W(15, 424) <= 0; flappy_W(15, 425) <= 0; flappy_W(15, 426) <= 1; flappy_W(15, 427) <= 1; flappy_W(15, 428) <= 1; flappy_W(15, 429) <= 1; flappy_W(15, 430) <= 1; flappy_W(15, 431) <= 1; flappy_W(15, 432) <= 1; flappy_W(15, 433) <= 1; flappy_W(15, 434) <= 1; flappy_W(15, 435) <= 1; flappy_W(15, 436) <= 1; flappy_W(15, 437) <= 1; flappy_W(15, 438) <= 0; flappy_W(15, 439) <= 0; flappy_W(15, 440) <= 0; flappy_W(15, 441) <= 0; flappy_W(15, 442) <= 0; flappy_W(15, 443) <= 0; flappy_W(15, 444) <= 0; flappy_W(15, 445) <= 0; flappy_W(15, 446) <= 0; flappy_W(15, 447) <= 0; flappy_W(15, 448) <= 0; flappy_W(15, 449) <= 0; flappy_W(15, 450) <= 0; flappy_W(15, 451) <= 0; flappy_W(15, 452) <= 0; flappy_W(15, 453) <= 0; flappy_W(15, 454) <= 0; flappy_W(15, 455) <= 0; flappy_W(15, 456) <= 0; flappy_W(15, 457) <= 0; flappy_W(15, 458) <= 0; flappy_W(15, 459) <= 0; flappy_W(15, 460) <= 0; flappy_W(15, 461) <= 0; flappy_W(15, 462) <= 0; flappy_W(15, 463) <= 0; flappy_W(15, 464) <= 0; flappy_W(15, 465) <= 0; flappy_W(15, 466) <= 0; flappy_W(15, 467) <= 0; flappy_W(15, 468) <= 1; flappy_W(15, 469) <= 1; flappy_W(15, 470) <= 1; flappy_W(15, 471) <= 1; flappy_W(15, 472) <= 1; flappy_W(15, 473) <= 1; flappy_W(15, 474) <= 1; flappy_W(15, 475) <= 1; flappy_W(15, 476) <= 1; flappy_W(15, 477) <= 1; flappy_W(15, 478) <= 1; flappy_W(15, 479) <= 1; flappy_W(15, 480) <= 0; flappy_W(15, 481) <= 0; flappy_W(15, 482) <= 0; flappy_W(15, 483) <= 0; flappy_W(15, 484) <= 0; flappy_W(15, 485) <= 0; flappy_W(15, 486) <= 0; flappy_W(15, 487) <= 0; flappy_W(15, 488) <= 0; flappy_W(15, 489) <= 0; flappy_W(15, 490) <= 0; flappy_W(15, 491) <= 0; flappy_W(15, 492) <= 0; flappy_W(15, 493) <= 0; flappy_W(15, 494) <= 0; flappy_W(15, 495) <= 0; flappy_W(15, 496) <= 0; flappy_W(15, 497) <= 0; flappy_W(15, 498) <= 0; flappy_W(15, 499) <= 0; flappy_W(15, 500) <= 0; flappy_W(15, 501) <= 0; flappy_W(15, 502) <= 0; flappy_W(15, 503) <= 0; flappy_W(15, 504) <= 0; flappy_W(15, 505) <= 0; flappy_W(15, 506) <= 0; flappy_W(15, 507) <= 0; flappy_W(15, 508) <= 0; flappy_W(15, 509) <= 0; flappy_W(15, 510) <= 1; flappy_W(15, 511) <= 1; flappy_W(15, 512) <= 1; flappy_W(15, 513) <= 1; flappy_W(15, 514) <= 1; flappy_W(15, 515) <= 1; flappy_W(15, 516) <= 1; flappy_W(15, 517) <= 1; flappy_W(15, 518) <= 1; flappy_W(15, 519) <= 1; flappy_W(15, 520) <= 1; flappy_W(15, 521) <= 1; flappy_W(15, 522) <= 0; flappy_W(15, 523) <= 0; flappy_W(15, 524) <= 0; flappy_W(15, 525) <= 0; flappy_W(15, 526) <= 0; flappy_W(15, 527) <= 0; flappy_W(15, 528) <= 0; flappy_W(15, 529) <= 0; flappy_W(15, 530) <= 0; flappy_W(15, 531) <= 0; flappy_W(15, 532) <= 0; flappy_W(15, 533) <= 0; flappy_W(15, 534) <= 1; flappy_W(15, 535) <= 1; flappy_W(15, 536) <= 1; flappy_W(15, 537) <= 1; flappy_W(15, 538) <= 1; flappy_W(15, 539) <= 1; flappy_W(15, 540) <= 1; flappy_W(15, 541) <= 1; flappy_W(15, 542) <= 1; flappy_W(15, 543) <= 1; flappy_W(15, 544) <= 1; flappy_W(15, 545) <= 1; flappy_W(15, 546) <= 0; flappy_W(15, 547) <= 0; flappy_W(15, 548) <= 0; flappy_W(15, 549) <= 0; flappy_W(15, 550) <= 0; flappy_W(15, 551) <= 0; flappy_W(15, 552) <= 0; flappy_W(15, 553) <= 0; flappy_W(15, 554) <= 0; flappy_W(15, 555) <= 0; flappy_W(15, 556) <= 0; flappy_W(15, 557) <= 0; flappy_W(15, 558) <= 0; flappy_W(15, 559) <= 0; flappy_W(15, 560) <= 0; flappy_W(15, 561) <= 0; flappy_W(15, 562) <= 0; flappy_W(15, 563) <= 0; flappy_W(15, 564) <= 1; flappy_W(15, 565) <= 1; flappy_W(15, 566) <= 1; flappy_W(15, 567) <= 1; flappy_W(15, 568) <= 1; flappy_W(15, 569) <= 1; flappy_W(15, 570) <= 1; flappy_W(15, 571) <= 1; flappy_W(15, 572) <= 1; flappy_W(15, 573) <= 1; flappy_W(15, 574) <= 1; flappy_W(15, 575) <= 1; flappy_W(15, 576) <= 0; flappy_W(15, 577) <= 0; flappy_W(15, 578) <= 0; flappy_W(15, 579) <= 0; flappy_W(15, 580) <= 0; flappy_W(15, 581) <= 0; flappy_W(15, 582) <= 0; flappy_W(15, 583) <= 0; flappy_W(15, 584) <= 0; flappy_W(15, 585) <= 0; flappy_W(15, 586) <= 0; flappy_W(15, 587) <= 0; flappy_W(15, 588) <= 1; flappy_W(15, 589) <= 1; flappy_W(15, 590) <= 1; flappy_W(15, 591) <= 1; flappy_W(15, 592) <= 1; flappy_W(15, 593) <= 1; 
flappy_W(16, 0) <= 0; flappy_W(16, 1) <= 0; flappy_W(16, 2) <= 0; flappy_W(16, 3) <= 0; flappy_W(16, 4) <= 0; flappy_W(16, 5) <= 0; flappy_W(16, 6) <= 1; flappy_W(16, 7) <= 1; flappy_W(16, 8) <= 1; flappy_W(16, 9) <= 1; flappy_W(16, 10) <= 1; flappy_W(16, 11) <= 1; flappy_W(16, 12) <= 1; flappy_W(16, 13) <= 1; flappy_W(16, 14) <= 1; flappy_W(16, 15) <= 1; flappy_W(16, 16) <= 1; flappy_W(16, 17) <= 1; flappy_W(16, 18) <= 0; flappy_W(16, 19) <= 0; flappy_W(16, 20) <= 0; flappy_W(16, 21) <= 0; flappy_W(16, 22) <= 0; flappy_W(16, 23) <= 0; flappy_W(16, 24) <= 0; flappy_W(16, 25) <= 0; flappy_W(16, 26) <= 0; flappy_W(16, 27) <= 0; flappy_W(16, 28) <= 0; flappy_W(16, 29) <= 0; flappy_W(16, 30) <= 0; flappy_W(16, 31) <= 0; flappy_W(16, 32) <= 0; flappy_W(16, 33) <= 0; flappy_W(16, 34) <= 0; flappy_W(16, 35) <= 0; flappy_W(16, 36) <= 1; flappy_W(16, 37) <= 1; flappy_W(16, 38) <= 1; flappy_W(16, 39) <= 1; flappy_W(16, 40) <= 1; flappy_W(16, 41) <= 1; flappy_W(16, 42) <= 0; flappy_W(16, 43) <= 0; flappy_W(16, 44) <= 0; flappy_W(16, 45) <= 0; flappy_W(16, 46) <= 0; flappy_W(16, 47) <= 0; flappy_W(16, 48) <= 0; flappy_W(16, 49) <= 0; flappy_W(16, 50) <= 0; flappy_W(16, 51) <= 0; flappy_W(16, 52) <= 0; flappy_W(16, 53) <= 0; flappy_W(16, 54) <= 0; flappy_W(16, 55) <= 0; flappy_W(16, 56) <= 0; flappy_W(16, 57) <= 0; flappy_W(16, 58) <= 0; flappy_W(16, 59) <= 0; flappy_W(16, 60) <= 1; flappy_W(16, 61) <= 1; flappy_W(16, 62) <= 1; flappy_W(16, 63) <= 1; flappy_W(16, 64) <= 1; flappy_W(16, 65) <= 1; flappy_W(16, 66) <= 1; flappy_W(16, 67) <= 1; flappy_W(16, 68) <= 1; flappy_W(16, 69) <= 1; flappy_W(16, 70) <= 1; flappy_W(16, 71) <= 1; flappy_W(16, 72) <= 0; flappy_W(16, 73) <= 0; flappy_W(16, 74) <= 0; flappy_W(16, 75) <= 0; flappy_W(16, 76) <= 0; flappy_W(16, 77) <= 0; flappy_W(16, 78) <= 0; flappy_W(16, 79) <= 0; flappy_W(16, 80) <= 0; flappy_W(16, 81) <= 0; flappy_W(16, 82) <= 0; flappy_W(16, 83) <= 0; flappy_W(16, 84) <= 0; flappy_W(16, 85) <= 0; flappy_W(16, 86) <= 0; flappy_W(16, 87) <= 0; flappy_W(16, 88) <= 0; flappy_W(16, 89) <= 0; flappy_W(16, 90) <= 0; flappy_W(16, 91) <= 0; flappy_W(16, 92) <= 0; flappy_W(16, 93) <= 0; flappy_W(16, 94) <= 0; flappy_W(16, 95) <= 0; flappy_W(16, 96) <= 0; flappy_W(16, 97) <= 0; flappy_W(16, 98) <= 0; flappy_W(16, 99) <= 0; flappy_W(16, 100) <= 0; flappy_W(16, 101) <= 0; flappy_W(16, 102) <= 0; flappy_W(16, 103) <= 0; flappy_W(16, 104) <= 0; flappy_W(16, 105) <= 0; flappy_W(16, 106) <= 0; flappy_W(16, 107) <= 0; flappy_W(16, 108) <= 0; flappy_W(16, 109) <= 0; flappy_W(16, 110) <= 0; flappy_W(16, 111) <= 0; flappy_W(16, 112) <= 0; flappy_W(16, 113) <= 0; flappy_W(16, 114) <= 1; flappy_W(16, 115) <= 1; flappy_W(16, 116) <= 1; flappy_W(16, 117) <= 1; flappy_W(16, 118) <= 1; flappy_W(16, 119) <= 1; flappy_W(16, 120) <= 1; flappy_W(16, 121) <= 1; flappy_W(16, 122) <= 1; flappy_W(16, 123) <= 1; flappy_W(16, 124) <= 1; flappy_W(16, 125) <= 1; flappy_W(16, 126) <= 0; flappy_W(16, 127) <= 0; flappy_W(16, 128) <= 0; flappy_W(16, 129) <= 0; flappy_W(16, 130) <= 0; flappy_W(16, 131) <= 0; flappy_W(16, 132) <= 1; flappy_W(16, 133) <= 1; flappy_W(16, 134) <= 1; flappy_W(16, 135) <= 1; flappy_W(16, 136) <= 1; flappy_W(16, 137) <= 1; flappy_W(16, 138) <= 1; flappy_W(16, 139) <= 1; flappy_W(16, 140) <= 1; flappy_W(16, 141) <= 1; flappy_W(16, 142) <= 1; flappy_W(16, 143) <= 1; flappy_W(16, 144) <= 0; flappy_W(16, 145) <= 0; flappy_W(16, 146) <= 0; flappy_W(16, 147) <= 0; flappy_W(16, 148) <= 0; flappy_W(16, 149) <= 0; flappy_W(16, 150) <= 0; flappy_W(16, 151) <= 0; flappy_W(16, 152) <= 0; flappy_W(16, 153) <= 0; flappy_W(16, 154) <= 0; flappy_W(16, 155) <= 0; flappy_W(16, 156) <= 0; flappy_W(16, 157) <= 0; flappy_W(16, 158) <= 0; flappy_W(16, 159) <= 0; flappy_W(16, 160) <= 0; flappy_W(16, 161) <= 0; flappy_W(16, 162) <= 0; flappy_W(16, 163) <= 0; flappy_W(16, 164) <= 0; flappy_W(16, 165) <= 0; flappy_W(16, 166) <= 0; flappy_W(16, 167) <= 0; flappy_W(16, 168) <= 1; flappy_W(16, 169) <= 1; flappy_W(16, 170) <= 1; flappy_W(16, 171) <= 1; flappy_W(16, 172) <= 1; flappy_W(16, 173) <= 1; flappy_W(16, 174) <= 1; flappy_W(16, 175) <= 1; flappy_W(16, 176) <= 1; flappy_W(16, 177) <= 1; flappy_W(16, 178) <= 1; flappy_W(16, 179) <= 1; flappy_W(16, 180) <= 0; flappy_W(16, 181) <= 0; flappy_W(16, 182) <= 0; flappy_W(16, 183) <= 0; flappy_W(16, 184) <= 0; flappy_W(16, 185) <= 0; flappy_W(16, 186) <= 0; flappy_W(16, 187) <= 0; flappy_W(16, 188) <= 0; flappy_W(16, 189) <= 0; flappy_W(16, 190) <= 0; flappy_W(16, 191) <= 0; flappy_W(16, 192) <= 1; flappy_W(16, 193) <= 1; flappy_W(16, 194) <= 1; flappy_W(16, 195) <= 1; flappy_W(16, 196) <= 1; flappy_W(16, 197) <= 1; flappy_W(16, 198) <= 1; flappy_W(16, 199) <= 1; flappy_W(16, 200) <= 1; flappy_W(16, 201) <= 1; flappy_W(16, 202) <= 1; flappy_W(16, 203) <= 1; flappy_W(16, 204) <= 0; flappy_W(16, 205) <= 0; flappy_W(16, 206) <= 0; flappy_W(16, 207) <= 0; flappy_W(16, 208) <= 0; flappy_W(16, 209) <= 0; flappy_W(16, 210) <= 0; flappy_W(16, 211) <= 0; flappy_W(16, 212) <= 0; flappy_W(16, 213) <= 0; flappy_W(16, 214) <= 0; flappy_W(16, 215) <= 0; flappy_W(16, 216) <= 0; flappy_W(16, 217) <= 0; flappy_W(16, 218) <= 0; flappy_W(16, 219) <= 0; flappy_W(16, 220) <= 0; flappy_W(16, 221) <= 0; flappy_W(16, 222) <= 1; flappy_W(16, 223) <= 1; flappy_W(16, 224) <= 1; flappy_W(16, 225) <= 1; flappy_W(16, 226) <= 1; flappy_W(16, 227) <= 1; flappy_W(16, 228) <= 1; flappy_W(16, 229) <= 1; flappy_W(16, 230) <= 1; flappy_W(16, 231) <= 1; flappy_W(16, 232) <= 1; flappy_W(16, 233) <= 1; flappy_W(16, 234) <= 0; flappy_W(16, 235) <= 0; flappy_W(16, 236) <= 0; flappy_W(16, 237) <= 0; flappy_W(16, 238) <= 0; flappy_W(16, 239) <= 0; flappy_W(16, 240) <= 0; flappy_W(16, 241) <= 0; flappy_W(16, 242) <= 0; flappy_W(16, 243) <= 0; flappy_W(16, 244) <= 0; flappy_W(16, 245) <= 0; flappy_W(16, 246) <= 1; flappy_W(16, 247) <= 1; flappy_W(16, 248) <= 1; flappy_W(16, 249) <= 1; flappy_W(16, 250) <= 1; flappy_W(16, 251) <= 1; flappy_W(16, 252) <= 1; flappy_W(16, 253) <= 1; flappy_W(16, 254) <= 1; flappy_W(16, 255) <= 1; flappy_W(16, 256) <= 1; flappy_W(16, 257) <= 1; flappy_W(16, 258) <= 0; flappy_W(16, 259) <= 0; flappy_W(16, 260) <= 0; flappy_W(16, 261) <= 0; flappy_W(16, 262) <= 0; flappy_W(16, 263) <= 0; flappy_W(16, 264) <= 0; flappy_W(16, 265) <= 0; flappy_W(16, 266) <= 0; flappy_W(16, 267) <= 0; flappy_W(16, 268) <= 0; flappy_W(16, 269) <= 0; flappy_W(16, 270) <= 1; flappy_W(16, 271) <= 1; flappy_W(16, 272) <= 1; flappy_W(16, 273) <= 1; flappy_W(16, 274) <= 1; flappy_W(16, 275) <= 1; flappy_W(16, 276) <= 1; flappy_W(16, 277) <= 1; flappy_W(16, 278) <= 1; flappy_W(16, 279) <= 1; flappy_W(16, 280) <= 1; flappy_W(16, 281) <= 1; flappy_W(16, 282) <= 0; flappy_W(16, 283) <= 0; flappy_W(16, 284) <= 0; flappy_W(16, 285) <= 0; flappy_W(16, 286) <= 0; flappy_W(16, 287) <= 0; flappy_W(16, 288) <= 0; flappy_W(16, 289) <= 0; flappy_W(16, 290) <= 0; flappy_W(16, 291) <= 0; flappy_W(16, 292) <= 0; flappy_W(16, 293) <= 0; flappy_W(16, 294) <= 0; flappy_W(16, 295) <= 0; flappy_W(16, 296) <= 0; flappy_W(16, 297) <= 0; flappy_W(16, 298) <= 0; flappy_W(16, 299) <= 0; flappy_W(16, 300) <= 0; flappy_W(16, 301) <= 0; flappy_W(16, 302) <= 0; flappy_W(16, 303) <= 0; flappy_W(16, 304) <= 0; flappy_W(16, 305) <= 0; flappy_W(16, 306) <= 1; flappy_W(16, 307) <= 1; flappy_W(16, 308) <= 1; flappy_W(16, 309) <= 1; flappy_W(16, 310) <= 1; flappy_W(16, 311) <= 1; flappy_W(16, 312) <= 1; flappy_W(16, 313) <= 1; flappy_W(16, 314) <= 1; flappy_W(16, 315) <= 1; flappy_W(16, 316) <= 1; flappy_W(16, 317) <= 1; flappy_W(16, 318) <= 0; flappy_W(16, 319) <= 0; flappy_W(16, 320) <= 0; flappy_W(16, 321) <= 0; flappy_W(16, 322) <= 0; flappy_W(16, 323) <= 0; flappy_W(16, 324) <= 0; flappy_W(16, 325) <= 0; flappy_W(16, 326) <= 0; flappy_W(16, 327) <= 0; flappy_W(16, 328) <= 0; flappy_W(16, 329) <= 0; flappy_W(16, 330) <= 0; flappy_W(16, 331) <= 0; flappy_W(16, 332) <= 0; flappy_W(16, 333) <= 0; flappy_W(16, 334) <= 0; flappy_W(16, 335) <= 0; flappy_W(16, 336) <= 0; flappy_W(16, 337) <= 0; flappy_W(16, 338) <= 0; flappy_W(16, 339) <= 0; flappy_W(16, 340) <= 0; flappy_W(16, 341) <= 0; flappy_W(16, 342) <= 0; flappy_W(16, 343) <= 0; flappy_W(16, 344) <= 0; flappy_W(16, 345) <= 0; flappy_W(16, 346) <= 0; flappy_W(16, 347) <= 0; flappy_W(16, 348) <= 0; flappy_W(16, 349) <= 0; flappy_W(16, 350) <= 0; flappy_W(16, 351) <= 0; flappy_W(16, 352) <= 0; flappy_W(16, 353) <= 0; flappy_W(16, 354) <= 0; flappy_W(16, 355) <= 0; flappy_W(16, 356) <= 0; flappy_W(16, 357) <= 0; flappy_W(16, 358) <= 0; flappy_W(16, 359) <= 0; flappy_W(16, 360) <= 0; flappy_W(16, 361) <= 0; flappy_W(16, 362) <= 0; flappy_W(16, 363) <= 0; flappy_W(16, 364) <= 0; flappy_W(16, 365) <= 0; flappy_W(16, 366) <= 0; flappy_W(16, 367) <= 0; flappy_W(16, 368) <= 0; flappy_W(16, 369) <= 0; flappy_W(16, 370) <= 0; flappy_W(16, 371) <= 0; flappy_W(16, 372) <= 0; flappy_W(16, 373) <= 0; flappy_W(16, 374) <= 0; flappy_W(16, 375) <= 0; flappy_W(16, 376) <= 0; flappy_W(16, 377) <= 0; flappy_W(16, 378) <= 0; flappy_W(16, 379) <= 0; flappy_W(16, 380) <= 0; flappy_W(16, 381) <= 0; flappy_W(16, 382) <= 0; flappy_W(16, 383) <= 0; flappy_W(16, 384) <= 0; flappy_W(16, 385) <= 0; flappy_W(16, 386) <= 0; flappy_W(16, 387) <= 0; flappy_W(16, 388) <= 0; flappy_W(16, 389) <= 0; flappy_W(16, 390) <= 0; flappy_W(16, 391) <= 0; flappy_W(16, 392) <= 0; flappy_W(16, 393) <= 0; flappy_W(16, 394) <= 0; flappy_W(16, 395) <= 0; flappy_W(16, 396) <= 0; flappy_W(16, 397) <= 0; flappy_W(16, 398) <= 0; flappy_W(16, 399) <= 0; flappy_W(16, 400) <= 0; flappy_W(16, 401) <= 0; flappy_W(16, 402) <= 1; flappy_W(16, 403) <= 1; flappy_W(16, 404) <= 1; flappy_W(16, 405) <= 1; flappy_W(16, 406) <= 1; flappy_W(16, 407) <= 1; flappy_W(16, 408) <= 1; flappy_W(16, 409) <= 1; flappy_W(16, 410) <= 1; flappy_W(16, 411) <= 1; flappy_W(16, 412) <= 1; flappy_W(16, 413) <= 1; flappy_W(16, 414) <= 0; flappy_W(16, 415) <= 0; flappy_W(16, 416) <= 0; flappy_W(16, 417) <= 0; flappy_W(16, 418) <= 0; flappy_W(16, 419) <= 0; flappy_W(16, 420) <= 0; flappy_W(16, 421) <= 0; flappy_W(16, 422) <= 0; flappy_W(16, 423) <= 0; flappy_W(16, 424) <= 0; flappy_W(16, 425) <= 0; flappy_W(16, 426) <= 1; flappy_W(16, 427) <= 1; flappy_W(16, 428) <= 1; flappy_W(16, 429) <= 1; flappy_W(16, 430) <= 1; flappy_W(16, 431) <= 1; flappy_W(16, 432) <= 1; flappy_W(16, 433) <= 1; flappy_W(16, 434) <= 1; flappy_W(16, 435) <= 1; flappy_W(16, 436) <= 1; flappy_W(16, 437) <= 1; flappy_W(16, 438) <= 0; flappy_W(16, 439) <= 0; flappy_W(16, 440) <= 0; flappy_W(16, 441) <= 0; flappy_W(16, 442) <= 0; flappy_W(16, 443) <= 0; flappy_W(16, 444) <= 0; flappy_W(16, 445) <= 0; flappy_W(16, 446) <= 0; flappy_W(16, 447) <= 0; flappy_W(16, 448) <= 0; flappy_W(16, 449) <= 0; flappy_W(16, 450) <= 0; flappy_W(16, 451) <= 0; flappy_W(16, 452) <= 0; flappy_W(16, 453) <= 0; flappy_W(16, 454) <= 0; flappy_W(16, 455) <= 0; flappy_W(16, 456) <= 0; flappy_W(16, 457) <= 0; flappy_W(16, 458) <= 0; flappy_W(16, 459) <= 0; flappy_W(16, 460) <= 0; flappy_W(16, 461) <= 0; flappy_W(16, 462) <= 0; flappy_W(16, 463) <= 0; flappy_W(16, 464) <= 0; flappy_W(16, 465) <= 0; flappy_W(16, 466) <= 0; flappy_W(16, 467) <= 0; flappy_W(16, 468) <= 1; flappy_W(16, 469) <= 1; flappy_W(16, 470) <= 1; flappy_W(16, 471) <= 1; flappy_W(16, 472) <= 1; flappy_W(16, 473) <= 1; flappy_W(16, 474) <= 1; flappy_W(16, 475) <= 1; flappy_W(16, 476) <= 1; flappy_W(16, 477) <= 1; flappy_W(16, 478) <= 1; flappy_W(16, 479) <= 1; flappy_W(16, 480) <= 0; flappy_W(16, 481) <= 0; flappy_W(16, 482) <= 0; flappy_W(16, 483) <= 0; flappy_W(16, 484) <= 0; flappy_W(16, 485) <= 0; flappy_W(16, 486) <= 0; flappy_W(16, 487) <= 0; flappy_W(16, 488) <= 0; flappy_W(16, 489) <= 0; flappy_W(16, 490) <= 0; flappy_W(16, 491) <= 0; flappy_W(16, 492) <= 0; flappy_W(16, 493) <= 0; flappy_W(16, 494) <= 0; flappy_W(16, 495) <= 0; flappy_W(16, 496) <= 0; flappy_W(16, 497) <= 0; flappy_W(16, 498) <= 0; flappy_W(16, 499) <= 0; flappy_W(16, 500) <= 0; flappy_W(16, 501) <= 0; flappy_W(16, 502) <= 0; flappy_W(16, 503) <= 0; flappy_W(16, 504) <= 0; flappy_W(16, 505) <= 0; flappy_W(16, 506) <= 0; flappy_W(16, 507) <= 0; flappy_W(16, 508) <= 0; flappy_W(16, 509) <= 0; flappy_W(16, 510) <= 1; flappy_W(16, 511) <= 1; flappy_W(16, 512) <= 1; flappy_W(16, 513) <= 1; flappy_W(16, 514) <= 1; flappy_W(16, 515) <= 1; flappy_W(16, 516) <= 1; flappy_W(16, 517) <= 1; flappy_W(16, 518) <= 1; flappy_W(16, 519) <= 1; flappy_W(16, 520) <= 1; flappy_W(16, 521) <= 1; flappy_W(16, 522) <= 0; flappy_W(16, 523) <= 0; flappy_W(16, 524) <= 0; flappy_W(16, 525) <= 0; flappy_W(16, 526) <= 0; flappy_W(16, 527) <= 0; flappy_W(16, 528) <= 0; flappy_W(16, 529) <= 0; flappy_W(16, 530) <= 0; flappy_W(16, 531) <= 0; flappy_W(16, 532) <= 0; flappy_W(16, 533) <= 0; flappy_W(16, 534) <= 1; flappy_W(16, 535) <= 1; flappy_W(16, 536) <= 1; flappy_W(16, 537) <= 1; flappy_W(16, 538) <= 1; flappy_W(16, 539) <= 1; flappy_W(16, 540) <= 1; flappy_W(16, 541) <= 1; flappy_W(16, 542) <= 1; flappy_W(16, 543) <= 1; flappy_W(16, 544) <= 1; flappy_W(16, 545) <= 1; flappy_W(16, 546) <= 0; flappy_W(16, 547) <= 0; flappy_W(16, 548) <= 0; flappy_W(16, 549) <= 0; flappy_W(16, 550) <= 0; flappy_W(16, 551) <= 0; flappy_W(16, 552) <= 0; flappy_W(16, 553) <= 0; flappy_W(16, 554) <= 0; flappy_W(16, 555) <= 0; flappy_W(16, 556) <= 0; flappy_W(16, 557) <= 0; flappy_W(16, 558) <= 0; flappy_W(16, 559) <= 0; flappy_W(16, 560) <= 0; flappy_W(16, 561) <= 0; flappy_W(16, 562) <= 0; flappy_W(16, 563) <= 0; flappy_W(16, 564) <= 1; flappy_W(16, 565) <= 1; flappy_W(16, 566) <= 1; flappy_W(16, 567) <= 1; flappy_W(16, 568) <= 1; flappy_W(16, 569) <= 1; flappy_W(16, 570) <= 1; flappy_W(16, 571) <= 1; flappy_W(16, 572) <= 1; flappy_W(16, 573) <= 1; flappy_W(16, 574) <= 1; flappy_W(16, 575) <= 1; flappy_W(16, 576) <= 0; flappy_W(16, 577) <= 0; flappy_W(16, 578) <= 0; flappy_W(16, 579) <= 0; flappy_W(16, 580) <= 0; flappy_W(16, 581) <= 0; flappy_W(16, 582) <= 0; flappy_W(16, 583) <= 0; flappy_W(16, 584) <= 0; flappy_W(16, 585) <= 0; flappy_W(16, 586) <= 0; flappy_W(16, 587) <= 0; flappy_W(16, 588) <= 1; flappy_W(16, 589) <= 1; flappy_W(16, 590) <= 1; flappy_W(16, 591) <= 1; flappy_W(16, 592) <= 1; flappy_W(16, 593) <= 1; 
flappy_W(17, 0) <= 0; flappy_W(17, 1) <= 0; flappy_W(17, 2) <= 0; flappy_W(17, 3) <= 0; flappy_W(17, 4) <= 0; flappy_W(17, 5) <= 0; flappy_W(17, 6) <= 1; flappy_W(17, 7) <= 1; flappy_W(17, 8) <= 1; flappy_W(17, 9) <= 1; flappy_W(17, 10) <= 1; flappy_W(17, 11) <= 1; flappy_W(17, 12) <= 1; flappy_W(17, 13) <= 1; flappy_W(17, 14) <= 1; flappy_W(17, 15) <= 1; flappy_W(17, 16) <= 1; flappy_W(17, 17) <= 1; flappy_W(17, 18) <= 0; flappy_W(17, 19) <= 0; flappy_W(17, 20) <= 0; flappy_W(17, 21) <= 0; flappy_W(17, 22) <= 0; flappy_W(17, 23) <= 0; flappy_W(17, 24) <= 0; flappy_W(17, 25) <= 0; flappy_W(17, 26) <= 0; flappy_W(17, 27) <= 0; flappy_W(17, 28) <= 0; flappy_W(17, 29) <= 0; flappy_W(17, 30) <= 0; flappy_W(17, 31) <= 0; flappy_W(17, 32) <= 0; flappy_W(17, 33) <= 0; flappy_W(17, 34) <= 0; flappy_W(17, 35) <= 0; flappy_W(17, 36) <= 1; flappy_W(17, 37) <= 1; flappy_W(17, 38) <= 1; flappy_W(17, 39) <= 1; flappy_W(17, 40) <= 1; flappy_W(17, 41) <= 1; flappy_W(17, 42) <= 0; flappy_W(17, 43) <= 0; flappy_W(17, 44) <= 0; flappy_W(17, 45) <= 0; flappy_W(17, 46) <= 0; flappy_W(17, 47) <= 0; flappy_W(17, 48) <= 0; flappy_W(17, 49) <= 0; flappy_W(17, 50) <= 0; flappy_W(17, 51) <= 0; flappy_W(17, 52) <= 0; flappy_W(17, 53) <= 0; flappy_W(17, 54) <= 0; flappy_W(17, 55) <= 0; flappy_W(17, 56) <= 0; flappy_W(17, 57) <= 0; flappy_W(17, 58) <= 0; flappy_W(17, 59) <= 0; flappy_W(17, 60) <= 1; flappy_W(17, 61) <= 1; flappy_W(17, 62) <= 1; flappy_W(17, 63) <= 1; flappy_W(17, 64) <= 1; flappy_W(17, 65) <= 1; flappy_W(17, 66) <= 1; flappy_W(17, 67) <= 1; flappy_W(17, 68) <= 1; flappy_W(17, 69) <= 1; flappy_W(17, 70) <= 1; flappy_W(17, 71) <= 1; flappy_W(17, 72) <= 0; flappy_W(17, 73) <= 0; flappy_W(17, 74) <= 0; flappy_W(17, 75) <= 0; flappy_W(17, 76) <= 0; flappy_W(17, 77) <= 0; flappy_W(17, 78) <= 0; flappy_W(17, 79) <= 0; flappy_W(17, 80) <= 0; flappy_W(17, 81) <= 0; flappy_W(17, 82) <= 0; flappy_W(17, 83) <= 0; flappy_W(17, 84) <= 0; flappy_W(17, 85) <= 0; flappy_W(17, 86) <= 0; flappy_W(17, 87) <= 0; flappy_W(17, 88) <= 0; flappy_W(17, 89) <= 0; flappy_W(17, 90) <= 0; flappy_W(17, 91) <= 0; flappy_W(17, 92) <= 0; flappy_W(17, 93) <= 0; flappy_W(17, 94) <= 0; flappy_W(17, 95) <= 0; flappy_W(17, 96) <= 0; flappy_W(17, 97) <= 0; flappy_W(17, 98) <= 0; flappy_W(17, 99) <= 0; flappy_W(17, 100) <= 0; flappy_W(17, 101) <= 0; flappy_W(17, 102) <= 0; flappy_W(17, 103) <= 0; flappy_W(17, 104) <= 0; flappy_W(17, 105) <= 0; flappy_W(17, 106) <= 0; flappy_W(17, 107) <= 0; flappy_W(17, 108) <= 0; flappy_W(17, 109) <= 0; flappy_W(17, 110) <= 0; flappy_W(17, 111) <= 0; flappy_W(17, 112) <= 0; flappy_W(17, 113) <= 0; flappy_W(17, 114) <= 1; flappy_W(17, 115) <= 1; flappy_W(17, 116) <= 1; flappy_W(17, 117) <= 1; flappy_W(17, 118) <= 1; flappy_W(17, 119) <= 1; flappy_W(17, 120) <= 1; flappy_W(17, 121) <= 1; flappy_W(17, 122) <= 1; flappy_W(17, 123) <= 1; flappy_W(17, 124) <= 1; flappy_W(17, 125) <= 1; flappy_W(17, 126) <= 0; flappy_W(17, 127) <= 0; flappy_W(17, 128) <= 0; flappy_W(17, 129) <= 0; flappy_W(17, 130) <= 0; flappy_W(17, 131) <= 0; flappy_W(17, 132) <= 1; flappy_W(17, 133) <= 1; flappy_W(17, 134) <= 1; flappy_W(17, 135) <= 1; flappy_W(17, 136) <= 1; flappy_W(17, 137) <= 1; flappy_W(17, 138) <= 1; flappy_W(17, 139) <= 1; flappy_W(17, 140) <= 1; flappy_W(17, 141) <= 1; flappy_W(17, 142) <= 1; flappy_W(17, 143) <= 1; flappy_W(17, 144) <= 0; flappy_W(17, 145) <= 0; flappy_W(17, 146) <= 0; flappy_W(17, 147) <= 0; flappy_W(17, 148) <= 0; flappy_W(17, 149) <= 0; flappy_W(17, 150) <= 0; flappy_W(17, 151) <= 0; flappy_W(17, 152) <= 0; flappy_W(17, 153) <= 0; flappy_W(17, 154) <= 0; flappy_W(17, 155) <= 0; flappy_W(17, 156) <= 0; flappy_W(17, 157) <= 0; flappy_W(17, 158) <= 0; flappy_W(17, 159) <= 0; flappy_W(17, 160) <= 0; flappy_W(17, 161) <= 0; flappy_W(17, 162) <= 0; flappy_W(17, 163) <= 0; flappy_W(17, 164) <= 0; flappy_W(17, 165) <= 0; flappy_W(17, 166) <= 0; flappy_W(17, 167) <= 0; flappy_W(17, 168) <= 1; flappy_W(17, 169) <= 1; flappy_W(17, 170) <= 1; flappy_W(17, 171) <= 1; flappy_W(17, 172) <= 1; flappy_W(17, 173) <= 1; flappy_W(17, 174) <= 1; flappy_W(17, 175) <= 1; flappy_W(17, 176) <= 1; flappy_W(17, 177) <= 1; flappy_W(17, 178) <= 1; flappy_W(17, 179) <= 1; flappy_W(17, 180) <= 0; flappy_W(17, 181) <= 0; flappy_W(17, 182) <= 0; flappy_W(17, 183) <= 0; flappy_W(17, 184) <= 0; flappy_W(17, 185) <= 0; flappy_W(17, 186) <= 0; flappy_W(17, 187) <= 0; flappy_W(17, 188) <= 0; flappy_W(17, 189) <= 0; flappy_W(17, 190) <= 0; flappy_W(17, 191) <= 0; flappy_W(17, 192) <= 1; flappy_W(17, 193) <= 1; flappy_W(17, 194) <= 1; flappy_W(17, 195) <= 1; flappy_W(17, 196) <= 1; flappy_W(17, 197) <= 1; flappy_W(17, 198) <= 1; flappy_W(17, 199) <= 1; flappy_W(17, 200) <= 1; flappy_W(17, 201) <= 1; flappy_W(17, 202) <= 1; flappy_W(17, 203) <= 1; flappy_W(17, 204) <= 0; flappy_W(17, 205) <= 0; flappy_W(17, 206) <= 0; flappy_W(17, 207) <= 0; flappy_W(17, 208) <= 0; flappy_W(17, 209) <= 0; flappy_W(17, 210) <= 0; flappy_W(17, 211) <= 0; flappy_W(17, 212) <= 0; flappy_W(17, 213) <= 0; flappy_W(17, 214) <= 0; flappy_W(17, 215) <= 0; flappy_W(17, 216) <= 0; flappy_W(17, 217) <= 0; flappy_W(17, 218) <= 0; flappy_W(17, 219) <= 0; flappy_W(17, 220) <= 0; flappy_W(17, 221) <= 0; flappy_W(17, 222) <= 1; flappy_W(17, 223) <= 1; flappy_W(17, 224) <= 1; flappy_W(17, 225) <= 1; flappy_W(17, 226) <= 1; flappy_W(17, 227) <= 1; flappy_W(17, 228) <= 1; flappy_W(17, 229) <= 1; flappy_W(17, 230) <= 1; flappy_W(17, 231) <= 1; flappy_W(17, 232) <= 1; flappy_W(17, 233) <= 1; flappy_W(17, 234) <= 0; flappy_W(17, 235) <= 0; flappy_W(17, 236) <= 0; flappy_W(17, 237) <= 0; flappy_W(17, 238) <= 0; flappy_W(17, 239) <= 0; flappy_W(17, 240) <= 0; flappy_W(17, 241) <= 0; flappy_W(17, 242) <= 0; flappy_W(17, 243) <= 0; flappy_W(17, 244) <= 0; flappy_W(17, 245) <= 0; flappy_W(17, 246) <= 1; flappy_W(17, 247) <= 1; flappy_W(17, 248) <= 1; flappy_W(17, 249) <= 1; flappy_W(17, 250) <= 1; flappy_W(17, 251) <= 1; flappy_W(17, 252) <= 1; flappy_W(17, 253) <= 1; flappy_W(17, 254) <= 1; flappy_W(17, 255) <= 1; flappy_W(17, 256) <= 1; flappy_W(17, 257) <= 1; flappy_W(17, 258) <= 0; flappy_W(17, 259) <= 0; flappy_W(17, 260) <= 0; flappy_W(17, 261) <= 0; flappy_W(17, 262) <= 0; flappy_W(17, 263) <= 0; flappy_W(17, 264) <= 0; flappy_W(17, 265) <= 0; flappy_W(17, 266) <= 0; flappy_W(17, 267) <= 0; flappy_W(17, 268) <= 0; flappy_W(17, 269) <= 0; flappy_W(17, 270) <= 1; flappy_W(17, 271) <= 1; flappy_W(17, 272) <= 1; flappy_W(17, 273) <= 1; flappy_W(17, 274) <= 1; flappy_W(17, 275) <= 1; flappy_W(17, 276) <= 1; flappy_W(17, 277) <= 1; flappy_W(17, 278) <= 1; flappy_W(17, 279) <= 1; flappy_W(17, 280) <= 1; flappy_W(17, 281) <= 1; flappy_W(17, 282) <= 0; flappy_W(17, 283) <= 0; flappy_W(17, 284) <= 0; flappy_W(17, 285) <= 0; flappy_W(17, 286) <= 0; flappy_W(17, 287) <= 0; flappy_W(17, 288) <= 0; flappy_W(17, 289) <= 0; flappy_W(17, 290) <= 0; flappy_W(17, 291) <= 0; flappy_W(17, 292) <= 0; flappy_W(17, 293) <= 0; flappy_W(17, 294) <= 0; flappy_W(17, 295) <= 0; flappy_W(17, 296) <= 0; flappy_W(17, 297) <= 0; flappy_W(17, 298) <= 0; flappy_W(17, 299) <= 0; flappy_W(17, 300) <= 0; flappy_W(17, 301) <= 0; flappy_W(17, 302) <= 0; flappy_W(17, 303) <= 0; flappy_W(17, 304) <= 0; flappy_W(17, 305) <= 0; flappy_W(17, 306) <= 1; flappy_W(17, 307) <= 1; flappy_W(17, 308) <= 1; flappy_W(17, 309) <= 1; flappy_W(17, 310) <= 1; flappy_W(17, 311) <= 1; flappy_W(17, 312) <= 1; flappy_W(17, 313) <= 1; flappy_W(17, 314) <= 1; flappy_W(17, 315) <= 1; flappy_W(17, 316) <= 1; flappy_W(17, 317) <= 1; flappy_W(17, 318) <= 0; flappy_W(17, 319) <= 0; flappy_W(17, 320) <= 0; flappy_W(17, 321) <= 0; flappy_W(17, 322) <= 0; flappy_W(17, 323) <= 0; flappy_W(17, 324) <= 0; flappy_W(17, 325) <= 0; flappy_W(17, 326) <= 0; flappy_W(17, 327) <= 0; flappy_W(17, 328) <= 0; flappy_W(17, 329) <= 0; flappy_W(17, 330) <= 0; flappy_W(17, 331) <= 0; flappy_W(17, 332) <= 0; flappy_W(17, 333) <= 0; flappy_W(17, 334) <= 0; flappy_W(17, 335) <= 0; flappy_W(17, 336) <= 0; flappy_W(17, 337) <= 0; flappy_W(17, 338) <= 0; flappy_W(17, 339) <= 0; flappy_W(17, 340) <= 0; flappy_W(17, 341) <= 0; flappy_W(17, 342) <= 0; flappy_W(17, 343) <= 0; flappy_W(17, 344) <= 0; flappy_W(17, 345) <= 0; flappy_W(17, 346) <= 0; flappy_W(17, 347) <= 0; flappy_W(17, 348) <= 0; flappy_W(17, 349) <= 0; flappy_W(17, 350) <= 0; flappy_W(17, 351) <= 0; flappy_W(17, 352) <= 0; flappy_W(17, 353) <= 0; flappy_W(17, 354) <= 0; flappy_W(17, 355) <= 0; flappy_W(17, 356) <= 0; flappy_W(17, 357) <= 0; flappy_W(17, 358) <= 0; flappy_W(17, 359) <= 0; flappy_W(17, 360) <= 0; flappy_W(17, 361) <= 0; flappy_W(17, 362) <= 0; flappy_W(17, 363) <= 0; flappy_W(17, 364) <= 0; flappy_W(17, 365) <= 0; flappy_W(17, 366) <= 0; flappy_W(17, 367) <= 0; flappy_W(17, 368) <= 0; flappy_W(17, 369) <= 0; flappy_W(17, 370) <= 0; flappy_W(17, 371) <= 0; flappy_W(17, 372) <= 0; flappy_W(17, 373) <= 0; flappy_W(17, 374) <= 0; flappy_W(17, 375) <= 0; flappy_W(17, 376) <= 0; flappy_W(17, 377) <= 0; flappy_W(17, 378) <= 0; flappy_W(17, 379) <= 0; flappy_W(17, 380) <= 0; flappy_W(17, 381) <= 0; flappy_W(17, 382) <= 0; flappy_W(17, 383) <= 0; flappy_W(17, 384) <= 0; flappy_W(17, 385) <= 0; flappy_W(17, 386) <= 0; flappy_W(17, 387) <= 0; flappy_W(17, 388) <= 0; flappy_W(17, 389) <= 0; flappy_W(17, 390) <= 0; flappy_W(17, 391) <= 0; flappy_W(17, 392) <= 0; flappy_W(17, 393) <= 0; flappy_W(17, 394) <= 0; flappy_W(17, 395) <= 0; flappy_W(17, 396) <= 0; flappy_W(17, 397) <= 0; flappy_W(17, 398) <= 0; flappy_W(17, 399) <= 0; flappy_W(17, 400) <= 0; flappy_W(17, 401) <= 0; flappy_W(17, 402) <= 1; flappy_W(17, 403) <= 1; flappy_W(17, 404) <= 1; flappy_W(17, 405) <= 1; flappy_W(17, 406) <= 1; flappy_W(17, 407) <= 1; flappy_W(17, 408) <= 1; flappy_W(17, 409) <= 1; flappy_W(17, 410) <= 1; flappy_W(17, 411) <= 1; flappy_W(17, 412) <= 1; flappy_W(17, 413) <= 1; flappy_W(17, 414) <= 0; flappy_W(17, 415) <= 0; flappy_W(17, 416) <= 0; flappy_W(17, 417) <= 0; flappy_W(17, 418) <= 0; flappy_W(17, 419) <= 0; flappy_W(17, 420) <= 0; flappy_W(17, 421) <= 0; flappy_W(17, 422) <= 0; flappy_W(17, 423) <= 0; flappy_W(17, 424) <= 0; flappy_W(17, 425) <= 0; flappy_W(17, 426) <= 1; flappy_W(17, 427) <= 1; flappy_W(17, 428) <= 1; flappy_W(17, 429) <= 1; flappy_W(17, 430) <= 1; flappy_W(17, 431) <= 1; flappy_W(17, 432) <= 1; flappy_W(17, 433) <= 1; flappy_W(17, 434) <= 1; flappy_W(17, 435) <= 1; flappy_W(17, 436) <= 1; flappy_W(17, 437) <= 1; flappy_W(17, 438) <= 0; flappy_W(17, 439) <= 0; flappy_W(17, 440) <= 0; flappy_W(17, 441) <= 0; flappy_W(17, 442) <= 0; flappy_W(17, 443) <= 0; flappy_W(17, 444) <= 0; flappy_W(17, 445) <= 0; flappy_W(17, 446) <= 0; flappy_W(17, 447) <= 0; flappy_W(17, 448) <= 0; flappy_W(17, 449) <= 0; flappy_W(17, 450) <= 0; flappy_W(17, 451) <= 0; flappy_W(17, 452) <= 0; flappy_W(17, 453) <= 0; flappy_W(17, 454) <= 0; flappy_W(17, 455) <= 0; flappy_W(17, 456) <= 0; flappy_W(17, 457) <= 0; flappy_W(17, 458) <= 0; flappy_W(17, 459) <= 0; flappy_W(17, 460) <= 0; flappy_W(17, 461) <= 0; flappy_W(17, 462) <= 0; flappy_W(17, 463) <= 0; flappy_W(17, 464) <= 0; flappy_W(17, 465) <= 0; flappy_W(17, 466) <= 0; flappy_W(17, 467) <= 0; flappy_W(17, 468) <= 1; flappy_W(17, 469) <= 1; flappy_W(17, 470) <= 1; flappy_W(17, 471) <= 1; flappy_W(17, 472) <= 1; flappy_W(17, 473) <= 1; flappy_W(17, 474) <= 1; flappy_W(17, 475) <= 1; flappy_W(17, 476) <= 1; flappy_W(17, 477) <= 1; flappy_W(17, 478) <= 1; flappy_W(17, 479) <= 1; flappy_W(17, 480) <= 0; flappy_W(17, 481) <= 0; flappy_W(17, 482) <= 0; flappy_W(17, 483) <= 0; flappy_W(17, 484) <= 0; flappy_W(17, 485) <= 0; flappy_W(17, 486) <= 0; flappy_W(17, 487) <= 0; flappy_W(17, 488) <= 0; flappy_W(17, 489) <= 0; flappy_W(17, 490) <= 0; flappy_W(17, 491) <= 0; flappy_W(17, 492) <= 0; flappy_W(17, 493) <= 0; flappy_W(17, 494) <= 0; flappy_W(17, 495) <= 0; flappy_W(17, 496) <= 0; flappy_W(17, 497) <= 0; flappy_W(17, 498) <= 0; flappy_W(17, 499) <= 0; flappy_W(17, 500) <= 0; flappy_W(17, 501) <= 0; flappy_W(17, 502) <= 0; flappy_W(17, 503) <= 0; flappy_W(17, 504) <= 0; flappy_W(17, 505) <= 0; flappy_W(17, 506) <= 0; flappy_W(17, 507) <= 0; flappy_W(17, 508) <= 0; flappy_W(17, 509) <= 0; flappy_W(17, 510) <= 1; flappy_W(17, 511) <= 1; flappy_W(17, 512) <= 1; flappy_W(17, 513) <= 1; flappy_W(17, 514) <= 1; flappy_W(17, 515) <= 1; flappy_W(17, 516) <= 1; flappy_W(17, 517) <= 1; flappy_W(17, 518) <= 1; flappy_W(17, 519) <= 1; flappy_W(17, 520) <= 1; flappy_W(17, 521) <= 1; flappy_W(17, 522) <= 0; flappy_W(17, 523) <= 0; flappy_W(17, 524) <= 0; flappy_W(17, 525) <= 0; flappy_W(17, 526) <= 0; flappy_W(17, 527) <= 0; flappy_W(17, 528) <= 0; flappy_W(17, 529) <= 0; flappy_W(17, 530) <= 0; flappy_W(17, 531) <= 0; flappy_W(17, 532) <= 0; flappy_W(17, 533) <= 0; flappy_W(17, 534) <= 1; flappy_W(17, 535) <= 1; flappy_W(17, 536) <= 1; flappy_W(17, 537) <= 1; flappy_W(17, 538) <= 1; flappy_W(17, 539) <= 1; flappy_W(17, 540) <= 1; flappy_W(17, 541) <= 1; flappy_W(17, 542) <= 1; flappy_W(17, 543) <= 1; flappy_W(17, 544) <= 1; flappy_W(17, 545) <= 1; flappy_W(17, 546) <= 0; flappy_W(17, 547) <= 0; flappy_W(17, 548) <= 0; flappy_W(17, 549) <= 0; flappy_W(17, 550) <= 0; flappy_W(17, 551) <= 0; flappy_W(17, 552) <= 0; flappy_W(17, 553) <= 0; flappy_W(17, 554) <= 0; flappy_W(17, 555) <= 0; flappy_W(17, 556) <= 0; flappy_W(17, 557) <= 0; flappy_W(17, 558) <= 0; flappy_W(17, 559) <= 0; flappy_W(17, 560) <= 0; flappy_W(17, 561) <= 0; flappy_W(17, 562) <= 0; flappy_W(17, 563) <= 0; flappy_W(17, 564) <= 1; flappy_W(17, 565) <= 1; flappy_W(17, 566) <= 1; flappy_W(17, 567) <= 1; flappy_W(17, 568) <= 1; flappy_W(17, 569) <= 1; flappy_W(17, 570) <= 1; flappy_W(17, 571) <= 1; flappy_W(17, 572) <= 1; flappy_W(17, 573) <= 1; flappy_W(17, 574) <= 1; flappy_W(17, 575) <= 1; flappy_W(17, 576) <= 0; flappy_W(17, 577) <= 0; flappy_W(17, 578) <= 0; flappy_W(17, 579) <= 0; flappy_W(17, 580) <= 0; flappy_W(17, 581) <= 0; flappy_W(17, 582) <= 0; flappy_W(17, 583) <= 0; flappy_W(17, 584) <= 0; flappy_W(17, 585) <= 0; flappy_W(17, 586) <= 0; flappy_W(17, 587) <= 0; flappy_W(17, 588) <= 1; flappy_W(17, 589) <= 1; flappy_W(17, 590) <= 1; flappy_W(17, 591) <= 1; flappy_W(17, 592) <= 1; flappy_W(17, 593) <= 1; 
flappy_W(18, 0) <= 0; flappy_W(18, 1) <= 0; flappy_W(18, 2) <= 0; flappy_W(18, 3) <= 0; flappy_W(18, 4) <= 0; flappy_W(18, 5) <= 0; flappy_W(18, 6) <= 1; flappy_W(18, 7) <= 1; flappy_W(18, 8) <= 1; flappy_W(18, 9) <= 1; flappy_W(18, 10) <= 1; flappy_W(18, 11) <= 1; flappy_W(18, 12) <= 1; flappy_W(18, 13) <= 1; flappy_W(18, 14) <= 1; flappy_W(18, 15) <= 1; flappy_W(18, 16) <= 1; flappy_W(18, 17) <= 1; flappy_W(18, 18) <= 0; flappy_W(18, 19) <= 0; flappy_W(18, 20) <= 0; flappy_W(18, 21) <= 0; flappy_W(18, 22) <= 0; flappy_W(18, 23) <= 0; flappy_W(18, 24) <= 1; flappy_W(18, 25) <= 1; flappy_W(18, 26) <= 1; flappy_W(18, 27) <= 1; flappy_W(18, 28) <= 1; flappy_W(18, 29) <= 1; flappy_W(18, 30) <= 0; flappy_W(18, 31) <= 0; flappy_W(18, 32) <= 0; flappy_W(18, 33) <= 0; flappy_W(18, 34) <= 0; flappy_W(18, 35) <= 0; flappy_W(18, 36) <= 0; flappy_W(18, 37) <= 0; flappy_W(18, 38) <= 0; flappy_W(18, 39) <= 0; flappy_W(18, 40) <= 0; flappy_W(18, 41) <= 0; flappy_W(18, 42) <= 0; flappy_W(18, 43) <= 0; flappy_W(18, 44) <= 0; flappy_W(18, 45) <= 0; flappy_W(18, 46) <= 0; flappy_W(18, 47) <= 0; flappy_W(18, 48) <= 0; flappy_W(18, 49) <= 0; flappy_W(18, 50) <= 0; flappy_W(18, 51) <= 0; flappy_W(18, 52) <= 0; flappy_W(18, 53) <= 0; flappy_W(18, 54) <= 0; flappy_W(18, 55) <= 0; flappy_W(18, 56) <= 0; flappy_W(18, 57) <= 0; flappy_W(18, 58) <= 0; flappy_W(18, 59) <= 0; flappy_W(18, 60) <= 1; flappy_W(18, 61) <= 1; flappy_W(18, 62) <= 1; flappy_W(18, 63) <= 1; flappy_W(18, 64) <= 1; flappy_W(18, 65) <= 1; flappy_W(18, 66) <= 1; flappy_W(18, 67) <= 1; flappy_W(18, 68) <= 1; flappy_W(18, 69) <= 1; flappy_W(18, 70) <= 1; flappy_W(18, 71) <= 1; flappy_W(18, 72) <= 0; flappy_W(18, 73) <= 0; flappy_W(18, 74) <= 0; flappy_W(18, 75) <= 0; flappy_W(18, 76) <= 0; flappy_W(18, 77) <= 0; flappy_W(18, 78) <= 0; flappy_W(18, 79) <= 0; flappy_W(18, 80) <= 0; flappy_W(18, 81) <= 0; flappy_W(18, 82) <= 0; flappy_W(18, 83) <= 0; flappy_W(18, 84) <= 0; flappy_W(18, 85) <= 0; flappy_W(18, 86) <= 0; flappy_W(18, 87) <= 0; flappy_W(18, 88) <= 0; flappy_W(18, 89) <= 0; flappy_W(18, 90) <= 0; flappy_W(18, 91) <= 0; flappy_W(18, 92) <= 0; flappy_W(18, 93) <= 0; flappy_W(18, 94) <= 0; flappy_W(18, 95) <= 0; flappy_W(18, 96) <= 0; flappy_W(18, 97) <= 0; flappy_W(18, 98) <= 0; flappy_W(18, 99) <= 0; flappy_W(18, 100) <= 0; flappy_W(18, 101) <= 0; flappy_W(18, 102) <= 0; flappy_W(18, 103) <= 0; flappy_W(18, 104) <= 0; flappy_W(18, 105) <= 0; flappy_W(18, 106) <= 0; flappy_W(18, 107) <= 0; flappy_W(18, 108) <= 1; flappy_W(18, 109) <= 1; flappy_W(18, 110) <= 1; flappy_W(18, 111) <= 1; flappy_W(18, 112) <= 1; flappy_W(18, 113) <= 1; flappy_W(18, 114) <= 1; flappy_W(18, 115) <= 1; flappy_W(18, 116) <= 1; flappy_W(18, 117) <= 1; flappy_W(18, 118) <= 1; flappy_W(18, 119) <= 1; flappy_W(18, 120) <= 0; flappy_W(18, 121) <= 0; flappy_W(18, 122) <= 0; flappy_W(18, 123) <= 0; flappy_W(18, 124) <= 0; flappy_W(18, 125) <= 0; flappy_W(18, 126) <= 0; flappy_W(18, 127) <= 0; flappy_W(18, 128) <= 0; flappy_W(18, 129) <= 0; flappy_W(18, 130) <= 0; flappy_W(18, 131) <= 0; flappy_W(18, 132) <= 0; flappy_W(18, 133) <= 0; flappy_W(18, 134) <= 0; flappy_W(18, 135) <= 0; flappy_W(18, 136) <= 0; flappy_W(18, 137) <= 0; flappy_W(18, 138) <= 1; flappy_W(18, 139) <= 1; flappy_W(18, 140) <= 1; flappy_W(18, 141) <= 1; flappy_W(18, 142) <= 1; flappy_W(18, 143) <= 1; flappy_W(18, 144) <= 1; flappy_W(18, 145) <= 1; flappy_W(18, 146) <= 1; flappy_W(18, 147) <= 1; flappy_W(18, 148) <= 1; flappy_W(18, 149) <= 1; flappy_W(18, 150) <= 0; flappy_W(18, 151) <= 0; flappy_W(18, 152) <= 0; flappy_W(18, 153) <= 0; flappy_W(18, 154) <= 0; flappy_W(18, 155) <= 0; flappy_W(18, 156) <= 0; flappy_W(18, 157) <= 0; flappy_W(18, 158) <= 0; flappy_W(18, 159) <= 0; flappy_W(18, 160) <= 0; flappy_W(18, 161) <= 0; flappy_W(18, 162) <= 0; flappy_W(18, 163) <= 0; flappy_W(18, 164) <= 0; flappy_W(18, 165) <= 0; flappy_W(18, 166) <= 0; flappy_W(18, 167) <= 0; flappy_W(18, 168) <= 1; flappy_W(18, 169) <= 1; flappy_W(18, 170) <= 1; flappy_W(18, 171) <= 1; flappy_W(18, 172) <= 1; flappy_W(18, 173) <= 1; flappy_W(18, 174) <= 1; flappy_W(18, 175) <= 1; flappy_W(18, 176) <= 1; flappy_W(18, 177) <= 1; flappy_W(18, 178) <= 1; flappy_W(18, 179) <= 1; flappy_W(18, 180) <= 0; flappy_W(18, 181) <= 0; flappy_W(18, 182) <= 0; flappy_W(18, 183) <= 0; flappy_W(18, 184) <= 0; flappy_W(18, 185) <= 0; flappy_W(18, 186) <= 0; flappy_W(18, 187) <= 0; flappy_W(18, 188) <= 0; flappy_W(18, 189) <= 0; flappy_W(18, 190) <= 0; flappy_W(18, 191) <= 0; flappy_W(18, 192) <= 1; flappy_W(18, 193) <= 1; flappy_W(18, 194) <= 1; flappy_W(18, 195) <= 1; flappy_W(18, 196) <= 1; flappy_W(18, 197) <= 1; flappy_W(18, 198) <= 1; flappy_W(18, 199) <= 1; flappy_W(18, 200) <= 1; flappy_W(18, 201) <= 1; flappy_W(18, 202) <= 1; flappy_W(18, 203) <= 1; flappy_W(18, 204) <= 0; flappy_W(18, 205) <= 0; flappy_W(18, 206) <= 0; flappy_W(18, 207) <= 0; flappy_W(18, 208) <= 0; flappy_W(18, 209) <= 0; flappy_W(18, 210) <= 0; flappy_W(18, 211) <= 0; flappy_W(18, 212) <= 0; flappy_W(18, 213) <= 0; flappy_W(18, 214) <= 0; flappy_W(18, 215) <= 0; flappy_W(18, 216) <= 0; flappy_W(18, 217) <= 0; flappy_W(18, 218) <= 0; flappy_W(18, 219) <= 0; flappy_W(18, 220) <= 0; flappy_W(18, 221) <= 0; flappy_W(18, 222) <= 1; flappy_W(18, 223) <= 1; flappy_W(18, 224) <= 1; flappy_W(18, 225) <= 1; flappy_W(18, 226) <= 1; flappy_W(18, 227) <= 1; flappy_W(18, 228) <= 1; flappy_W(18, 229) <= 1; flappy_W(18, 230) <= 1; flappy_W(18, 231) <= 1; flappy_W(18, 232) <= 1; flappy_W(18, 233) <= 1; flappy_W(18, 234) <= 0; flappy_W(18, 235) <= 0; flappy_W(18, 236) <= 0; flappy_W(18, 237) <= 0; flappy_W(18, 238) <= 0; flappy_W(18, 239) <= 0; flappy_W(18, 240) <= 0; flappy_W(18, 241) <= 0; flappy_W(18, 242) <= 0; flappy_W(18, 243) <= 0; flappy_W(18, 244) <= 0; flappy_W(18, 245) <= 0; flappy_W(18, 246) <= 1; flappy_W(18, 247) <= 1; flappy_W(18, 248) <= 1; flappy_W(18, 249) <= 1; flappy_W(18, 250) <= 1; flappy_W(18, 251) <= 1; flappy_W(18, 252) <= 1; flappy_W(18, 253) <= 1; flappy_W(18, 254) <= 1; flappy_W(18, 255) <= 1; flappy_W(18, 256) <= 1; flappy_W(18, 257) <= 1; flappy_W(18, 258) <= 0; flappy_W(18, 259) <= 0; flappy_W(18, 260) <= 0; flappy_W(18, 261) <= 0; flappy_W(18, 262) <= 0; flappy_W(18, 263) <= 0; flappy_W(18, 264) <= 0; flappy_W(18, 265) <= 0; flappy_W(18, 266) <= 0; flappy_W(18, 267) <= 0; flappy_W(18, 268) <= 0; flappy_W(18, 269) <= 0; flappy_W(18, 270) <= 0; flappy_W(18, 271) <= 0; flappy_W(18, 272) <= 0; flappy_W(18, 273) <= 0; flappy_W(18, 274) <= 0; flappy_W(18, 275) <= 0; flappy_W(18, 276) <= 1; flappy_W(18, 277) <= 1; flappy_W(18, 278) <= 1; flappy_W(18, 279) <= 1; flappy_W(18, 280) <= 1; flappy_W(18, 281) <= 1; flappy_W(18, 282) <= 1; flappy_W(18, 283) <= 1; flappy_W(18, 284) <= 1; flappy_W(18, 285) <= 1; flappy_W(18, 286) <= 1; flappy_W(18, 287) <= 1; flappy_W(18, 288) <= 0; flappy_W(18, 289) <= 0; flappy_W(18, 290) <= 0; flappy_W(18, 291) <= 0; flappy_W(18, 292) <= 0; flappy_W(18, 293) <= 0; flappy_W(18, 294) <= 0; flappy_W(18, 295) <= 0; flappy_W(18, 296) <= 0; flappy_W(18, 297) <= 0; flappy_W(18, 298) <= 0; flappy_W(18, 299) <= 0; flappy_W(18, 300) <= 1; flappy_W(18, 301) <= 1; flappy_W(18, 302) <= 1; flappy_W(18, 303) <= 1; flappy_W(18, 304) <= 1; flappy_W(18, 305) <= 1; flappy_W(18, 306) <= 1; flappy_W(18, 307) <= 1; flappy_W(18, 308) <= 1; flappy_W(18, 309) <= 1; flappy_W(18, 310) <= 1; flappy_W(18, 311) <= 1; flappy_W(18, 312) <= 0; flappy_W(18, 313) <= 0; flappy_W(18, 314) <= 0; flappy_W(18, 315) <= 0; flappy_W(18, 316) <= 0; flappy_W(18, 317) <= 0; flappy_W(18, 318) <= 0; flappy_W(18, 319) <= 0; flappy_W(18, 320) <= 0; flappy_W(18, 321) <= 0; flappy_W(18, 322) <= 0; flappy_W(18, 323) <= 0; flappy_W(18, 324) <= 0; flappy_W(18, 325) <= 0; flappy_W(18, 326) <= 0; flappy_W(18, 327) <= 0; flappy_W(18, 328) <= 0; flappy_W(18, 329) <= 0; flappy_W(18, 330) <= 0; flappy_W(18, 331) <= 0; flappy_W(18, 332) <= 0; flappy_W(18, 333) <= 0; flappy_W(18, 334) <= 0; flappy_W(18, 335) <= 0; flappy_W(18, 336) <= 0; flappy_W(18, 337) <= 0; flappy_W(18, 338) <= 0; flappy_W(18, 339) <= 0; flappy_W(18, 340) <= 0; flappy_W(18, 341) <= 0; flappy_W(18, 342) <= 0; flappy_W(18, 343) <= 0; flappy_W(18, 344) <= 0; flappy_W(18, 345) <= 0; flappy_W(18, 346) <= 0; flappy_W(18, 347) <= 0; flappy_W(18, 348) <= 0; flappy_W(18, 349) <= 0; flappy_W(18, 350) <= 0; flappy_W(18, 351) <= 0; flappy_W(18, 352) <= 0; flappy_W(18, 353) <= 0; flappy_W(18, 354) <= 0; flappy_W(18, 355) <= 0; flappy_W(18, 356) <= 0; flappy_W(18, 357) <= 0; flappy_W(18, 358) <= 0; flappy_W(18, 359) <= 0; flappy_W(18, 360) <= 0; flappy_W(18, 361) <= 0; flappy_W(18, 362) <= 0; flappy_W(18, 363) <= 0; flappy_W(18, 364) <= 0; flappy_W(18, 365) <= 0; flappy_W(18, 366) <= 0; flappy_W(18, 367) <= 0; flappy_W(18, 368) <= 0; flappy_W(18, 369) <= 0; flappy_W(18, 370) <= 0; flappy_W(18, 371) <= 0; flappy_W(18, 372) <= 0; flappy_W(18, 373) <= 0; flappy_W(18, 374) <= 0; flappy_W(18, 375) <= 0; flappy_W(18, 376) <= 0; flappy_W(18, 377) <= 0; flappy_W(18, 378) <= 0; flappy_W(18, 379) <= 0; flappy_W(18, 380) <= 0; flappy_W(18, 381) <= 0; flappy_W(18, 382) <= 0; flappy_W(18, 383) <= 0; flappy_W(18, 384) <= 0; flappy_W(18, 385) <= 0; flappy_W(18, 386) <= 0; flappy_W(18, 387) <= 0; flappy_W(18, 388) <= 0; flappy_W(18, 389) <= 0; flappy_W(18, 390) <= 0; flappy_W(18, 391) <= 0; flappy_W(18, 392) <= 0; flappy_W(18, 393) <= 0; flappy_W(18, 394) <= 0; flappy_W(18, 395) <= 0; flappy_W(18, 396) <= 0; flappy_W(18, 397) <= 0; flappy_W(18, 398) <= 0; flappy_W(18, 399) <= 0; flappy_W(18, 400) <= 0; flappy_W(18, 401) <= 0; flappy_W(18, 402) <= 1; flappy_W(18, 403) <= 1; flappy_W(18, 404) <= 1; flappy_W(18, 405) <= 1; flappy_W(18, 406) <= 1; flappy_W(18, 407) <= 1; flappy_W(18, 408) <= 1; flappy_W(18, 409) <= 1; flappy_W(18, 410) <= 1; flappy_W(18, 411) <= 1; flappy_W(18, 412) <= 1; flappy_W(18, 413) <= 1; flappy_W(18, 414) <= 0; flappy_W(18, 415) <= 0; flappy_W(18, 416) <= 0; flappy_W(18, 417) <= 0; flappy_W(18, 418) <= 0; flappy_W(18, 419) <= 0; flappy_W(18, 420) <= 0; flappy_W(18, 421) <= 0; flappy_W(18, 422) <= 0; flappy_W(18, 423) <= 0; flappy_W(18, 424) <= 0; flappy_W(18, 425) <= 0; flappy_W(18, 426) <= 1; flappy_W(18, 427) <= 1; flappy_W(18, 428) <= 1; flappy_W(18, 429) <= 1; flappy_W(18, 430) <= 1; flappy_W(18, 431) <= 1; flappy_W(18, 432) <= 1; flappy_W(18, 433) <= 1; flappy_W(18, 434) <= 1; flappy_W(18, 435) <= 1; flappy_W(18, 436) <= 1; flappy_W(18, 437) <= 1; flappy_W(18, 438) <= 0; flappy_W(18, 439) <= 0; flappy_W(18, 440) <= 0; flappy_W(18, 441) <= 0; flappy_W(18, 442) <= 0; flappy_W(18, 443) <= 0; flappy_W(18, 444) <= 0; flappy_W(18, 445) <= 0; flappy_W(18, 446) <= 0; flappy_W(18, 447) <= 0; flappy_W(18, 448) <= 0; flappy_W(18, 449) <= 0; flappy_W(18, 450) <= 0; flappy_W(18, 451) <= 0; flappy_W(18, 452) <= 0; flappy_W(18, 453) <= 0; flappy_W(18, 454) <= 0; flappy_W(18, 455) <= 0; flappy_W(18, 456) <= 0; flappy_W(18, 457) <= 0; flappy_W(18, 458) <= 0; flappy_W(18, 459) <= 0; flappy_W(18, 460) <= 0; flappy_W(18, 461) <= 0; flappy_W(18, 462) <= 0; flappy_W(18, 463) <= 0; flappy_W(18, 464) <= 0; flappy_W(18, 465) <= 0; flappy_W(18, 466) <= 0; flappy_W(18, 467) <= 0; flappy_W(18, 468) <= 1; flappy_W(18, 469) <= 1; flappy_W(18, 470) <= 1; flappy_W(18, 471) <= 1; flappy_W(18, 472) <= 1; flappy_W(18, 473) <= 1; flappy_W(18, 474) <= 1; flappy_W(18, 475) <= 1; flappy_W(18, 476) <= 1; flappy_W(18, 477) <= 1; flappy_W(18, 478) <= 1; flappy_W(18, 479) <= 1; flappy_W(18, 480) <= 0; flappy_W(18, 481) <= 0; flappy_W(18, 482) <= 0; flappy_W(18, 483) <= 0; flappy_W(18, 484) <= 0; flappy_W(18, 485) <= 0; flappy_W(18, 486) <= 0; flappy_W(18, 487) <= 0; flappy_W(18, 488) <= 0; flappy_W(18, 489) <= 0; flappy_W(18, 490) <= 0; flappy_W(18, 491) <= 0; flappy_W(18, 492) <= 0; flappy_W(18, 493) <= 0; flappy_W(18, 494) <= 0; flappy_W(18, 495) <= 0; flappy_W(18, 496) <= 0; flappy_W(18, 497) <= 0; flappy_W(18, 498) <= 0; flappy_W(18, 499) <= 0; flappy_W(18, 500) <= 0; flappy_W(18, 501) <= 0; flappy_W(18, 502) <= 0; flappy_W(18, 503) <= 0; flappy_W(18, 504) <= 0; flappy_W(18, 505) <= 0; flappy_W(18, 506) <= 0; flappy_W(18, 507) <= 0; flappy_W(18, 508) <= 0; flappy_W(18, 509) <= 0; flappy_W(18, 510) <= 1; flappy_W(18, 511) <= 1; flappy_W(18, 512) <= 1; flappy_W(18, 513) <= 1; flappy_W(18, 514) <= 1; flappy_W(18, 515) <= 1; flappy_W(18, 516) <= 1; flappy_W(18, 517) <= 1; flappy_W(18, 518) <= 1; flappy_W(18, 519) <= 1; flappy_W(18, 520) <= 1; flappy_W(18, 521) <= 1; flappy_W(18, 522) <= 0; flappy_W(18, 523) <= 0; flappy_W(18, 524) <= 0; flappy_W(18, 525) <= 0; flappy_W(18, 526) <= 0; flappy_W(18, 527) <= 0; flappy_W(18, 528) <= 0; flappy_W(18, 529) <= 0; flappy_W(18, 530) <= 0; flappy_W(18, 531) <= 0; flappy_W(18, 532) <= 0; flappy_W(18, 533) <= 0; flappy_W(18, 534) <= 1; flappy_W(18, 535) <= 1; flappy_W(18, 536) <= 1; flappy_W(18, 537) <= 1; flappy_W(18, 538) <= 1; flappy_W(18, 539) <= 1; flappy_W(18, 540) <= 1; flappy_W(18, 541) <= 1; flappy_W(18, 542) <= 1; flappy_W(18, 543) <= 1; flappy_W(18, 544) <= 1; flappy_W(18, 545) <= 1; flappy_W(18, 546) <= 0; flappy_W(18, 547) <= 0; flappy_W(18, 548) <= 0; flappy_W(18, 549) <= 0; flappy_W(18, 550) <= 0; flappy_W(18, 551) <= 0; flappy_W(18, 552) <= 0; flappy_W(18, 553) <= 0; flappy_W(18, 554) <= 0; flappy_W(18, 555) <= 0; flappy_W(18, 556) <= 0; flappy_W(18, 557) <= 0; flappy_W(18, 558) <= 0; flappy_W(18, 559) <= 0; flappy_W(18, 560) <= 0; flappy_W(18, 561) <= 0; flappy_W(18, 562) <= 0; flappy_W(18, 563) <= 0; flappy_W(18, 564) <= 1; flappy_W(18, 565) <= 1; flappy_W(18, 566) <= 1; flappy_W(18, 567) <= 1; flappy_W(18, 568) <= 1; flappy_W(18, 569) <= 1; flappy_W(18, 570) <= 1; flappy_W(18, 571) <= 1; flappy_W(18, 572) <= 1; flappy_W(18, 573) <= 1; flappy_W(18, 574) <= 1; flappy_W(18, 575) <= 1; flappy_W(18, 576) <= 0; flappy_W(18, 577) <= 0; flappy_W(18, 578) <= 0; flappy_W(18, 579) <= 0; flappy_W(18, 580) <= 0; flappy_W(18, 581) <= 0; flappy_W(18, 582) <= 0; flappy_W(18, 583) <= 0; flappy_W(18, 584) <= 0; flappy_W(18, 585) <= 0; flappy_W(18, 586) <= 0; flappy_W(18, 587) <= 0; flappy_W(18, 588) <= 1; flappy_W(18, 589) <= 1; flappy_W(18, 590) <= 1; flappy_W(18, 591) <= 1; flappy_W(18, 592) <= 1; flappy_W(18, 593) <= 1; 
flappy_W(19, 0) <= 0; flappy_W(19, 1) <= 0; flappy_W(19, 2) <= 0; flappy_W(19, 3) <= 0; flappy_W(19, 4) <= 0; flappy_W(19, 5) <= 0; flappy_W(19, 6) <= 1; flappy_W(19, 7) <= 1; flappy_W(19, 8) <= 1; flappy_W(19, 9) <= 1; flappy_W(19, 10) <= 1; flappy_W(19, 11) <= 1; flappy_W(19, 12) <= 1; flappy_W(19, 13) <= 1; flappy_W(19, 14) <= 1; flappy_W(19, 15) <= 1; flappy_W(19, 16) <= 1; flappy_W(19, 17) <= 1; flappy_W(19, 18) <= 0; flappy_W(19, 19) <= 0; flappy_W(19, 20) <= 0; flappy_W(19, 21) <= 0; flappy_W(19, 22) <= 0; flappy_W(19, 23) <= 0; flappy_W(19, 24) <= 1; flappy_W(19, 25) <= 1; flappy_W(19, 26) <= 1; flappy_W(19, 27) <= 1; flappy_W(19, 28) <= 1; flappy_W(19, 29) <= 1; flappy_W(19, 30) <= 0; flappy_W(19, 31) <= 0; flappy_W(19, 32) <= 0; flappy_W(19, 33) <= 0; flappy_W(19, 34) <= 0; flappy_W(19, 35) <= 0; flappy_W(19, 36) <= 0; flappy_W(19, 37) <= 0; flappy_W(19, 38) <= 0; flappy_W(19, 39) <= 0; flappy_W(19, 40) <= 0; flappy_W(19, 41) <= 0; flappy_W(19, 42) <= 0; flappy_W(19, 43) <= 0; flappy_W(19, 44) <= 0; flappy_W(19, 45) <= 0; flappy_W(19, 46) <= 0; flappy_W(19, 47) <= 0; flappy_W(19, 48) <= 0; flappy_W(19, 49) <= 0; flappy_W(19, 50) <= 0; flappy_W(19, 51) <= 0; flappy_W(19, 52) <= 0; flappy_W(19, 53) <= 0; flappy_W(19, 54) <= 0; flappy_W(19, 55) <= 0; flappy_W(19, 56) <= 0; flappy_W(19, 57) <= 0; flappy_W(19, 58) <= 0; flappy_W(19, 59) <= 0; flappy_W(19, 60) <= 1; flappy_W(19, 61) <= 1; flappy_W(19, 62) <= 1; flappy_W(19, 63) <= 1; flappy_W(19, 64) <= 1; flappy_W(19, 65) <= 1; flappy_W(19, 66) <= 1; flappy_W(19, 67) <= 1; flappy_W(19, 68) <= 1; flappy_W(19, 69) <= 1; flappy_W(19, 70) <= 1; flappy_W(19, 71) <= 1; flappy_W(19, 72) <= 0; flappy_W(19, 73) <= 0; flappy_W(19, 74) <= 0; flappy_W(19, 75) <= 0; flappy_W(19, 76) <= 0; flappy_W(19, 77) <= 0; flappy_W(19, 78) <= 0; flappy_W(19, 79) <= 0; flappy_W(19, 80) <= 0; flappy_W(19, 81) <= 0; flappy_W(19, 82) <= 0; flappy_W(19, 83) <= 0; flappy_W(19, 84) <= 0; flappy_W(19, 85) <= 0; flappy_W(19, 86) <= 0; flappy_W(19, 87) <= 0; flappy_W(19, 88) <= 0; flappy_W(19, 89) <= 0; flappy_W(19, 90) <= 0; flappy_W(19, 91) <= 0; flappy_W(19, 92) <= 0; flappy_W(19, 93) <= 0; flappy_W(19, 94) <= 0; flappy_W(19, 95) <= 0; flappy_W(19, 96) <= 0; flappy_W(19, 97) <= 0; flappy_W(19, 98) <= 0; flappy_W(19, 99) <= 0; flappy_W(19, 100) <= 0; flappy_W(19, 101) <= 0; flappy_W(19, 102) <= 0; flappy_W(19, 103) <= 0; flappy_W(19, 104) <= 0; flappy_W(19, 105) <= 0; flappy_W(19, 106) <= 0; flappy_W(19, 107) <= 0; flappy_W(19, 108) <= 1; flappy_W(19, 109) <= 1; flappy_W(19, 110) <= 1; flappy_W(19, 111) <= 1; flappy_W(19, 112) <= 1; flappy_W(19, 113) <= 1; flappy_W(19, 114) <= 1; flappy_W(19, 115) <= 1; flappy_W(19, 116) <= 1; flappy_W(19, 117) <= 1; flappy_W(19, 118) <= 1; flappy_W(19, 119) <= 1; flappy_W(19, 120) <= 0; flappy_W(19, 121) <= 0; flappy_W(19, 122) <= 0; flappy_W(19, 123) <= 0; flappy_W(19, 124) <= 0; flappy_W(19, 125) <= 0; flappy_W(19, 126) <= 0; flappy_W(19, 127) <= 0; flappy_W(19, 128) <= 0; flappy_W(19, 129) <= 0; flappy_W(19, 130) <= 0; flappy_W(19, 131) <= 0; flappy_W(19, 132) <= 0; flappy_W(19, 133) <= 0; flappy_W(19, 134) <= 0; flappy_W(19, 135) <= 0; flappy_W(19, 136) <= 0; flappy_W(19, 137) <= 0; flappy_W(19, 138) <= 1; flappy_W(19, 139) <= 1; flappy_W(19, 140) <= 1; flappy_W(19, 141) <= 1; flappy_W(19, 142) <= 1; flappy_W(19, 143) <= 1; flappy_W(19, 144) <= 1; flappy_W(19, 145) <= 1; flappy_W(19, 146) <= 1; flappy_W(19, 147) <= 1; flappy_W(19, 148) <= 1; flappy_W(19, 149) <= 1; flappy_W(19, 150) <= 0; flappy_W(19, 151) <= 0; flappy_W(19, 152) <= 0; flappy_W(19, 153) <= 0; flappy_W(19, 154) <= 0; flappy_W(19, 155) <= 0; flappy_W(19, 156) <= 0; flappy_W(19, 157) <= 0; flappy_W(19, 158) <= 0; flappy_W(19, 159) <= 0; flappy_W(19, 160) <= 0; flappy_W(19, 161) <= 0; flappy_W(19, 162) <= 0; flappy_W(19, 163) <= 0; flappy_W(19, 164) <= 0; flappy_W(19, 165) <= 0; flappy_W(19, 166) <= 0; flappy_W(19, 167) <= 0; flappy_W(19, 168) <= 1; flappy_W(19, 169) <= 1; flappy_W(19, 170) <= 1; flappy_W(19, 171) <= 1; flappy_W(19, 172) <= 1; flappy_W(19, 173) <= 1; flappy_W(19, 174) <= 1; flappy_W(19, 175) <= 1; flappy_W(19, 176) <= 1; flappy_W(19, 177) <= 1; flappy_W(19, 178) <= 1; flappy_W(19, 179) <= 1; flappy_W(19, 180) <= 0; flappy_W(19, 181) <= 0; flappy_W(19, 182) <= 0; flappy_W(19, 183) <= 0; flappy_W(19, 184) <= 0; flappy_W(19, 185) <= 0; flappy_W(19, 186) <= 0; flappy_W(19, 187) <= 0; flappy_W(19, 188) <= 0; flappy_W(19, 189) <= 0; flappy_W(19, 190) <= 0; flappy_W(19, 191) <= 0; flappy_W(19, 192) <= 1; flappy_W(19, 193) <= 1; flappy_W(19, 194) <= 1; flappy_W(19, 195) <= 1; flappy_W(19, 196) <= 1; flappy_W(19, 197) <= 1; flappy_W(19, 198) <= 1; flappy_W(19, 199) <= 1; flappy_W(19, 200) <= 1; flappy_W(19, 201) <= 1; flappy_W(19, 202) <= 1; flappy_W(19, 203) <= 1; flappy_W(19, 204) <= 0; flappy_W(19, 205) <= 0; flappy_W(19, 206) <= 0; flappy_W(19, 207) <= 0; flappy_W(19, 208) <= 0; flappy_W(19, 209) <= 0; flappy_W(19, 210) <= 0; flappy_W(19, 211) <= 0; flappy_W(19, 212) <= 0; flappy_W(19, 213) <= 0; flappy_W(19, 214) <= 0; flappy_W(19, 215) <= 0; flappy_W(19, 216) <= 0; flappy_W(19, 217) <= 0; flappy_W(19, 218) <= 0; flappy_W(19, 219) <= 0; flappy_W(19, 220) <= 0; flappy_W(19, 221) <= 0; flappy_W(19, 222) <= 1; flappy_W(19, 223) <= 1; flappy_W(19, 224) <= 1; flappy_W(19, 225) <= 1; flappy_W(19, 226) <= 1; flappy_W(19, 227) <= 1; flappy_W(19, 228) <= 1; flappy_W(19, 229) <= 1; flappy_W(19, 230) <= 1; flappy_W(19, 231) <= 1; flappy_W(19, 232) <= 1; flappy_W(19, 233) <= 1; flappy_W(19, 234) <= 0; flappy_W(19, 235) <= 0; flappy_W(19, 236) <= 0; flappy_W(19, 237) <= 0; flappy_W(19, 238) <= 0; flappy_W(19, 239) <= 0; flappy_W(19, 240) <= 0; flappy_W(19, 241) <= 0; flappy_W(19, 242) <= 0; flappy_W(19, 243) <= 0; flappy_W(19, 244) <= 0; flappy_W(19, 245) <= 0; flappy_W(19, 246) <= 1; flappy_W(19, 247) <= 1; flappy_W(19, 248) <= 1; flappy_W(19, 249) <= 1; flappy_W(19, 250) <= 1; flappy_W(19, 251) <= 1; flappy_W(19, 252) <= 1; flappy_W(19, 253) <= 1; flappy_W(19, 254) <= 1; flappy_W(19, 255) <= 1; flappy_W(19, 256) <= 1; flappy_W(19, 257) <= 1; flappy_W(19, 258) <= 0; flappy_W(19, 259) <= 0; flappy_W(19, 260) <= 0; flappy_W(19, 261) <= 0; flappy_W(19, 262) <= 0; flappy_W(19, 263) <= 0; flappy_W(19, 264) <= 0; flappy_W(19, 265) <= 0; flappy_W(19, 266) <= 0; flappy_W(19, 267) <= 0; flappy_W(19, 268) <= 0; flappy_W(19, 269) <= 0; flappy_W(19, 270) <= 0; flappy_W(19, 271) <= 0; flappy_W(19, 272) <= 0; flappy_W(19, 273) <= 0; flappy_W(19, 274) <= 0; flappy_W(19, 275) <= 0; flappy_W(19, 276) <= 1; flappy_W(19, 277) <= 1; flappy_W(19, 278) <= 1; flappy_W(19, 279) <= 1; flappy_W(19, 280) <= 1; flappy_W(19, 281) <= 1; flappy_W(19, 282) <= 1; flappy_W(19, 283) <= 1; flappy_W(19, 284) <= 1; flappy_W(19, 285) <= 1; flappy_W(19, 286) <= 1; flappy_W(19, 287) <= 1; flappy_W(19, 288) <= 0; flappy_W(19, 289) <= 0; flappy_W(19, 290) <= 0; flappy_W(19, 291) <= 0; flappy_W(19, 292) <= 0; flappy_W(19, 293) <= 0; flappy_W(19, 294) <= 0; flappy_W(19, 295) <= 0; flappy_W(19, 296) <= 0; flappy_W(19, 297) <= 0; flappy_W(19, 298) <= 0; flappy_W(19, 299) <= 0; flappy_W(19, 300) <= 1; flappy_W(19, 301) <= 1; flappy_W(19, 302) <= 1; flappy_W(19, 303) <= 1; flappy_W(19, 304) <= 1; flappy_W(19, 305) <= 1; flappy_W(19, 306) <= 1; flappy_W(19, 307) <= 1; flappy_W(19, 308) <= 1; flappy_W(19, 309) <= 1; flappy_W(19, 310) <= 1; flappy_W(19, 311) <= 1; flappy_W(19, 312) <= 0; flappy_W(19, 313) <= 0; flappy_W(19, 314) <= 0; flappy_W(19, 315) <= 0; flappy_W(19, 316) <= 0; flappy_W(19, 317) <= 0; flappy_W(19, 318) <= 0; flappy_W(19, 319) <= 0; flappy_W(19, 320) <= 0; flappy_W(19, 321) <= 0; flappy_W(19, 322) <= 0; flappy_W(19, 323) <= 0; flappy_W(19, 324) <= 0; flappy_W(19, 325) <= 0; flappy_W(19, 326) <= 0; flappy_W(19, 327) <= 0; flappy_W(19, 328) <= 0; flappy_W(19, 329) <= 0; flappy_W(19, 330) <= 0; flappy_W(19, 331) <= 0; flappy_W(19, 332) <= 0; flappy_W(19, 333) <= 0; flappy_W(19, 334) <= 0; flappy_W(19, 335) <= 0; flappy_W(19, 336) <= 0; flappy_W(19, 337) <= 0; flappy_W(19, 338) <= 0; flappy_W(19, 339) <= 0; flappy_W(19, 340) <= 0; flappy_W(19, 341) <= 0; flappy_W(19, 342) <= 0; flappy_W(19, 343) <= 0; flappy_W(19, 344) <= 0; flappy_W(19, 345) <= 0; flappy_W(19, 346) <= 0; flappy_W(19, 347) <= 0; flappy_W(19, 348) <= 0; flappy_W(19, 349) <= 0; flappy_W(19, 350) <= 0; flappy_W(19, 351) <= 0; flappy_W(19, 352) <= 0; flappy_W(19, 353) <= 0; flappy_W(19, 354) <= 0; flappy_W(19, 355) <= 0; flappy_W(19, 356) <= 0; flappy_W(19, 357) <= 0; flappy_W(19, 358) <= 0; flappy_W(19, 359) <= 0; flappy_W(19, 360) <= 0; flappy_W(19, 361) <= 0; flappy_W(19, 362) <= 0; flappy_W(19, 363) <= 0; flappy_W(19, 364) <= 0; flappy_W(19, 365) <= 0; flappy_W(19, 366) <= 0; flappy_W(19, 367) <= 0; flappy_W(19, 368) <= 0; flappy_W(19, 369) <= 0; flappy_W(19, 370) <= 0; flappy_W(19, 371) <= 0; flappy_W(19, 372) <= 0; flappy_W(19, 373) <= 0; flappy_W(19, 374) <= 0; flappy_W(19, 375) <= 0; flappy_W(19, 376) <= 0; flappy_W(19, 377) <= 0; flappy_W(19, 378) <= 0; flappy_W(19, 379) <= 0; flappy_W(19, 380) <= 0; flappy_W(19, 381) <= 0; flappy_W(19, 382) <= 0; flappy_W(19, 383) <= 0; flappy_W(19, 384) <= 0; flappy_W(19, 385) <= 0; flappy_W(19, 386) <= 0; flappy_W(19, 387) <= 0; flappy_W(19, 388) <= 0; flappy_W(19, 389) <= 0; flappy_W(19, 390) <= 0; flappy_W(19, 391) <= 0; flappy_W(19, 392) <= 0; flappy_W(19, 393) <= 0; flappy_W(19, 394) <= 0; flappy_W(19, 395) <= 0; flappy_W(19, 396) <= 0; flappy_W(19, 397) <= 0; flappy_W(19, 398) <= 0; flappy_W(19, 399) <= 0; flappy_W(19, 400) <= 0; flappy_W(19, 401) <= 0; flappy_W(19, 402) <= 1; flappy_W(19, 403) <= 1; flappy_W(19, 404) <= 1; flappy_W(19, 405) <= 1; flappy_W(19, 406) <= 1; flappy_W(19, 407) <= 1; flappy_W(19, 408) <= 1; flappy_W(19, 409) <= 1; flappy_W(19, 410) <= 1; flappy_W(19, 411) <= 1; flappy_W(19, 412) <= 1; flappy_W(19, 413) <= 1; flappy_W(19, 414) <= 0; flappy_W(19, 415) <= 0; flappy_W(19, 416) <= 0; flappy_W(19, 417) <= 0; flappy_W(19, 418) <= 0; flappy_W(19, 419) <= 0; flappy_W(19, 420) <= 0; flappy_W(19, 421) <= 0; flappy_W(19, 422) <= 0; flappy_W(19, 423) <= 0; flappy_W(19, 424) <= 0; flappy_W(19, 425) <= 0; flappy_W(19, 426) <= 1; flappy_W(19, 427) <= 1; flappy_W(19, 428) <= 1; flappy_W(19, 429) <= 1; flappy_W(19, 430) <= 1; flappy_W(19, 431) <= 1; flappy_W(19, 432) <= 1; flappy_W(19, 433) <= 1; flappy_W(19, 434) <= 1; flappy_W(19, 435) <= 1; flappy_W(19, 436) <= 1; flappy_W(19, 437) <= 1; flappy_W(19, 438) <= 0; flappy_W(19, 439) <= 0; flappy_W(19, 440) <= 0; flappy_W(19, 441) <= 0; flappy_W(19, 442) <= 0; flappy_W(19, 443) <= 0; flappy_W(19, 444) <= 0; flappy_W(19, 445) <= 0; flappy_W(19, 446) <= 0; flappy_W(19, 447) <= 0; flappy_W(19, 448) <= 0; flappy_W(19, 449) <= 0; flappy_W(19, 450) <= 0; flappy_W(19, 451) <= 0; flappy_W(19, 452) <= 0; flappy_W(19, 453) <= 0; flappy_W(19, 454) <= 0; flappy_W(19, 455) <= 0; flappy_W(19, 456) <= 0; flappy_W(19, 457) <= 0; flappy_W(19, 458) <= 0; flappy_W(19, 459) <= 0; flappy_W(19, 460) <= 0; flappy_W(19, 461) <= 0; flappy_W(19, 462) <= 0; flappy_W(19, 463) <= 0; flappy_W(19, 464) <= 0; flappy_W(19, 465) <= 0; flappy_W(19, 466) <= 0; flappy_W(19, 467) <= 0; flappy_W(19, 468) <= 1; flappy_W(19, 469) <= 1; flappy_W(19, 470) <= 1; flappy_W(19, 471) <= 1; flappy_W(19, 472) <= 1; flappy_W(19, 473) <= 1; flappy_W(19, 474) <= 1; flappy_W(19, 475) <= 1; flappy_W(19, 476) <= 1; flappy_W(19, 477) <= 1; flappy_W(19, 478) <= 1; flappy_W(19, 479) <= 1; flappy_W(19, 480) <= 0; flappy_W(19, 481) <= 0; flappy_W(19, 482) <= 0; flappy_W(19, 483) <= 0; flappy_W(19, 484) <= 0; flappy_W(19, 485) <= 0; flappy_W(19, 486) <= 0; flappy_W(19, 487) <= 0; flappy_W(19, 488) <= 0; flappy_W(19, 489) <= 0; flappy_W(19, 490) <= 0; flappy_W(19, 491) <= 0; flappy_W(19, 492) <= 0; flappy_W(19, 493) <= 0; flappy_W(19, 494) <= 0; flappy_W(19, 495) <= 0; flappy_W(19, 496) <= 0; flappy_W(19, 497) <= 0; flappy_W(19, 498) <= 0; flappy_W(19, 499) <= 0; flappy_W(19, 500) <= 0; flappy_W(19, 501) <= 0; flappy_W(19, 502) <= 0; flappy_W(19, 503) <= 0; flappy_W(19, 504) <= 0; flappy_W(19, 505) <= 0; flappy_W(19, 506) <= 0; flappy_W(19, 507) <= 0; flappy_W(19, 508) <= 0; flappy_W(19, 509) <= 0; flappy_W(19, 510) <= 1; flappy_W(19, 511) <= 1; flappy_W(19, 512) <= 1; flappy_W(19, 513) <= 1; flappy_W(19, 514) <= 1; flappy_W(19, 515) <= 1; flappy_W(19, 516) <= 1; flappy_W(19, 517) <= 1; flappy_W(19, 518) <= 1; flappy_W(19, 519) <= 1; flappy_W(19, 520) <= 1; flappy_W(19, 521) <= 1; flappy_W(19, 522) <= 0; flappy_W(19, 523) <= 0; flappy_W(19, 524) <= 0; flappy_W(19, 525) <= 0; flappy_W(19, 526) <= 0; flappy_W(19, 527) <= 0; flappy_W(19, 528) <= 0; flappy_W(19, 529) <= 0; flappy_W(19, 530) <= 0; flappy_W(19, 531) <= 0; flappy_W(19, 532) <= 0; flappy_W(19, 533) <= 0; flappy_W(19, 534) <= 1; flappy_W(19, 535) <= 1; flappy_W(19, 536) <= 1; flappy_W(19, 537) <= 1; flappy_W(19, 538) <= 1; flappy_W(19, 539) <= 1; flappy_W(19, 540) <= 1; flappy_W(19, 541) <= 1; flappy_W(19, 542) <= 1; flappy_W(19, 543) <= 1; flappy_W(19, 544) <= 1; flappy_W(19, 545) <= 1; flappy_W(19, 546) <= 0; flappy_W(19, 547) <= 0; flappy_W(19, 548) <= 0; flappy_W(19, 549) <= 0; flappy_W(19, 550) <= 0; flappy_W(19, 551) <= 0; flappy_W(19, 552) <= 0; flappy_W(19, 553) <= 0; flappy_W(19, 554) <= 0; flappy_W(19, 555) <= 0; flappy_W(19, 556) <= 0; flappy_W(19, 557) <= 0; flappy_W(19, 558) <= 0; flappy_W(19, 559) <= 0; flappy_W(19, 560) <= 0; flappy_W(19, 561) <= 0; flappy_W(19, 562) <= 0; flappy_W(19, 563) <= 0; flappy_W(19, 564) <= 1; flappy_W(19, 565) <= 1; flappy_W(19, 566) <= 1; flappy_W(19, 567) <= 1; flappy_W(19, 568) <= 1; flappy_W(19, 569) <= 1; flappy_W(19, 570) <= 1; flappy_W(19, 571) <= 1; flappy_W(19, 572) <= 1; flappy_W(19, 573) <= 1; flappy_W(19, 574) <= 1; flappy_W(19, 575) <= 1; flappy_W(19, 576) <= 0; flappy_W(19, 577) <= 0; flappy_W(19, 578) <= 0; flappy_W(19, 579) <= 0; flappy_W(19, 580) <= 0; flappy_W(19, 581) <= 0; flappy_W(19, 582) <= 0; flappy_W(19, 583) <= 0; flappy_W(19, 584) <= 0; flappy_W(19, 585) <= 0; flappy_W(19, 586) <= 0; flappy_W(19, 587) <= 0; flappy_W(19, 588) <= 1; flappy_W(19, 589) <= 1; flappy_W(19, 590) <= 1; flappy_W(19, 591) <= 1; flappy_W(19, 592) <= 1; flappy_W(19, 593) <= 1; 
flappy_W(20, 0) <= 0; flappy_W(20, 1) <= 0; flappy_W(20, 2) <= 0; flappy_W(20, 3) <= 0; flappy_W(20, 4) <= 0; flappy_W(20, 5) <= 0; flappy_W(20, 6) <= 1; flappy_W(20, 7) <= 1; flappy_W(20, 8) <= 1; flappy_W(20, 9) <= 1; flappy_W(20, 10) <= 1; flappy_W(20, 11) <= 1; flappy_W(20, 12) <= 1; flappy_W(20, 13) <= 1; flappy_W(20, 14) <= 1; flappy_W(20, 15) <= 1; flappy_W(20, 16) <= 1; flappy_W(20, 17) <= 1; flappy_W(20, 18) <= 0; flappy_W(20, 19) <= 0; flappy_W(20, 20) <= 0; flappy_W(20, 21) <= 0; flappy_W(20, 22) <= 0; flappy_W(20, 23) <= 0; flappy_W(20, 24) <= 1; flappy_W(20, 25) <= 1; flappy_W(20, 26) <= 1; flappy_W(20, 27) <= 1; flappy_W(20, 28) <= 1; flappy_W(20, 29) <= 1; flappy_W(20, 30) <= 0; flappy_W(20, 31) <= 0; flappy_W(20, 32) <= 0; flappy_W(20, 33) <= 0; flappy_W(20, 34) <= 0; flappy_W(20, 35) <= 0; flappy_W(20, 36) <= 0; flappy_W(20, 37) <= 0; flappy_W(20, 38) <= 0; flappy_W(20, 39) <= 0; flappy_W(20, 40) <= 0; flappy_W(20, 41) <= 0; flappy_W(20, 42) <= 0; flappy_W(20, 43) <= 0; flappy_W(20, 44) <= 0; flappy_W(20, 45) <= 0; flappy_W(20, 46) <= 0; flappy_W(20, 47) <= 0; flappy_W(20, 48) <= 0; flappy_W(20, 49) <= 0; flappy_W(20, 50) <= 0; flappy_W(20, 51) <= 0; flappy_W(20, 52) <= 0; flappy_W(20, 53) <= 0; flappy_W(20, 54) <= 0; flappy_W(20, 55) <= 0; flappy_W(20, 56) <= 0; flappy_W(20, 57) <= 0; flappy_W(20, 58) <= 0; flappy_W(20, 59) <= 0; flappy_W(20, 60) <= 1; flappy_W(20, 61) <= 1; flappy_W(20, 62) <= 1; flappy_W(20, 63) <= 1; flappy_W(20, 64) <= 1; flappy_W(20, 65) <= 1; flappy_W(20, 66) <= 1; flappy_W(20, 67) <= 1; flappy_W(20, 68) <= 1; flappy_W(20, 69) <= 1; flappy_W(20, 70) <= 1; flappy_W(20, 71) <= 1; flappy_W(20, 72) <= 0; flappy_W(20, 73) <= 0; flappy_W(20, 74) <= 0; flappy_W(20, 75) <= 0; flappy_W(20, 76) <= 0; flappy_W(20, 77) <= 0; flappy_W(20, 78) <= 0; flappy_W(20, 79) <= 0; flappy_W(20, 80) <= 0; flappy_W(20, 81) <= 0; flappy_W(20, 82) <= 0; flappy_W(20, 83) <= 0; flappy_W(20, 84) <= 0; flappy_W(20, 85) <= 0; flappy_W(20, 86) <= 0; flappy_W(20, 87) <= 0; flappy_W(20, 88) <= 0; flappy_W(20, 89) <= 0; flappy_W(20, 90) <= 0; flappy_W(20, 91) <= 0; flappy_W(20, 92) <= 0; flappy_W(20, 93) <= 0; flappy_W(20, 94) <= 0; flappy_W(20, 95) <= 0; flappy_W(20, 96) <= 0; flappy_W(20, 97) <= 0; flappy_W(20, 98) <= 0; flappy_W(20, 99) <= 0; flappy_W(20, 100) <= 0; flappy_W(20, 101) <= 0; flappy_W(20, 102) <= 0; flappy_W(20, 103) <= 0; flappy_W(20, 104) <= 0; flappy_W(20, 105) <= 0; flappy_W(20, 106) <= 0; flappy_W(20, 107) <= 0; flappy_W(20, 108) <= 1; flappy_W(20, 109) <= 1; flappy_W(20, 110) <= 1; flappy_W(20, 111) <= 1; flappy_W(20, 112) <= 1; flappy_W(20, 113) <= 1; flappy_W(20, 114) <= 1; flappy_W(20, 115) <= 1; flappy_W(20, 116) <= 1; flappy_W(20, 117) <= 1; flappy_W(20, 118) <= 1; flappy_W(20, 119) <= 1; flappy_W(20, 120) <= 0; flappy_W(20, 121) <= 0; flappy_W(20, 122) <= 0; flappy_W(20, 123) <= 0; flappy_W(20, 124) <= 0; flappy_W(20, 125) <= 0; flappy_W(20, 126) <= 0; flappy_W(20, 127) <= 0; flappy_W(20, 128) <= 0; flappy_W(20, 129) <= 0; flappy_W(20, 130) <= 0; flappy_W(20, 131) <= 0; flappy_W(20, 132) <= 0; flappy_W(20, 133) <= 0; flappy_W(20, 134) <= 0; flappy_W(20, 135) <= 0; flappy_W(20, 136) <= 0; flappy_W(20, 137) <= 0; flappy_W(20, 138) <= 1; flappy_W(20, 139) <= 1; flappy_W(20, 140) <= 1; flappy_W(20, 141) <= 1; flappy_W(20, 142) <= 1; flappy_W(20, 143) <= 1; flappy_W(20, 144) <= 1; flappy_W(20, 145) <= 1; flappy_W(20, 146) <= 1; flappy_W(20, 147) <= 1; flappy_W(20, 148) <= 1; flappy_W(20, 149) <= 1; flappy_W(20, 150) <= 0; flappy_W(20, 151) <= 0; flappy_W(20, 152) <= 0; flappy_W(20, 153) <= 0; flappy_W(20, 154) <= 0; flappy_W(20, 155) <= 0; flappy_W(20, 156) <= 0; flappy_W(20, 157) <= 0; flappy_W(20, 158) <= 0; flappy_W(20, 159) <= 0; flappy_W(20, 160) <= 0; flappy_W(20, 161) <= 0; flappy_W(20, 162) <= 0; flappy_W(20, 163) <= 0; flappy_W(20, 164) <= 0; flappy_W(20, 165) <= 0; flappy_W(20, 166) <= 0; flappy_W(20, 167) <= 0; flappy_W(20, 168) <= 1; flappy_W(20, 169) <= 1; flappy_W(20, 170) <= 1; flappy_W(20, 171) <= 1; flappy_W(20, 172) <= 1; flappy_W(20, 173) <= 1; flappy_W(20, 174) <= 1; flappy_W(20, 175) <= 1; flappy_W(20, 176) <= 1; flappy_W(20, 177) <= 1; flappy_W(20, 178) <= 1; flappy_W(20, 179) <= 1; flappy_W(20, 180) <= 0; flappy_W(20, 181) <= 0; flappy_W(20, 182) <= 0; flappy_W(20, 183) <= 0; flappy_W(20, 184) <= 0; flappy_W(20, 185) <= 0; flappy_W(20, 186) <= 0; flappy_W(20, 187) <= 0; flappy_W(20, 188) <= 0; flappy_W(20, 189) <= 0; flappy_W(20, 190) <= 0; flappy_W(20, 191) <= 0; flappy_W(20, 192) <= 1; flappy_W(20, 193) <= 1; flappy_W(20, 194) <= 1; flappy_W(20, 195) <= 1; flappy_W(20, 196) <= 1; flappy_W(20, 197) <= 1; flappy_W(20, 198) <= 1; flappy_W(20, 199) <= 1; flappy_W(20, 200) <= 1; flappy_W(20, 201) <= 1; flappy_W(20, 202) <= 1; flappy_W(20, 203) <= 1; flappy_W(20, 204) <= 0; flappy_W(20, 205) <= 0; flappy_W(20, 206) <= 0; flappy_W(20, 207) <= 0; flappy_W(20, 208) <= 0; flappy_W(20, 209) <= 0; flappy_W(20, 210) <= 0; flappy_W(20, 211) <= 0; flappy_W(20, 212) <= 0; flappy_W(20, 213) <= 0; flappy_W(20, 214) <= 0; flappy_W(20, 215) <= 0; flappy_W(20, 216) <= 0; flappy_W(20, 217) <= 0; flappy_W(20, 218) <= 0; flappy_W(20, 219) <= 0; flappy_W(20, 220) <= 0; flappy_W(20, 221) <= 0; flappy_W(20, 222) <= 1; flappy_W(20, 223) <= 1; flappy_W(20, 224) <= 1; flappy_W(20, 225) <= 1; flappy_W(20, 226) <= 1; flappy_W(20, 227) <= 1; flappy_W(20, 228) <= 1; flappy_W(20, 229) <= 1; flappy_W(20, 230) <= 1; flappy_W(20, 231) <= 1; flappy_W(20, 232) <= 1; flappy_W(20, 233) <= 1; flappy_W(20, 234) <= 0; flappy_W(20, 235) <= 0; flappy_W(20, 236) <= 0; flappy_W(20, 237) <= 0; flappy_W(20, 238) <= 0; flappy_W(20, 239) <= 0; flappy_W(20, 240) <= 0; flappy_W(20, 241) <= 0; flappy_W(20, 242) <= 0; flappy_W(20, 243) <= 0; flappy_W(20, 244) <= 0; flappy_W(20, 245) <= 0; flappy_W(20, 246) <= 1; flappy_W(20, 247) <= 1; flappy_W(20, 248) <= 1; flappy_W(20, 249) <= 1; flappy_W(20, 250) <= 1; flappy_W(20, 251) <= 1; flappy_W(20, 252) <= 1; flappy_W(20, 253) <= 1; flappy_W(20, 254) <= 1; flappy_W(20, 255) <= 1; flappy_W(20, 256) <= 1; flappy_W(20, 257) <= 1; flappy_W(20, 258) <= 0; flappy_W(20, 259) <= 0; flappy_W(20, 260) <= 0; flappy_W(20, 261) <= 0; flappy_W(20, 262) <= 0; flappy_W(20, 263) <= 0; flappy_W(20, 264) <= 0; flappy_W(20, 265) <= 0; flappy_W(20, 266) <= 0; flappy_W(20, 267) <= 0; flappy_W(20, 268) <= 0; flappy_W(20, 269) <= 0; flappy_W(20, 270) <= 0; flappy_W(20, 271) <= 0; flappy_W(20, 272) <= 0; flappy_W(20, 273) <= 0; flappy_W(20, 274) <= 0; flappy_W(20, 275) <= 0; flappy_W(20, 276) <= 1; flappy_W(20, 277) <= 1; flappy_W(20, 278) <= 1; flappy_W(20, 279) <= 1; flappy_W(20, 280) <= 1; flappy_W(20, 281) <= 1; flappy_W(20, 282) <= 1; flappy_W(20, 283) <= 1; flappy_W(20, 284) <= 1; flappy_W(20, 285) <= 1; flappy_W(20, 286) <= 1; flappy_W(20, 287) <= 1; flappy_W(20, 288) <= 0; flappy_W(20, 289) <= 0; flappy_W(20, 290) <= 0; flappy_W(20, 291) <= 0; flappy_W(20, 292) <= 0; flappy_W(20, 293) <= 0; flappy_W(20, 294) <= 0; flappy_W(20, 295) <= 0; flappy_W(20, 296) <= 0; flappy_W(20, 297) <= 0; flappy_W(20, 298) <= 0; flappy_W(20, 299) <= 0; flappy_W(20, 300) <= 1; flappy_W(20, 301) <= 1; flappy_W(20, 302) <= 1; flappy_W(20, 303) <= 1; flappy_W(20, 304) <= 1; flappy_W(20, 305) <= 1; flappy_W(20, 306) <= 1; flappy_W(20, 307) <= 1; flappy_W(20, 308) <= 1; flappy_W(20, 309) <= 1; flappy_W(20, 310) <= 1; flappy_W(20, 311) <= 1; flappy_W(20, 312) <= 0; flappy_W(20, 313) <= 0; flappy_W(20, 314) <= 0; flappy_W(20, 315) <= 0; flappy_W(20, 316) <= 0; flappy_W(20, 317) <= 0; flappy_W(20, 318) <= 0; flappy_W(20, 319) <= 0; flappy_W(20, 320) <= 0; flappy_W(20, 321) <= 0; flappy_W(20, 322) <= 0; flappy_W(20, 323) <= 0; flappy_W(20, 324) <= 0; flappy_W(20, 325) <= 0; flappy_W(20, 326) <= 0; flappy_W(20, 327) <= 0; flappy_W(20, 328) <= 0; flappy_W(20, 329) <= 0; flappy_W(20, 330) <= 0; flappy_W(20, 331) <= 0; flappy_W(20, 332) <= 0; flappy_W(20, 333) <= 0; flappy_W(20, 334) <= 0; flappy_W(20, 335) <= 0; flappy_W(20, 336) <= 0; flappy_W(20, 337) <= 0; flappy_W(20, 338) <= 0; flappy_W(20, 339) <= 0; flappy_W(20, 340) <= 0; flappy_W(20, 341) <= 0; flappy_W(20, 342) <= 0; flappy_W(20, 343) <= 0; flappy_W(20, 344) <= 0; flappy_W(20, 345) <= 0; flappy_W(20, 346) <= 0; flappy_W(20, 347) <= 0; flappy_W(20, 348) <= 0; flappy_W(20, 349) <= 0; flappy_W(20, 350) <= 0; flappy_W(20, 351) <= 0; flappy_W(20, 352) <= 0; flappy_W(20, 353) <= 0; flappy_W(20, 354) <= 0; flappy_W(20, 355) <= 0; flappy_W(20, 356) <= 0; flappy_W(20, 357) <= 0; flappy_W(20, 358) <= 0; flappy_W(20, 359) <= 0; flappy_W(20, 360) <= 0; flappy_W(20, 361) <= 0; flappy_W(20, 362) <= 0; flappy_W(20, 363) <= 0; flappy_W(20, 364) <= 0; flappy_W(20, 365) <= 0; flappy_W(20, 366) <= 0; flappy_W(20, 367) <= 0; flappy_W(20, 368) <= 0; flappy_W(20, 369) <= 0; flappy_W(20, 370) <= 0; flappy_W(20, 371) <= 0; flappy_W(20, 372) <= 0; flappy_W(20, 373) <= 0; flappy_W(20, 374) <= 0; flappy_W(20, 375) <= 0; flappy_W(20, 376) <= 0; flappy_W(20, 377) <= 0; flappy_W(20, 378) <= 0; flappy_W(20, 379) <= 0; flappy_W(20, 380) <= 0; flappy_W(20, 381) <= 0; flappy_W(20, 382) <= 0; flappy_W(20, 383) <= 0; flappy_W(20, 384) <= 0; flappy_W(20, 385) <= 0; flappy_W(20, 386) <= 0; flappy_W(20, 387) <= 0; flappy_W(20, 388) <= 0; flappy_W(20, 389) <= 0; flappy_W(20, 390) <= 0; flappy_W(20, 391) <= 0; flappy_W(20, 392) <= 0; flappy_W(20, 393) <= 0; flappy_W(20, 394) <= 0; flappy_W(20, 395) <= 0; flappy_W(20, 396) <= 0; flappy_W(20, 397) <= 0; flappy_W(20, 398) <= 0; flappy_W(20, 399) <= 0; flappy_W(20, 400) <= 0; flappy_W(20, 401) <= 0; flappy_W(20, 402) <= 1; flappy_W(20, 403) <= 1; flappy_W(20, 404) <= 1; flappy_W(20, 405) <= 1; flappy_W(20, 406) <= 1; flappy_W(20, 407) <= 1; flappy_W(20, 408) <= 1; flappy_W(20, 409) <= 1; flappy_W(20, 410) <= 1; flappy_W(20, 411) <= 1; flappy_W(20, 412) <= 1; flappy_W(20, 413) <= 1; flappy_W(20, 414) <= 0; flappy_W(20, 415) <= 0; flappy_W(20, 416) <= 0; flappy_W(20, 417) <= 0; flappy_W(20, 418) <= 0; flappy_W(20, 419) <= 0; flappy_W(20, 420) <= 0; flappy_W(20, 421) <= 0; flappy_W(20, 422) <= 0; flappy_W(20, 423) <= 0; flappy_W(20, 424) <= 0; flappy_W(20, 425) <= 0; flappy_W(20, 426) <= 1; flappy_W(20, 427) <= 1; flappy_W(20, 428) <= 1; flappy_W(20, 429) <= 1; flappy_W(20, 430) <= 1; flappy_W(20, 431) <= 1; flappy_W(20, 432) <= 1; flappy_W(20, 433) <= 1; flappy_W(20, 434) <= 1; flappy_W(20, 435) <= 1; flappy_W(20, 436) <= 1; flappy_W(20, 437) <= 1; flappy_W(20, 438) <= 0; flappy_W(20, 439) <= 0; flappy_W(20, 440) <= 0; flappy_W(20, 441) <= 0; flappy_W(20, 442) <= 0; flappy_W(20, 443) <= 0; flappy_W(20, 444) <= 0; flappy_W(20, 445) <= 0; flappy_W(20, 446) <= 0; flappy_W(20, 447) <= 0; flappy_W(20, 448) <= 0; flappy_W(20, 449) <= 0; flappy_W(20, 450) <= 0; flappy_W(20, 451) <= 0; flappy_W(20, 452) <= 0; flappy_W(20, 453) <= 0; flappy_W(20, 454) <= 0; flappy_W(20, 455) <= 0; flappy_W(20, 456) <= 0; flappy_W(20, 457) <= 0; flappy_W(20, 458) <= 0; flappy_W(20, 459) <= 0; flappy_W(20, 460) <= 0; flappy_W(20, 461) <= 0; flappy_W(20, 462) <= 0; flappy_W(20, 463) <= 0; flappy_W(20, 464) <= 0; flappy_W(20, 465) <= 0; flappy_W(20, 466) <= 0; flappy_W(20, 467) <= 0; flappy_W(20, 468) <= 1; flappy_W(20, 469) <= 1; flappy_W(20, 470) <= 1; flappy_W(20, 471) <= 1; flappy_W(20, 472) <= 1; flappy_W(20, 473) <= 1; flappy_W(20, 474) <= 1; flappy_W(20, 475) <= 1; flappy_W(20, 476) <= 1; flappy_W(20, 477) <= 1; flappy_W(20, 478) <= 1; flappy_W(20, 479) <= 1; flappy_W(20, 480) <= 0; flappy_W(20, 481) <= 0; flappy_W(20, 482) <= 0; flappy_W(20, 483) <= 0; flappy_W(20, 484) <= 0; flappy_W(20, 485) <= 0; flappy_W(20, 486) <= 0; flappy_W(20, 487) <= 0; flappy_W(20, 488) <= 0; flappy_W(20, 489) <= 0; flappy_W(20, 490) <= 0; flappy_W(20, 491) <= 0; flappy_W(20, 492) <= 0; flappy_W(20, 493) <= 0; flappy_W(20, 494) <= 0; flappy_W(20, 495) <= 0; flappy_W(20, 496) <= 0; flappy_W(20, 497) <= 0; flappy_W(20, 498) <= 0; flappy_W(20, 499) <= 0; flappy_W(20, 500) <= 0; flappy_W(20, 501) <= 0; flappy_W(20, 502) <= 0; flappy_W(20, 503) <= 0; flappy_W(20, 504) <= 0; flappy_W(20, 505) <= 0; flappy_W(20, 506) <= 0; flappy_W(20, 507) <= 0; flappy_W(20, 508) <= 0; flappy_W(20, 509) <= 0; flappy_W(20, 510) <= 1; flappy_W(20, 511) <= 1; flappy_W(20, 512) <= 1; flappy_W(20, 513) <= 1; flappy_W(20, 514) <= 1; flappy_W(20, 515) <= 1; flappy_W(20, 516) <= 1; flappy_W(20, 517) <= 1; flappy_W(20, 518) <= 1; flappy_W(20, 519) <= 1; flappy_W(20, 520) <= 1; flappy_W(20, 521) <= 1; flappy_W(20, 522) <= 0; flappy_W(20, 523) <= 0; flappy_W(20, 524) <= 0; flappy_W(20, 525) <= 0; flappy_W(20, 526) <= 0; flappy_W(20, 527) <= 0; flappy_W(20, 528) <= 0; flappy_W(20, 529) <= 0; flappy_W(20, 530) <= 0; flappy_W(20, 531) <= 0; flappy_W(20, 532) <= 0; flappy_W(20, 533) <= 0; flappy_W(20, 534) <= 1; flappy_W(20, 535) <= 1; flappy_W(20, 536) <= 1; flappy_W(20, 537) <= 1; flappy_W(20, 538) <= 1; flappy_W(20, 539) <= 1; flappy_W(20, 540) <= 1; flappy_W(20, 541) <= 1; flappy_W(20, 542) <= 1; flappy_W(20, 543) <= 1; flappy_W(20, 544) <= 1; flappy_W(20, 545) <= 1; flappy_W(20, 546) <= 0; flappy_W(20, 547) <= 0; flappy_W(20, 548) <= 0; flappy_W(20, 549) <= 0; flappy_W(20, 550) <= 0; flappy_W(20, 551) <= 0; flappy_W(20, 552) <= 0; flappy_W(20, 553) <= 0; flappy_W(20, 554) <= 0; flappy_W(20, 555) <= 0; flappy_W(20, 556) <= 0; flappy_W(20, 557) <= 0; flappy_W(20, 558) <= 0; flappy_W(20, 559) <= 0; flappy_W(20, 560) <= 0; flappy_W(20, 561) <= 0; flappy_W(20, 562) <= 0; flappy_W(20, 563) <= 0; flappy_W(20, 564) <= 1; flappy_W(20, 565) <= 1; flappy_W(20, 566) <= 1; flappy_W(20, 567) <= 1; flappy_W(20, 568) <= 1; flappy_W(20, 569) <= 1; flappy_W(20, 570) <= 1; flappy_W(20, 571) <= 1; flappy_W(20, 572) <= 1; flappy_W(20, 573) <= 1; flappy_W(20, 574) <= 1; flappy_W(20, 575) <= 1; flappy_W(20, 576) <= 0; flappy_W(20, 577) <= 0; flappy_W(20, 578) <= 0; flappy_W(20, 579) <= 0; flappy_W(20, 580) <= 0; flappy_W(20, 581) <= 0; flappy_W(20, 582) <= 0; flappy_W(20, 583) <= 0; flappy_W(20, 584) <= 0; flappy_W(20, 585) <= 0; flappy_W(20, 586) <= 0; flappy_W(20, 587) <= 0; flappy_W(20, 588) <= 1; flappy_W(20, 589) <= 1; flappy_W(20, 590) <= 1; flappy_W(20, 591) <= 1; flappy_W(20, 592) <= 1; flappy_W(20, 593) <= 1; 
flappy_W(21, 0) <= 0; flappy_W(21, 1) <= 0; flappy_W(21, 2) <= 0; flappy_W(21, 3) <= 0; flappy_W(21, 4) <= 0; flappy_W(21, 5) <= 0; flappy_W(21, 6) <= 1; flappy_W(21, 7) <= 1; flappy_W(21, 8) <= 1; flappy_W(21, 9) <= 1; flappy_W(21, 10) <= 1; flappy_W(21, 11) <= 1; flappy_W(21, 12) <= 1; flappy_W(21, 13) <= 1; flappy_W(21, 14) <= 1; flappy_W(21, 15) <= 1; flappy_W(21, 16) <= 1; flappy_W(21, 17) <= 1; flappy_W(21, 18) <= 0; flappy_W(21, 19) <= 0; flappy_W(21, 20) <= 0; flappy_W(21, 21) <= 0; flappy_W(21, 22) <= 0; flappy_W(21, 23) <= 0; flappy_W(21, 24) <= 1; flappy_W(21, 25) <= 1; flappy_W(21, 26) <= 1; flappy_W(21, 27) <= 1; flappy_W(21, 28) <= 1; flappy_W(21, 29) <= 1; flappy_W(21, 30) <= 0; flappy_W(21, 31) <= 0; flappy_W(21, 32) <= 0; flappy_W(21, 33) <= 0; flappy_W(21, 34) <= 0; flappy_W(21, 35) <= 0; flappy_W(21, 36) <= 0; flappy_W(21, 37) <= 0; flappy_W(21, 38) <= 0; flappy_W(21, 39) <= 0; flappy_W(21, 40) <= 0; flappy_W(21, 41) <= 0; flappy_W(21, 42) <= 0; flappy_W(21, 43) <= 0; flappy_W(21, 44) <= 0; flappy_W(21, 45) <= 0; flappy_W(21, 46) <= 0; flappy_W(21, 47) <= 0; flappy_W(21, 48) <= 0; flappy_W(21, 49) <= 0; flappy_W(21, 50) <= 0; flappy_W(21, 51) <= 0; flappy_W(21, 52) <= 0; flappy_W(21, 53) <= 0; flappy_W(21, 54) <= 0; flappy_W(21, 55) <= 0; flappy_W(21, 56) <= 0; flappy_W(21, 57) <= 0; flappy_W(21, 58) <= 0; flappy_W(21, 59) <= 0; flappy_W(21, 60) <= 1; flappy_W(21, 61) <= 1; flappy_W(21, 62) <= 1; flappy_W(21, 63) <= 1; flappy_W(21, 64) <= 1; flappy_W(21, 65) <= 1; flappy_W(21, 66) <= 1; flappy_W(21, 67) <= 1; flappy_W(21, 68) <= 1; flappy_W(21, 69) <= 1; flappy_W(21, 70) <= 1; flappy_W(21, 71) <= 1; flappy_W(21, 72) <= 0; flappy_W(21, 73) <= 0; flappy_W(21, 74) <= 0; flappy_W(21, 75) <= 0; flappy_W(21, 76) <= 0; flappy_W(21, 77) <= 0; flappy_W(21, 78) <= 0; flappy_W(21, 79) <= 0; flappy_W(21, 80) <= 0; flappy_W(21, 81) <= 0; flappy_W(21, 82) <= 0; flappy_W(21, 83) <= 0; flappy_W(21, 84) <= 0; flappy_W(21, 85) <= 0; flappy_W(21, 86) <= 0; flappy_W(21, 87) <= 0; flappy_W(21, 88) <= 0; flappy_W(21, 89) <= 0; flappy_W(21, 90) <= 0; flappy_W(21, 91) <= 0; flappy_W(21, 92) <= 0; flappy_W(21, 93) <= 0; flappy_W(21, 94) <= 0; flappy_W(21, 95) <= 0; flappy_W(21, 96) <= 0; flappy_W(21, 97) <= 0; flappy_W(21, 98) <= 0; flappy_W(21, 99) <= 0; flappy_W(21, 100) <= 0; flappy_W(21, 101) <= 0; flappy_W(21, 102) <= 0; flappy_W(21, 103) <= 0; flappy_W(21, 104) <= 0; flappy_W(21, 105) <= 0; flappy_W(21, 106) <= 0; flappy_W(21, 107) <= 0; flappy_W(21, 108) <= 1; flappy_W(21, 109) <= 1; flappy_W(21, 110) <= 1; flappy_W(21, 111) <= 1; flappy_W(21, 112) <= 1; flappy_W(21, 113) <= 1; flappy_W(21, 114) <= 1; flappy_W(21, 115) <= 1; flappy_W(21, 116) <= 1; flappy_W(21, 117) <= 1; flappy_W(21, 118) <= 1; flappy_W(21, 119) <= 1; flappy_W(21, 120) <= 0; flappy_W(21, 121) <= 0; flappy_W(21, 122) <= 0; flappy_W(21, 123) <= 0; flappy_W(21, 124) <= 0; flappy_W(21, 125) <= 0; flappy_W(21, 126) <= 0; flappy_W(21, 127) <= 0; flappy_W(21, 128) <= 0; flappy_W(21, 129) <= 0; flappy_W(21, 130) <= 0; flappy_W(21, 131) <= 0; flappy_W(21, 132) <= 0; flappy_W(21, 133) <= 0; flappy_W(21, 134) <= 0; flappy_W(21, 135) <= 0; flappy_W(21, 136) <= 0; flappy_W(21, 137) <= 0; flappy_W(21, 138) <= 1; flappy_W(21, 139) <= 1; flappy_W(21, 140) <= 1; flappy_W(21, 141) <= 1; flappy_W(21, 142) <= 1; flappy_W(21, 143) <= 1; flappy_W(21, 144) <= 1; flappy_W(21, 145) <= 1; flappy_W(21, 146) <= 1; flappy_W(21, 147) <= 1; flappy_W(21, 148) <= 1; flappy_W(21, 149) <= 1; flappy_W(21, 150) <= 0; flappy_W(21, 151) <= 0; flappy_W(21, 152) <= 0; flappy_W(21, 153) <= 0; flappy_W(21, 154) <= 0; flappy_W(21, 155) <= 0; flappy_W(21, 156) <= 0; flappy_W(21, 157) <= 0; flappy_W(21, 158) <= 0; flappy_W(21, 159) <= 0; flappy_W(21, 160) <= 0; flappy_W(21, 161) <= 0; flappy_W(21, 162) <= 0; flappy_W(21, 163) <= 0; flappy_W(21, 164) <= 0; flappy_W(21, 165) <= 0; flappy_W(21, 166) <= 0; flappy_W(21, 167) <= 0; flappy_W(21, 168) <= 1; flappy_W(21, 169) <= 1; flappy_W(21, 170) <= 1; flappy_W(21, 171) <= 1; flappy_W(21, 172) <= 1; flappy_W(21, 173) <= 1; flappy_W(21, 174) <= 1; flappy_W(21, 175) <= 1; flappy_W(21, 176) <= 1; flappy_W(21, 177) <= 1; flappy_W(21, 178) <= 1; flappy_W(21, 179) <= 1; flappy_W(21, 180) <= 0; flappy_W(21, 181) <= 0; flappy_W(21, 182) <= 0; flappy_W(21, 183) <= 0; flappy_W(21, 184) <= 0; flappy_W(21, 185) <= 0; flappy_W(21, 186) <= 0; flappy_W(21, 187) <= 0; flappy_W(21, 188) <= 0; flappy_W(21, 189) <= 0; flappy_W(21, 190) <= 0; flappy_W(21, 191) <= 0; flappy_W(21, 192) <= 1; flappy_W(21, 193) <= 1; flappy_W(21, 194) <= 1; flappy_W(21, 195) <= 1; flappy_W(21, 196) <= 1; flappy_W(21, 197) <= 1; flappy_W(21, 198) <= 1; flappy_W(21, 199) <= 1; flappy_W(21, 200) <= 1; flappy_W(21, 201) <= 1; flappy_W(21, 202) <= 1; flappy_W(21, 203) <= 1; flappy_W(21, 204) <= 0; flappy_W(21, 205) <= 0; flappy_W(21, 206) <= 0; flappy_W(21, 207) <= 0; flappy_W(21, 208) <= 0; flappy_W(21, 209) <= 0; flappy_W(21, 210) <= 0; flappy_W(21, 211) <= 0; flappy_W(21, 212) <= 0; flappy_W(21, 213) <= 0; flappy_W(21, 214) <= 0; flappy_W(21, 215) <= 0; flappy_W(21, 216) <= 0; flappy_W(21, 217) <= 0; flappy_W(21, 218) <= 0; flappy_W(21, 219) <= 0; flappy_W(21, 220) <= 0; flappy_W(21, 221) <= 0; flappy_W(21, 222) <= 1; flappy_W(21, 223) <= 1; flappy_W(21, 224) <= 1; flappy_W(21, 225) <= 1; flappy_W(21, 226) <= 1; flappy_W(21, 227) <= 1; flappy_W(21, 228) <= 1; flappy_W(21, 229) <= 1; flappy_W(21, 230) <= 1; flappy_W(21, 231) <= 1; flappy_W(21, 232) <= 1; flappy_W(21, 233) <= 1; flappy_W(21, 234) <= 0; flappy_W(21, 235) <= 0; flappy_W(21, 236) <= 0; flappy_W(21, 237) <= 0; flappy_W(21, 238) <= 0; flappy_W(21, 239) <= 0; flappy_W(21, 240) <= 0; flappy_W(21, 241) <= 0; flappy_W(21, 242) <= 0; flappy_W(21, 243) <= 0; flappy_W(21, 244) <= 0; flappy_W(21, 245) <= 0; flappy_W(21, 246) <= 1; flappy_W(21, 247) <= 1; flappy_W(21, 248) <= 1; flappy_W(21, 249) <= 1; flappy_W(21, 250) <= 1; flappy_W(21, 251) <= 1; flappy_W(21, 252) <= 1; flappy_W(21, 253) <= 1; flappy_W(21, 254) <= 1; flappy_W(21, 255) <= 1; flappy_W(21, 256) <= 1; flappy_W(21, 257) <= 1; flappy_W(21, 258) <= 0; flappy_W(21, 259) <= 0; flappy_W(21, 260) <= 0; flappy_W(21, 261) <= 0; flappy_W(21, 262) <= 0; flappy_W(21, 263) <= 0; flappy_W(21, 264) <= 0; flappy_W(21, 265) <= 0; flappy_W(21, 266) <= 0; flappy_W(21, 267) <= 0; flappy_W(21, 268) <= 0; flappy_W(21, 269) <= 0; flappy_W(21, 270) <= 0; flappy_W(21, 271) <= 0; flappy_W(21, 272) <= 0; flappy_W(21, 273) <= 0; flappy_W(21, 274) <= 0; flappy_W(21, 275) <= 0; flappy_W(21, 276) <= 1; flappy_W(21, 277) <= 1; flappy_W(21, 278) <= 1; flappy_W(21, 279) <= 1; flappy_W(21, 280) <= 1; flappy_W(21, 281) <= 1; flappy_W(21, 282) <= 1; flappy_W(21, 283) <= 1; flappy_W(21, 284) <= 1; flappy_W(21, 285) <= 1; flappy_W(21, 286) <= 1; flappy_W(21, 287) <= 1; flappy_W(21, 288) <= 0; flappy_W(21, 289) <= 0; flappy_W(21, 290) <= 0; flappy_W(21, 291) <= 0; flappy_W(21, 292) <= 0; flappy_W(21, 293) <= 0; flappy_W(21, 294) <= 0; flappy_W(21, 295) <= 0; flappy_W(21, 296) <= 0; flappy_W(21, 297) <= 0; flappy_W(21, 298) <= 0; flappy_W(21, 299) <= 0; flappy_W(21, 300) <= 1; flappy_W(21, 301) <= 1; flappy_W(21, 302) <= 1; flappy_W(21, 303) <= 1; flappy_W(21, 304) <= 1; flappy_W(21, 305) <= 1; flappy_W(21, 306) <= 1; flappy_W(21, 307) <= 1; flappy_W(21, 308) <= 1; flappy_W(21, 309) <= 1; flappy_W(21, 310) <= 1; flappy_W(21, 311) <= 1; flappy_W(21, 312) <= 0; flappy_W(21, 313) <= 0; flappy_W(21, 314) <= 0; flappy_W(21, 315) <= 0; flappy_W(21, 316) <= 0; flappy_W(21, 317) <= 0; flappy_W(21, 318) <= 0; flappy_W(21, 319) <= 0; flappy_W(21, 320) <= 0; flappy_W(21, 321) <= 0; flappy_W(21, 322) <= 0; flappy_W(21, 323) <= 0; flappy_W(21, 324) <= 0; flappy_W(21, 325) <= 0; flappy_W(21, 326) <= 0; flappy_W(21, 327) <= 0; flappy_W(21, 328) <= 0; flappy_W(21, 329) <= 0; flappy_W(21, 330) <= 0; flappy_W(21, 331) <= 0; flappy_W(21, 332) <= 0; flappy_W(21, 333) <= 0; flappy_W(21, 334) <= 0; flappy_W(21, 335) <= 0; flappy_W(21, 336) <= 0; flappy_W(21, 337) <= 0; flappy_W(21, 338) <= 0; flappy_W(21, 339) <= 0; flappy_W(21, 340) <= 0; flappy_W(21, 341) <= 0; flappy_W(21, 342) <= 0; flappy_W(21, 343) <= 0; flappy_W(21, 344) <= 0; flappy_W(21, 345) <= 0; flappy_W(21, 346) <= 0; flappy_W(21, 347) <= 0; flappy_W(21, 348) <= 0; flappy_W(21, 349) <= 0; flappy_W(21, 350) <= 0; flappy_W(21, 351) <= 0; flappy_W(21, 352) <= 0; flappy_W(21, 353) <= 0; flappy_W(21, 354) <= 0; flappy_W(21, 355) <= 0; flappy_W(21, 356) <= 0; flappy_W(21, 357) <= 0; flappy_W(21, 358) <= 0; flappy_W(21, 359) <= 0; flappy_W(21, 360) <= 0; flappy_W(21, 361) <= 0; flappy_W(21, 362) <= 0; flappy_W(21, 363) <= 0; flappy_W(21, 364) <= 0; flappy_W(21, 365) <= 0; flappy_W(21, 366) <= 0; flappy_W(21, 367) <= 0; flappy_W(21, 368) <= 0; flappy_W(21, 369) <= 0; flappy_W(21, 370) <= 0; flappy_W(21, 371) <= 0; flappy_W(21, 372) <= 0; flappy_W(21, 373) <= 0; flappy_W(21, 374) <= 0; flappy_W(21, 375) <= 0; flappy_W(21, 376) <= 0; flappy_W(21, 377) <= 0; flappy_W(21, 378) <= 0; flappy_W(21, 379) <= 0; flappy_W(21, 380) <= 0; flappy_W(21, 381) <= 0; flappy_W(21, 382) <= 0; flappy_W(21, 383) <= 0; flappy_W(21, 384) <= 0; flappy_W(21, 385) <= 0; flappy_W(21, 386) <= 0; flappy_W(21, 387) <= 0; flappy_W(21, 388) <= 0; flappy_W(21, 389) <= 0; flappy_W(21, 390) <= 0; flappy_W(21, 391) <= 0; flappy_W(21, 392) <= 0; flappy_W(21, 393) <= 0; flappy_W(21, 394) <= 0; flappy_W(21, 395) <= 0; flappy_W(21, 396) <= 0; flappy_W(21, 397) <= 0; flappy_W(21, 398) <= 0; flappy_W(21, 399) <= 0; flappy_W(21, 400) <= 0; flappy_W(21, 401) <= 0; flappy_W(21, 402) <= 1; flappy_W(21, 403) <= 1; flappy_W(21, 404) <= 1; flappy_W(21, 405) <= 1; flappy_W(21, 406) <= 1; flappy_W(21, 407) <= 1; flappy_W(21, 408) <= 1; flappy_W(21, 409) <= 1; flappy_W(21, 410) <= 1; flappy_W(21, 411) <= 1; flappy_W(21, 412) <= 1; flappy_W(21, 413) <= 1; flappy_W(21, 414) <= 0; flappy_W(21, 415) <= 0; flappy_W(21, 416) <= 0; flappy_W(21, 417) <= 0; flappy_W(21, 418) <= 0; flappy_W(21, 419) <= 0; flappy_W(21, 420) <= 0; flappy_W(21, 421) <= 0; flappy_W(21, 422) <= 0; flappy_W(21, 423) <= 0; flappy_W(21, 424) <= 0; flappy_W(21, 425) <= 0; flappy_W(21, 426) <= 1; flappy_W(21, 427) <= 1; flappy_W(21, 428) <= 1; flappy_W(21, 429) <= 1; flappy_W(21, 430) <= 1; flappy_W(21, 431) <= 1; flappy_W(21, 432) <= 1; flappy_W(21, 433) <= 1; flappy_W(21, 434) <= 1; flappy_W(21, 435) <= 1; flappy_W(21, 436) <= 1; flappy_W(21, 437) <= 1; flappy_W(21, 438) <= 0; flappy_W(21, 439) <= 0; flappy_W(21, 440) <= 0; flappy_W(21, 441) <= 0; flappy_W(21, 442) <= 0; flappy_W(21, 443) <= 0; flappy_W(21, 444) <= 0; flappy_W(21, 445) <= 0; flappy_W(21, 446) <= 0; flappy_W(21, 447) <= 0; flappy_W(21, 448) <= 0; flappy_W(21, 449) <= 0; flappy_W(21, 450) <= 0; flappy_W(21, 451) <= 0; flappy_W(21, 452) <= 0; flappy_W(21, 453) <= 0; flappy_W(21, 454) <= 0; flappy_W(21, 455) <= 0; flappy_W(21, 456) <= 0; flappy_W(21, 457) <= 0; flappy_W(21, 458) <= 0; flappy_W(21, 459) <= 0; flappy_W(21, 460) <= 0; flappy_W(21, 461) <= 0; flappy_W(21, 462) <= 0; flappy_W(21, 463) <= 0; flappy_W(21, 464) <= 0; flappy_W(21, 465) <= 0; flappy_W(21, 466) <= 0; flappy_W(21, 467) <= 0; flappy_W(21, 468) <= 1; flappy_W(21, 469) <= 1; flappy_W(21, 470) <= 1; flappy_W(21, 471) <= 1; flappy_W(21, 472) <= 1; flappy_W(21, 473) <= 1; flappy_W(21, 474) <= 1; flappy_W(21, 475) <= 1; flappy_W(21, 476) <= 1; flappy_W(21, 477) <= 1; flappy_W(21, 478) <= 1; flappy_W(21, 479) <= 1; flappy_W(21, 480) <= 0; flappy_W(21, 481) <= 0; flappy_W(21, 482) <= 0; flappy_W(21, 483) <= 0; flappy_W(21, 484) <= 0; flappy_W(21, 485) <= 0; flappy_W(21, 486) <= 0; flappy_W(21, 487) <= 0; flappy_W(21, 488) <= 0; flappy_W(21, 489) <= 0; flappy_W(21, 490) <= 0; flappy_W(21, 491) <= 0; flappy_W(21, 492) <= 0; flappy_W(21, 493) <= 0; flappy_W(21, 494) <= 0; flappy_W(21, 495) <= 0; flappy_W(21, 496) <= 0; flappy_W(21, 497) <= 0; flappy_W(21, 498) <= 0; flappy_W(21, 499) <= 0; flappy_W(21, 500) <= 0; flappy_W(21, 501) <= 0; flappy_W(21, 502) <= 0; flappy_W(21, 503) <= 0; flappy_W(21, 504) <= 0; flappy_W(21, 505) <= 0; flappy_W(21, 506) <= 0; flappy_W(21, 507) <= 0; flappy_W(21, 508) <= 0; flappy_W(21, 509) <= 0; flappy_W(21, 510) <= 1; flappy_W(21, 511) <= 1; flappy_W(21, 512) <= 1; flappy_W(21, 513) <= 1; flappy_W(21, 514) <= 1; flappy_W(21, 515) <= 1; flappy_W(21, 516) <= 1; flappy_W(21, 517) <= 1; flappy_W(21, 518) <= 1; flappy_W(21, 519) <= 1; flappy_W(21, 520) <= 1; flappy_W(21, 521) <= 1; flappy_W(21, 522) <= 0; flappy_W(21, 523) <= 0; flappy_W(21, 524) <= 0; flappy_W(21, 525) <= 0; flappy_W(21, 526) <= 0; flappy_W(21, 527) <= 0; flappy_W(21, 528) <= 0; flappy_W(21, 529) <= 0; flappy_W(21, 530) <= 0; flappy_W(21, 531) <= 0; flappy_W(21, 532) <= 0; flappy_W(21, 533) <= 0; flappy_W(21, 534) <= 1; flappy_W(21, 535) <= 1; flappy_W(21, 536) <= 1; flappy_W(21, 537) <= 1; flappy_W(21, 538) <= 1; flappy_W(21, 539) <= 1; flappy_W(21, 540) <= 1; flappy_W(21, 541) <= 1; flappy_W(21, 542) <= 1; flappy_W(21, 543) <= 1; flappy_W(21, 544) <= 1; flappy_W(21, 545) <= 1; flappy_W(21, 546) <= 0; flappy_W(21, 547) <= 0; flappy_W(21, 548) <= 0; flappy_W(21, 549) <= 0; flappy_W(21, 550) <= 0; flappy_W(21, 551) <= 0; flappy_W(21, 552) <= 0; flappy_W(21, 553) <= 0; flappy_W(21, 554) <= 0; flappy_W(21, 555) <= 0; flappy_W(21, 556) <= 0; flappy_W(21, 557) <= 0; flappy_W(21, 558) <= 0; flappy_W(21, 559) <= 0; flappy_W(21, 560) <= 0; flappy_W(21, 561) <= 0; flappy_W(21, 562) <= 0; flappy_W(21, 563) <= 0; flappy_W(21, 564) <= 1; flappy_W(21, 565) <= 1; flappy_W(21, 566) <= 1; flappy_W(21, 567) <= 1; flappy_W(21, 568) <= 1; flappy_W(21, 569) <= 1; flappy_W(21, 570) <= 1; flappy_W(21, 571) <= 1; flappy_W(21, 572) <= 1; flappy_W(21, 573) <= 1; flappy_W(21, 574) <= 1; flappy_W(21, 575) <= 1; flappy_W(21, 576) <= 0; flappy_W(21, 577) <= 0; flappy_W(21, 578) <= 0; flappy_W(21, 579) <= 0; flappy_W(21, 580) <= 0; flappy_W(21, 581) <= 0; flappy_W(21, 582) <= 0; flappy_W(21, 583) <= 0; flappy_W(21, 584) <= 0; flappy_W(21, 585) <= 0; flappy_W(21, 586) <= 0; flappy_W(21, 587) <= 0; flappy_W(21, 588) <= 1; flappy_W(21, 589) <= 1; flappy_W(21, 590) <= 1; flappy_W(21, 591) <= 1; flappy_W(21, 592) <= 1; flappy_W(21, 593) <= 1; 
flappy_W(22, 0) <= 0; flappy_W(22, 1) <= 0; flappy_W(22, 2) <= 0; flappy_W(22, 3) <= 0; flappy_W(22, 4) <= 0; flappy_W(22, 5) <= 0; flappy_W(22, 6) <= 1; flappy_W(22, 7) <= 1; flappy_W(22, 8) <= 1; flappy_W(22, 9) <= 1; flappy_W(22, 10) <= 1; flappy_W(22, 11) <= 1; flappy_W(22, 12) <= 1; flappy_W(22, 13) <= 1; flappy_W(22, 14) <= 1; flappy_W(22, 15) <= 1; flappy_W(22, 16) <= 1; flappy_W(22, 17) <= 1; flappy_W(22, 18) <= 0; flappy_W(22, 19) <= 0; flappy_W(22, 20) <= 0; flappy_W(22, 21) <= 0; flappy_W(22, 22) <= 0; flappy_W(22, 23) <= 0; flappy_W(22, 24) <= 1; flappy_W(22, 25) <= 1; flappy_W(22, 26) <= 1; flappy_W(22, 27) <= 1; flappy_W(22, 28) <= 1; flappy_W(22, 29) <= 1; flappy_W(22, 30) <= 0; flappy_W(22, 31) <= 0; flappy_W(22, 32) <= 0; flappy_W(22, 33) <= 0; flappy_W(22, 34) <= 0; flappy_W(22, 35) <= 0; flappy_W(22, 36) <= 0; flappy_W(22, 37) <= 0; flappy_W(22, 38) <= 0; flappy_W(22, 39) <= 0; flappy_W(22, 40) <= 0; flappy_W(22, 41) <= 0; flappy_W(22, 42) <= 0; flappy_W(22, 43) <= 0; flappy_W(22, 44) <= 0; flappy_W(22, 45) <= 0; flappy_W(22, 46) <= 0; flappy_W(22, 47) <= 0; flappy_W(22, 48) <= 0; flappy_W(22, 49) <= 0; flappy_W(22, 50) <= 0; flappy_W(22, 51) <= 0; flappy_W(22, 52) <= 0; flappy_W(22, 53) <= 0; flappy_W(22, 54) <= 0; flappy_W(22, 55) <= 0; flappy_W(22, 56) <= 0; flappy_W(22, 57) <= 0; flappy_W(22, 58) <= 0; flappy_W(22, 59) <= 0; flappy_W(22, 60) <= 1; flappy_W(22, 61) <= 1; flappy_W(22, 62) <= 1; flappy_W(22, 63) <= 1; flappy_W(22, 64) <= 1; flappy_W(22, 65) <= 1; flappy_W(22, 66) <= 1; flappy_W(22, 67) <= 1; flappy_W(22, 68) <= 1; flappy_W(22, 69) <= 1; flappy_W(22, 70) <= 1; flappy_W(22, 71) <= 1; flappy_W(22, 72) <= 0; flappy_W(22, 73) <= 0; flappy_W(22, 74) <= 0; flappy_W(22, 75) <= 0; flappy_W(22, 76) <= 0; flappy_W(22, 77) <= 0; flappy_W(22, 78) <= 0; flappy_W(22, 79) <= 0; flappy_W(22, 80) <= 0; flappy_W(22, 81) <= 0; flappy_W(22, 82) <= 0; flappy_W(22, 83) <= 0; flappy_W(22, 84) <= 0; flappy_W(22, 85) <= 0; flappy_W(22, 86) <= 0; flappy_W(22, 87) <= 0; flappy_W(22, 88) <= 0; flappy_W(22, 89) <= 0; flappy_W(22, 90) <= 0; flappy_W(22, 91) <= 0; flappy_W(22, 92) <= 0; flappy_W(22, 93) <= 0; flappy_W(22, 94) <= 0; flappy_W(22, 95) <= 0; flappy_W(22, 96) <= 0; flappy_W(22, 97) <= 0; flappy_W(22, 98) <= 0; flappy_W(22, 99) <= 0; flappy_W(22, 100) <= 0; flappy_W(22, 101) <= 0; flappy_W(22, 102) <= 0; flappy_W(22, 103) <= 0; flappy_W(22, 104) <= 0; flappy_W(22, 105) <= 0; flappy_W(22, 106) <= 0; flappy_W(22, 107) <= 0; flappy_W(22, 108) <= 1; flappy_W(22, 109) <= 1; flappy_W(22, 110) <= 1; flappy_W(22, 111) <= 1; flappy_W(22, 112) <= 1; flappy_W(22, 113) <= 1; flappy_W(22, 114) <= 1; flappy_W(22, 115) <= 1; flappy_W(22, 116) <= 1; flappy_W(22, 117) <= 1; flappy_W(22, 118) <= 1; flappy_W(22, 119) <= 1; flappy_W(22, 120) <= 0; flappy_W(22, 121) <= 0; flappy_W(22, 122) <= 0; flappy_W(22, 123) <= 0; flappy_W(22, 124) <= 0; flappy_W(22, 125) <= 0; flappy_W(22, 126) <= 0; flappy_W(22, 127) <= 0; flappy_W(22, 128) <= 0; flappy_W(22, 129) <= 0; flappy_W(22, 130) <= 0; flappy_W(22, 131) <= 0; flappy_W(22, 132) <= 0; flappy_W(22, 133) <= 0; flappy_W(22, 134) <= 0; flappy_W(22, 135) <= 0; flappy_W(22, 136) <= 0; flappy_W(22, 137) <= 0; flappy_W(22, 138) <= 1; flappy_W(22, 139) <= 1; flappy_W(22, 140) <= 1; flappy_W(22, 141) <= 1; flappy_W(22, 142) <= 1; flappy_W(22, 143) <= 1; flappy_W(22, 144) <= 1; flappy_W(22, 145) <= 1; flappy_W(22, 146) <= 1; flappy_W(22, 147) <= 1; flappy_W(22, 148) <= 1; flappy_W(22, 149) <= 1; flappy_W(22, 150) <= 0; flappy_W(22, 151) <= 0; flappy_W(22, 152) <= 0; flappy_W(22, 153) <= 0; flappy_W(22, 154) <= 0; flappy_W(22, 155) <= 0; flappy_W(22, 156) <= 0; flappy_W(22, 157) <= 0; flappy_W(22, 158) <= 0; flappy_W(22, 159) <= 0; flappy_W(22, 160) <= 0; flappy_W(22, 161) <= 0; flappy_W(22, 162) <= 0; flappy_W(22, 163) <= 0; flappy_W(22, 164) <= 0; flappy_W(22, 165) <= 0; flappy_W(22, 166) <= 0; flappy_W(22, 167) <= 0; flappy_W(22, 168) <= 1; flappy_W(22, 169) <= 1; flappy_W(22, 170) <= 1; flappy_W(22, 171) <= 1; flappy_W(22, 172) <= 1; flappy_W(22, 173) <= 1; flappy_W(22, 174) <= 1; flappy_W(22, 175) <= 1; flappy_W(22, 176) <= 1; flappy_W(22, 177) <= 1; flappy_W(22, 178) <= 1; flappy_W(22, 179) <= 1; flappy_W(22, 180) <= 0; flappy_W(22, 181) <= 0; flappy_W(22, 182) <= 0; flappy_W(22, 183) <= 0; flappy_W(22, 184) <= 0; flappy_W(22, 185) <= 0; flappy_W(22, 186) <= 0; flappy_W(22, 187) <= 0; flappy_W(22, 188) <= 0; flappy_W(22, 189) <= 0; flappy_W(22, 190) <= 0; flappy_W(22, 191) <= 0; flappy_W(22, 192) <= 1; flappy_W(22, 193) <= 1; flappy_W(22, 194) <= 1; flappy_W(22, 195) <= 1; flappy_W(22, 196) <= 1; flappy_W(22, 197) <= 1; flappy_W(22, 198) <= 1; flappy_W(22, 199) <= 1; flappy_W(22, 200) <= 1; flappy_W(22, 201) <= 1; flappy_W(22, 202) <= 1; flappy_W(22, 203) <= 1; flappy_W(22, 204) <= 0; flappy_W(22, 205) <= 0; flappy_W(22, 206) <= 0; flappy_W(22, 207) <= 0; flappy_W(22, 208) <= 0; flappy_W(22, 209) <= 0; flappy_W(22, 210) <= 0; flappy_W(22, 211) <= 0; flappy_W(22, 212) <= 0; flappy_W(22, 213) <= 0; flappy_W(22, 214) <= 0; flappy_W(22, 215) <= 0; flappy_W(22, 216) <= 0; flappy_W(22, 217) <= 0; flappy_W(22, 218) <= 0; flappy_W(22, 219) <= 0; flappy_W(22, 220) <= 0; flappy_W(22, 221) <= 0; flappy_W(22, 222) <= 1; flappy_W(22, 223) <= 1; flappy_W(22, 224) <= 1; flappy_W(22, 225) <= 1; flappy_W(22, 226) <= 1; flappy_W(22, 227) <= 1; flappy_W(22, 228) <= 1; flappy_W(22, 229) <= 1; flappy_W(22, 230) <= 1; flappy_W(22, 231) <= 1; flappy_W(22, 232) <= 1; flappy_W(22, 233) <= 1; flappy_W(22, 234) <= 0; flappy_W(22, 235) <= 0; flappy_W(22, 236) <= 0; flappy_W(22, 237) <= 0; flappy_W(22, 238) <= 0; flappy_W(22, 239) <= 0; flappy_W(22, 240) <= 0; flappy_W(22, 241) <= 0; flappy_W(22, 242) <= 0; flappy_W(22, 243) <= 0; flappy_W(22, 244) <= 0; flappy_W(22, 245) <= 0; flappy_W(22, 246) <= 1; flappy_W(22, 247) <= 1; flappy_W(22, 248) <= 1; flappy_W(22, 249) <= 1; flappy_W(22, 250) <= 1; flappy_W(22, 251) <= 1; flappy_W(22, 252) <= 1; flappy_W(22, 253) <= 1; flappy_W(22, 254) <= 1; flappy_W(22, 255) <= 1; flappy_W(22, 256) <= 1; flappy_W(22, 257) <= 1; flappy_W(22, 258) <= 0; flappy_W(22, 259) <= 0; flappy_W(22, 260) <= 0; flappy_W(22, 261) <= 0; flappy_W(22, 262) <= 0; flappy_W(22, 263) <= 0; flappy_W(22, 264) <= 0; flappy_W(22, 265) <= 0; flappy_W(22, 266) <= 0; flappy_W(22, 267) <= 0; flappy_W(22, 268) <= 0; flappy_W(22, 269) <= 0; flappy_W(22, 270) <= 0; flappy_W(22, 271) <= 0; flappy_W(22, 272) <= 0; flappy_W(22, 273) <= 0; flappy_W(22, 274) <= 0; flappy_W(22, 275) <= 0; flappy_W(22, 276) <= 1; flappy_W(22, 277) <= 1; flappy_W(22, 278) <= 1; flappy_W(22, 279) <= 1; flappy_W(22, 280) <= 1; flappy_W(22, 281) <= 1; flappy_W(22, 282) <= 1; flappy_W(22, 283) <= 1; flappy_W(22, 284) <= 1; flappy_W(22, 285) <= 1; flappy_W(22, 286) <= 1; flappy_W(22, 287) <= 1; flappy_W(22, 288) <= 0; flappy_W(22, 289) <= 0; flappy_W(22, 290) <= 0; flappy_W(22, 291) <= 0; flappy_W(22, 292) <= 0; flappy_W(22, 293) <= 0; flappy_W(22, 294) <= 0; flappy_W(22, 295) <= 0; flappy_W(22, 296) <= 0; flappy_W(22, 297) <= 0; flappy_W(22, 298) <= 0; flappy_W(22, 299) <= 0; flappy_W(22, 300) <= 1; flappy_W(22, 301) <= 1; flappy_W(22, 302) <= 1; flappy_W(22, 303) <= 1; flappy_W(22, 304) <= 1; flappy_W(22, 305) <= 1; flappy_W(22, 306) <= 1; flappy_W(22, 307) <= 1; flappy_W(22, 308) <= 1; flappy_W(22, 309) <= 1; flappy_W(22, 310) <= 1; flappy_W(22, 311) <= 1; flappy_W(22, 312) <= 0; flappy_W(22, 313) <= 0; flappy_W(22, 314) <= 0; flappy_W(22, 315) <= 0; flappy_W(22, 316) <= 0; flappy_W(22, 317) <= 0; flappy_W(22, 318) <= 0; flappy_W(22, 319) <= 0; flappy_W(22, 320) <= 0; flappy_W(22, 321) <= 0; flappy_W(22, 322) <= 0; flappy_W(22, 323) <= 0; flappy_W(22, 324) <= 0; flappy_W(22, 325) <= 0; flappy_W(22, 326) <= 0; flappy_W(22, 327) <= 0; flappy_W(22, 328) <= 0; flappy_W(22, 329) <= 0; flappy_W(22, 330) <= 0; flappy_W(22, 331) <= 0; flappy_W(22, 332) <= 0; flappy_W(22, 333) <= 0; flappy_W(22, 334) <= 0; flappy_W(22, 335) <= 0; flappy_W(22, 336) <= 0; flappy_W(22, 337) <= 0; flappy_W(22, 338) <= 0; flappy_W(22, 339) <= 0; flappy_W(22, 340) <= 0; flappy_W(22, 341) <= 0; flappy_W(22, 342) <= 0; flappy_W(22, 343) <= 0; flappy_W(22, 344) <= 0; flappy_W(22, 345) <= 0; flappy_W(22, 346) <= 0; flappy_W(22, 347) <= 0; flappy_W(22, 348) <= 0; flappy_W(22, 349) <= 0; flappy_W(22, 350) <= 0; flappy_W(22, 351) <= 0; flappy_W(22, 352) <= 0; flappy_W(22, 353) <= 0; flappy_W(22, 354) <= 0; flappy_W(22, 355) <= 0; flappy_W(22, 356) <= 0; flappy_W(22, 357) <= 0; flappy_W(22, 358) <= 0; flappy_W(22, 359) <= 0; flappy_W(22, 360) <= 0; flappy_W(22, 361) <= 0; flappy_W(22, 362) <= 0; flappy_W(22, 363) <= 0; flappy_W(22, 364) <= 0; flappy_W(22, 365) <= 0; flappy_W(22, 366) <= 0; flappy_W(22, 367) <= 0; flappy_W(22, 368) <= 0; flappy_W(22, 369) <= 0; flappy_W(22, 370) <= 0; flappy_W(22, 371) <= 0; flappy_W(22, 372) <= 0; flappy_W(22, 373) <= 0; flappy_W(22, 374) <= 0; flappy_W(22, 375) <= 0; flappy_W(22, 376) <= 0; flappy_W(22, 377) <= 0; flappy_W(22, 378) <= 0; flappy_W(22, 379) <= 0; flappy_W(22, 380) <= 0; flappy_W(22, 381) <= 0; flappy_W(22, 382) <= 0; flappy_W(22, 383) <= 0; flappy_W(22, 384) <= 0; flappy_W(22, 385) <= 0; flappy_W(22, 386) <= 0; flappy_W(22, 387) <= 0; flappy_W(22, 388) <= 0; flappy_W(22, 389) <= 0; flappy_W(22, 390) <= 0; flappy_W(22, 391) <= 0; flappy_W(22, 392) <= 0; flappy_W(22, 393) <= 0; flappy_W(22, 394) <= 0; flappy_W(22, 395) <= 0; flappy_W(22, 396) <= 0; flappy_W(22, 397) <= 0; flappy_W(22, 398) <= 0; flappy_W(22, 399) <= 0; flappy_W(22, 400) <= 0; flappy_W(22, 401) <= 0; flappy_W(22, 402) <= 1; flappy_W(22, 403) <= 1; flappy_W(22, 404) <= 1; flappy_W(22, 405) <= 1; flappy_W(22, 406) <= 1; flappy_W(22, 407) <= 1; flappy_W(22, 408) <= 1; flappy_W(22, 409) <= 1; flappy_W(22, 410) <= 1; flappy_W(22, 411) <= 1; flappy_W(22, 412) <= 1; flappy_W(22, 413) <= 1; flappy_W(22, 414) <= 0; flappy_W(22, 415) <= 0; flappy_W(22, 416) <= 0; flappy_W(22, 417) <= 0; flappy_W(22, 418) <= 0; flappy_W(22, 419) <= 0; flappy_W(22, 420) <= 0; flappy_W(22, 421) <= 0; flappy_W(22, 422) <= 0; flappy_W(22, 423) <= 0; flappy_W(22, 424) <= 0; flappy_W(22, 425) <= 0; flappy_W(22, 426) <= 1; flappy_W(22, 427) <= 1; flappy_W(22, 428) <= 1; flappy_W(22, 429) <= 1; flappy_W(22, 430) <= 1; flappy_W(22, 431) <= 1; flappy_W(22, 432) <= 1; flappy_W(22, 433) <= 1; flappy_W(22, 434) <= 1; flappy_W(22, 435) <= 1; flappy_W(22, 436) <= 1; flappy_W(22, 437) <= 1; flappy_W(22, 438) <= 0; flappy_W(22, 439) <= 0; flappy_W(22, 440) <= 0; flappy_W(22, 441) <= 0; flappy_W(22, 442) <= 0; flappy_W(22, 443) <= 0; flappy_W(22, 444) <= 0; flappy_W(22, 445) <= 0; flappy_W(22, 446) <= 0; flappy_W(22, 447) <= 0; flappy_W(22, 448) <= 0; flappy_W(22, 449) <= 0; flappy_W(22, 450) <= 0; flappy_W(22, 451) <= 0; flappy_W(22, 452) <= 0; flappy_W(22, 453) <= 0; flappy_W(22, 454) <= 0; flappy_W(22, 455) <= 0; flappy_W(22, 456) <= 0; flappy_W(22, 457) <= 0; flappy_W(22, 458) <= 0; flappy_W(22, 459) <= 0; flappy_W(22, 460) <= 0; flappy_W(22, 461) <= 0; flappy_W(22, 462) <= 0; flappy_W(22, 463) <= 0; flappy_W(22, 464) <= 0; flappy_W(22, 465) <= 0; flappy_W(22, 466) <= 0; flappy_W(22, 467) <= 0; flappy_W(22, 468) <= 1; flappy_W(22, 469) <= 1; flappy_W(22, 470) <= 1; flappy_W(22, 471) <= 1; flappy_W(22, 472) <= 1; flappy_W(22, 473) <= 1; flappy_W(22, 474) <= 1; flappy_W(22, 475) <= 1; flappy_W(22, 476) <= 1; flappy_W(22, 477) <= 1; flappy_W(22, 478) <= 1; flappy_W(22, 479) <= 1; flappy_W(22, 480) <= 0; flappy_W(22, 481) <= 0; flappy_W(22, 482) <= 0; flappy_W(22, 483) <= 0; flappy_W(22, 484) <= 0; flappy_W(22, 485) <= 0; flappy_W(22, 486) <= 0; flappy_W(22, 487) <= 0; flappy_W(22, 488) <= 0; flappy_W(22, 489) <= 0; flappy_W(22, 490) <= 0; flappy_W(22, 491) <= 0; flappy_W(22, 492) <= 0; flappy_W(22, 493) <= 0; flappy_W(22, 494) <= 0; flappy_W(22, 495) <= 0; flappy_W(22, 496) <= 0; flappy_W(22, 497) <= 0; flappy_W(22, 498) <= 0; flappy_W(22, 499) <= 0; flappy_W(22, 500) <= 0; flappy_W(22, 501) <= 0; flappy_W(22, 502) <= 0; flappy_W(22, 503) <= 0; flappy_W(22, 504) <= 0; flappy_W(22, 505) <= 0; flappy_W(22, 506) <= 0; flappy_W(22, 507) <= 0; flappy_W(22, 508) <= 0; flappy_W(22, 509) <= 0; flappy_W(22, 510) <= 1; flappy_W(22, 511) <= 1; flappy_W(22, 512) <= 1; flappy_W(22, 513) <= 1; flappy_W(22, 514) <= 1; flappy_W(22, 515) <= 1; flappy_W(22, 516) <= 1; flappy_W(22, 517) <= 1; flappy_W(22, 518) <= 1; flappy_W(22, 519) <= 1; flappy_W(22, 520) <= 1; flappy_W(22, 521) <= 1; flappy_W(22, 522) <= 0; flappy_W(22, 523) <= 0; flappy_W(22, 524) <= 0; flappy_W(22, 525) <= 0; flappy_W(22, 526) <= 0; flappy_W(22, 527) <= 0; flappy_W(22, 528) <= 0; flappy_W(22, 529) <= 0; flappy_W(22, 530) <= 0; flappy_W(22, 531) <= 0; flappy_W(22, 532) <= 0; flappy_W(22, 533) <= 0; flappy_W(22, 534) <= 1; flappy_W(22, 535) <= 1; flappy_W(22, 536) <= 1; flappy_W(22, 537) <= 1; flappy_W(22, 538) <= 1; flappy_W(22, 539) <= 1; flappy_W(22, 540) <= 1; flappy_W(22, 541) <= 1; flappy_W(22, 542) <= 1; flappy_W(22, 543) <= 1; flappy_W(22, 544) <= 1; flappy_W(22, 545) <= 1; flappy_W(22, 546) <= 0; flappy_W(22, 547) <= 0; flappy_W(22, 548) <= 0; flappy_W(22, 549) <= 0; flappy_W(22, 550) <= 0; flappy_W(22, 551) <= 0; flappy_W(22, 552) <= 0; flappy_W(22, 553) <= 0; flappy_W(22, 554) <= 0; flappy_W(22, 555) <= 0; flappy_W(22, 556) <= 0; flappy_W(22, 557) <= 0; flappy_W(22, 558) <= 0; flappy_W(22, 559) <= 0; flappy_W(22, 560) <= 0; flappy_W(22, 561) <= 0; flappy_W(22, 562) <= 0; flappy_W(22, 563) <= 0; flappy_W(22, 564) <= 1; flappy_W(22, 565) <= 1; flappy_W(22, 566) <= 1; flappy_W(22, 567) <= 1; flappy_W(22, 568) <= 1; flappy_W(22, 569) <= 1; flappy_W(22, 570) <= 1; flappy_W(22, 571) <= 1; flappy_W(22, 572) <= 1; flappy_W(22, 573) <= 1; flappy_W(22, 574) <= 1; flappy_W(22, 575) <= 1; flappy_W(22, 576) <= 0; flappy_W(22, 577) <= 0; flappy_W(22, 578) <= 0; flappy_W(22, 579) <= 0; flappy_W(22, 580) <= 0; flappy_W(22, 581) <= 0; flappy_W(22, 582) <= 0; flappy_W(22, 583) <= 0; flappy_W(22, 584) <= 0; flappy_W(22, 585) <= 0; flappy_W(22, 586) <= 0; flappy_W(22, 587) <= 0; flappy_W(22, 588) <= 1; flappy_W(22, 589) <= 1; flappy_W(22, 590) <= 1; flappy_W(22, 591) <= 1; flappy_W(22, 592) <= 1; flappy_W(22, 593) <= 1; 
flappy_W(23, 0) <= 0; flappy_W(23, 1) <= 0; flappy_W(23, 2) <= 0; flappy_W(23, 3) <= 0; flappy_W(23, 4) <= 0; flappy_W(23, 5) <= 0; flappy_W(23, 6) <= 1; flappy_W(23, 7) <= 1; flappy_W(23, 8) <= 1; flappy_W(23, 9) <= 1; flappy_W(23, 10) <= 1; flappy_W(23, 11) <= 1; flappy_W(23, 12) <= 1; flappy_W(23, 13) <= 1; flappy_W(23, 14) <= 1; flappy_W(23, 15) <= 1; flappy_W(23, 16) <= 1; flappy_W(23, 17) <= 1; flappy_W(23, 18) <= 0; flappy_W(23, 19) <= 0; flappy_W(23, 20) <= 0; flappy_W(23, 21) <= 0; flappy_W(23, 22) <= 0; flappy_W(23, 23) <= 0; flappy_W(23, 24) <= 1; flappy_W(23, 25) <= 1; flappy_W(23, 26) <= 1; flappy_W(23, 27) <= 1; flappy_W(23, 28) <= 1; flappy_W(23, 29) <= 1; flappy_W(23, 30) <= 0; flappy_W(23, 31) <= 0; flappy_W(23, 32) <= 0; flappy_W(23, 33) <= 0; flappy_W(23, 34) <= 0; flappy_W(23, 35) <= 0; flappy_W(23, 36) <= 0; flappy_W(23, 37) <= 0; flappy_W(23, 38) <= 0; flappy_W(23, 39) <= 0; flappy_W(23, 40) <= 0; flappy_W(23, 41) <= 0; flappy_W(23, 42) <= 0; flappy_W(23, 43) <= 0; flappy_W(23, 44) <= 0; flappy_W(23, 45) <= 0; flappy_W(23, 46) <= 0; flappy_W(23, 47) <= 0; flappy_W(23, 48) <= 0; flappy_W(23, 49) <= 0; flappy_W(23, 50) <= 0; flappy_W(23, 51) <= 0; flappy_W(23, 52) <= 0; flappy_W(23, 53) <= 0; flappy_W(23, 54) <= 0; flappy_W(23, 55) <= 0; flappy_W(23, 56) <= 0; flappy_W(23, 57) <= 0; flappy_W(23, 58) <= 0; flappy_W(23, 59) <= 0; flappy_W(23, 60) <= 1; flappy_W(23, 61) <= 1; flappy_W(23, 62) <= 1; flappy_W(23, 63) <= 1; flappy_W(23, 64) <= 1; flappy_W(23, 65) <= 1; flappy_W(23, 66) <= 1; flappy_W(23, 67) <= 1; flappy_W(23, 68) <= 1; flappy_W(23, 69) <= 1; flappy_W(23, 70) <= 1; flappy_W(23, 71) <= 1; flappy_W(23, 72) <= 0; flappy_W(23, 73) <= 0; flappy_W(23, 74) <= 0; flappy_W(23, 75) <= 0; flappy_W(23, 76) <= 0; flappy_W(23, 77) <= 0; flappy_W(23, 78) <= 0; flappy_W(23, 79) <= 0; flappy_W(23, 80) <= 0; flappy_W(23, 81) <= 0; flappy_W(23, 82) <= 0; flappy_W(23, 83) <= 0; flappy_W(23, 84) <= 0; flappy_W(23, 85) <= 0; flappy_W(23, 86) <= 0; flappy_W(23, 87) <= 0; flappy_W(23, 88) <= 0; flappy_W(23, 89) <= 0; flappy_W(23, 90) <= 0; flappy_W(23, 91) <= 0; flappy_W(23, 92) <= 0; flappy_W(23, 93) <= 0; flappy_W(23, 94) <= 0; flappy_W(23, 95) <= 0; flappy_W(23, 96) <= 0; flappy_W(23, 97) <= 0; flappy_W(23, 98) <= 0; flappy_W(23, 99) <= 0; flappy_W(23, 100) <= 0; flappy_W(23, 101) <= 0; flappy_W(23, 102) <= 0; flappy_W(23, 103) <= 0; flappy_W(23, 104) <= 0; flappy_W(23, 105) <= 0; flappy_W(23, 106) <= 0; flappy_W(23, 107) <= 0; flappy_W(23, 108) <= 1; flappy_W(23, 109) <= 1; flappy_W(23, 110) <= 1; flappy_W(23, 111) <= 1; flappy_W(23, 112) <= 1; flappy_W(23, 113) <= 1; flappy_W(23, 114) <= 1; flappy_W(23, 115) <= 1; flappy_W(23, 116) <= 1; flappy_W(23, 117) <= 1; flappy_W(23, 118) <= 1; flappy_W(23, 119) <= 1; flappy_W(23, 120) <= 0; flappy_W(23, 121) <= 0; flappy_W(23, 122) <= 0; flappy_W(23, 123) <= 0; flappy_W(23, 124) <= 0; flappy_W(23, 125) <= 0; flappy_W(23, 126) <= 0; flappy_W(23, 127) <= 0; flappy_W(23, 128) <= 0; flappy_W(23, 129) <= 0; flappy_W(23, 130) <= 0; flappy_W(23, 131) <= 0; flappy_W(23, 132) <= 0; flappy_W(23, 133) <= 0; flappy_W(23, 134) <= 0; flappy_W(23, 135) <= 0; flappy_W(23, 136) <= 0; flappy_W(23, 137) <= 0; flappy_W(23, 138) <= 1; flappy_W(23, 139) <= 1; flappy_W(23, 140) <= 1; flappy_W(23, 141) <= 1; flappy_W(23, 142) <= 1; flappy_W(23, 143) <= 1; flappy_W(23, 144) <= 1; flappy_W(23, 145) <= 1; flappy_W(23, 146) <= 1; flappy_W(23, 147) <= 1; flappy_W(23, 148) <= 1; flappy_W(23, 149) <= 1; flappy_W(23, 150) <= 0; flappy_W(23, 151) <= 0; flappy_W(23, 152) <= 0; flappy_W(23, 153) <= 0; flappy_W(23, 154) <= 0; flappy_W(23, 155) <= 0; flappy_W(23, 156) <= 0; flappy_W(23, 157) <= 0; flappy_W(23, 158) <= 0; flappy_W(23, 159) <= 0; flappy_W(23, 160) <= 0; flappy_W(23, 161) <= 0; flappy_W(23, 162) <= 0; flappy_W(23, 163) <= 0; flappy_W(23, 164) <= 0; flappy_W(23, 165) <= 0; flappy_W(23, 166) <= 0; flappy_W(23, 167) <= 0; flappy_W(23, 168) <= 1; flappy_W(23, 169) <= 1; flappy_W(23, 170) <= 1; flappy_W(23, 171) <= 1; flappy_W(23, 172) <= 1; flappy_W(23, 173) <= 1; flappy_W(23, 174) <= 1; flappy_W(23, 175) <= 1; flappy_W(23, 176) <= 1; flappy_W(23, 177) <= 1; flappy_W(23, 178) <= 1; flappy_W(23, 179) <= 1; flappy_W(23, 180) <= 0; flappy_W(23, 181) <= 0; flappy_W(23, 182) <= 0; flappy_W(23, 183) <= 0; flappy_W(23, 184) <= 0; flappy_W(23, 185) <= 0; flappy_W(23, 186) <= 0; flappy_W(23, 187) <= 0; flappy_W(23, 188) <= 0; flappy_W(23, 189) <= 0; flappy_W(23, 190) <= 0; flappy_W(23, 191) <= 0; flappy_W(23, 192) <= 1; flappy_W(23, 193) <= 1; flappy_W(23, 194) <= 1; flappy_W(23, 195) <= 1; flappy_W(23, 196) <= 1; flappy_W(23, 197) <= 1; flappy_W(23, 198) <= 1; flappy_W(23, 199) <= 1; flappy_W(23, 200) <= 1; flappy_W(23, 201) <= 1; flappy_W(23, 202) <= 1; flappy_W(23, 203) <= 1; flappy_W(23, 204) <= 0; flappy_W(23, 205) <= 0; flappy_W(23, 206) <= 0; flappy_W(23, 207) <= 0; flappy_W(23, 208) <= 0; flappy_W(23, 209) <= 0; flappy_W(23, 210) <= 0; flappy_W(23, 211) <= 0; flappy_W(23, 212) <= 0; flappy_W(23, 213) <= 0; flappy_W(23, 214) <= 0; flappy_W(23, 215) <= 0; flappy_W(23, 216) <= 0; flappy_W(23, 217) <= 0; flappy_W(23, 218) <= 0; flappy_W(23, 219) <= 0; flappy_W(23, 220) <= 0; flappy_W(23, 221) <= 0; flappy_W(23, 222) <= 1; flappy_W(23, 223) <= 1; flappy_W(23, 224) <= 1; flappy_W(23, 225) <= 1; flappy_W(23, 226) <= 1; flappy_W(23, 227) <= 1; flappy_W(23, 228) <= 1; flappy_W(23, 229) <= 1; flappy_W(23, 230) <= 1; flappy_W(23, 231) <= 1; flappy_W(23, 232) <= 1; flappy_W(23, 233) <= 1; flappy_W(23, 234) <= 0; flappy_W(23, 235) <= 0; flappy_W(23, 236) <= 0; flappy_W(23, 237) <= 0; flappy_W(23, 238) <= 0; flappy_W(23, 239) <= 0; flappy_W(23, 240) <= 0; flappy_W(23, 241) <= 0; flappy_W(23, 242) <= 0; flappy_W(23, 243) <= 0; flappy_W(23, 244) <= 0; flappy_W(23, 245) <= 0; flappy_W(23, 246) <= 1; flappy_W(23, 247) <= 1; flappy_W(23, 248) <= 1; flappy_W(23, 249) <= 1; flappy_W(23, 250) <= 1; flappy_W(23, 251) <= 1; flappy_W(23, 252) <= 1; flappy_W(23, 253) <= 1; flappy_W(23, 254) <= 1; flappy_W(23, 255) <= 1; flappy_W(23, 256) <= 1; flappy_W(23, 257) <= 1; flappy_W(23, 258) <= 0; flappy_W(23, 259) <= 0; flappy_W(23, 260) <= 0; flappy_W(23, 261) <= 0; flappy_W(23, 262) <= 0; flappy_W(23, 263) <= 0; flappy_W(23, 264) <= 0; flappy_W(23, 265) <= 0; flappy_W(23, 266) <= 0; flappy_W(23, 267) <= 0; flappy_W(23, 268) <= 0; flappy_W(23, 269) <= 0; flappy_W(23, 270) <= 0; flappy_W(23, 271) <= 0; flappy_W(23, 272) <= 0; flappy_W(23, 273) <= 0; flappy_W(23, 274) <= 0; flappy_W(23, 275) <= 0; flappy_W(23, 276) <= 1; flappy_W(23, 277) <= 1; flappy_W(23, 278) <= 1; flappy_W(23, 279) <= 1; flappy_W(23, 280) <= 1; flappy_W(23, 281) <= 1; flappy_W(23, 282) <= 1; flappy_W(23, 283) <= 1; flappy_W(23, 284) <= 1; flappy_W(23, 285) <= 1; flappy_W(23, 286) <= 1; flappy_W(23, 287) <= 1; flappy_W(23, 288) <= 0; flappy_W(23, 289) <= 0; flappy_W(23, 290) <= 0; flappy_W(23, 291) <= 0; flappy_W(23, 292) <= 0; flappy_W(23, 293) <= 0; flappy_W(23, 294) <= 0; flappy_W(23, 295) <= 0; flappy_W(23, 296) <= 0; flappy_W(23, 297) <= 0; flappy_W(23, 298) <= 0; flappy_W(23, 299) <= 0; flappy_W(23, 300) <= 1; flappy_W(23, 301) <= 1; flappy_W(23, 302) <= 1; flappy_W(23, 303) <= 1; flappy_W(23, 304) <= 1; flappy_W(23, 305) <= 1; flappy_W(23, 306) <= 1; flappy_W(23, 307) <= 1; flappy_W(23, 308) <= 1; flappy_W(23, 309) <= 1; flappy_W(23, 310) <= 1; flappy_W(23, 311) <= 1; flappy_W(23, 312) <= 0; flappy_W(23, 313) <= 0; flappy_W(23, 314) <= 0; flappy_W(23, 315) <= 0; flappy_W(23, 316) <= 0; flappy_W(23, 317) <= 0; flappy_W(23, 318) <= 0; flappy_W(23, 319) <= 0; flappy_W(23, 320) <= 0; flappy_W(23, 321) <= 0; flappy_W(23, 322) <= 0; flappy_W(23, 323) <= 0; flappy_W(23, 324) <= 0; flappy_W(23, 325) <= 0; flappy_W(23, 326) <= 0; flappy_W(23, 327) <= 0; flappy_W(23, 328) <= 0; flappy_W(23, 329) <= 0; flappy_W(23, 330) <= 0; flappy_W(23, 331) <= 0; flappy_W(23, 332) <= 0; flappy_W(23, 333) <= 0; flappy_W(23, 334) <= 0; flappy_W(23, 335) <= 0; flappy_W(23, 336) <= 0; flappy_W(23, 337) <= 0; flappy_W(23, 338) <= 0; flappy_W(23, 339) <= 0; flappy_W(23, 340) <= 0; flappy_W(23, 341) <= 0; flappy_W(23, 342) <= 0; flappy_W(23, 343) <= 0; flappy_W(23, 344) <= 0; flappy_W(23, 345) <= 0; flappy_W(23, 346) <= 0; flappy_W(23, 347) <= 0; flappy_W(23, 348) <= 0; flappy_W(23, 349) <= 0; flappy_W(23, 350) <= 0; flappy_W(23, 351) <= 0; flappy_W(23, 352) <= 0; flappy_W(23, 353) <= 0; flappy_W(23, 354) <= 0; flappy_W(23, 355) <= 0; flappy_W(23, 356) <= 0; flappy_W(23, 357) <= 0; flappy_W(23, 358) <= 0; flappy_W(23, 359) <= 0; flappy_W(23, 360) <= 0; flappy_W(23, 361) <= 0; flappy_W(23, 362) <= 0; flappy_W(23, 363) <= 0; flappy_W(23, 364) <= 0; flappy_W(23, 365) <= 0; flappy_W(23, 366) <= 0; flappy_W(23, 367) <= 0; flappy_W(23, 368) <= 0; flappy_W(23, 369) <= 0; flappy_W(23, 370) <= 0; flappy_W(23, 371) <= 0; flappy_W(23, 372) <= 0; flappy_W(23, 373) <= 0; flappy_W(23, 374) <= 0; flappy_W(23, 375) <= 0; flappy_W(23, 376) <= 0; flappy_W(23, 377) <= 0; flappy_W(23, 378) <= 0; flappy_W(23, 379) <= 0; flappy_W(23, 380) <= 0; flappy_W(23, 381) <= 0; flappy_W(23, 382) <= 0; flappy_W(23, 383) <= 0; flappy_W(23, 384) <= 0; flappy_W(23, 385) <= 0; flappy_W(23, 386) <= 0; flappy_W(23, 387) <= 0; flappy_W(23, 388) <= 0; flappy_W(23, 389) <= 0; flappy_W(23, 390) <= 0; flappy_W(23, 391) <= 0; flappy_W(23, 392) <= 0; flappy_W(23, 393) <= 0; flappy_W(23, 394) <= 0; flappy_W(23, 395) <= 0; flappy_W(23, 396) <= 0; flappy_W(23, 397) <= 0; flappy_W(23, 398) <= 0; flappy_W(23, 399) <= 0; flappy_W(23, 400) <= 0; flappy_W(23, 401) <= 0; flappy_W(23, 402) <= 1; flappy_W(23, 403) <= 1; flappy_W(23, 404) <= 1; flappy_W(23, 405) <= 1; flappy_W(23, 406) <= 1; flappy_W(23, 407) <= 1; flappy_W(23, 408) <= 1; flappy_W(23, 409) <= 1; flappy_W(23, 410) <= 1; flappy_W(23, 411) <= 1; flappy_W(23, 412) <= 1; flappy_W(23, 413) <= 1; flappy_W(23, 414) <= 0; flappy_W(23, 415) <= 0; flappy_W(23, 416) <= 0; flappy_W(23, 417) <= 0; flappy_W(23, 418) <= 0; flappy_W(23, 419) <= 0; flappy_W(23, 420) <= 0; flappy_W(23, 421) <= 0; flappy_W(23, 422) <= 0; flappy_W(23, 423) <= 0; flappy_W(23, 424) <= 0; flappy_W(23, 425) <= 0; flappy_W(23, 426) <= 1; flappy_W(23, 427) <= 1; flappy_W(23, 428) <= 1; flappy_W(23, 429) <= 1; flappy_W(23, 430) <= 1; flappy_W(23, 431) <= 1; flappy_W(23, 432) <= 1; flappy_W(23, 433) <= 1; flappy_W(23, 434) <= 1; flappy_W(23, 435) <= 1; flappy_W(23, 436) <= 1; flappy_W(23, 437) <= 1; flappy_W(23, 438) <= 0; flappy_W(23, 439) <= 0; flappy_W(23, 440) <= 0; flappy_W(23, 441) <= 0; flappy_W(23, 442) <= 0; flappy_W(23, 443) <= 0; flappy_W(23, 444) <= 0; flappy_W(23, 445) <= 0; flappy_W(23, 446) <= 0; flappy_W(23, 447) <= 0; flappy_W(23, 448) <= 0; flappy_W(23, 449) <= 0; flappy_W(23, 450) <= 0; flappy_W(23, 451) <= 0; flappy_W(23, 452) <= 0; flappy_W(23, 453) <= 0; flappy_W(23, 454) <= 0; flappy_W(23, 455) <= 0; flappy_W(23, 456) <= 0; flappy_W(23, 457) <= 0; flappy_W(23, 458) <= 0; flappy_W(23, 459) <= 0; flappy_W(23, 460) <= 0; flappy_W(23, 461) <= 0; flappy_W(23, 462) <= 0; flappy_W(23, 463) <= 0; flappy_W(23, 464) <= 0; flappy_W(23, 465) <= 0; flappy_W(23, 466) <= 0; flappy_W(23, 467) <= 0; flappy_W(23, 468) <= 1; flappy_W(23, 469) <= 1; flappy_W(23, 470) <= 1; flappy_W(23, 471) <= 1; flappy_W(23, 472) <= 1; flappy_W(23, 473) <= 1; flappy_W(23, 474) <= 1; flappy_W(23, 475) <= 1; flappy_W(23, 476) <= 1; flappy_W(23, 477) <= 1; flappy_W(23, 478) <= 1; flappy_W(23, 479) <= 1; flappy_W(23, 480) <= 0; flappy_W(23, 481) <= 0; flappy_W(23, 482) <= 0; flappy_W(23, 483) <= 0; flappy_W(23, 484) <= 0; flappy_W(23, 485) <= 0; flappy_W(23, 486) <= 0; flappy_W(23, 487) <= 0; flappy_W(23, 488) <= 0; flappy_W(23, 489) <= 0; flappy_W(23, 490) <= 0; flappy_W(23, 491) <= 0; flappy_W(23, 492) <= 0; flappy_W(23, 493) <= 0; flappy_W(23, 494) <= 0; flappy_W(23, 495) <= 0; flappy_W(23, 496) <= 0; flappy_W(23, 497) <= 0; flappy_W(23, 498) <= 0; flappy_W(23, 499) <= 0; flappy_W(23, 500) <= 0; flappy_W(23, 501) <= 0; flappy_W(23, 502) <= 0; flappy_W(23, 503) <= 0; flappy_W(23, 504) <= 0; flappy_W(23, 505) <= 0; flappy_W(23, 506) <= 0; flappy_W(23, 507) <= 0; flappy_W(23, 508) <= 0; flappy_W(23, 509) <= 0; flappy_W(23, 510) <= 1; flappy_W(23, 511) <= 1; flappy_W(23, 512) <= 1; flappy_W(23, 513) <= 1; flappy_W(23, 514) <= 1; flappy_W(23, 515) <= 1; flappy_W(23, 516) <= 1; flappy_W(23, 517) <= 1; flappy_W(23, 518) <= 1; flappy_W(23, 519) <= 1; flappy_W(23, 520) <= 1; flappy_W(23, 521) <= 1; flappy_W(23, 522) <= 0; flappy_W(23, 523) <= 0; flappy_W(23, 524) <= 0; flappy_W(23, 525) <= 0; flappy_W(23, 526) <= 0; flappy_W(23, 527) <= 0; flappy_W(23, 528) <= 0; flappy_W(23, 529) <= 0; flappy_W(23, 530) <= 0; flappy_W(23, 531) <= 0; flappy_W(23, 532) <= 0; flappy_W(23, 533) <= 0; flappy_W(23, 534) <= 1; flappy_W(23, 535) <= 1; flappy_W(23, 536) <= 1; flappy_W(23, 537) <= 1; flappy_W(23, 538) <= 1; flappy_W(23, 539) <= 1; flappy_W(23, 540) <= 1; flappy_W(23, 541) <= 1; flappy_W(23, 542) <= 1; flappy_W(23, 543) <= 1; flappy_W(23, 544) <= 1; flappy_W(23, 545) <= 1; flappy_W(23, 546) <= 0; flappy_W(23, 547) <= 0; flappy_W(23, 548) <= 0; flappy_W(23, 549) <= 0; flappy_W(23, 550) <= 0; flappy_W(23, 551) <= 0; flappy_W(23, 552) <= 0; flappy_W(23, 553) <= 0; flappy_W(23, 554) <= 0; flappy_W(23, 555) <= 0; flappy_W(23, 556) <= 0; flappy_W(23, 557) <= 0; flappy_W(23, 558) <= 0; flappy_W(23, 559) <= 0; flappy_W(23, 560) <= 0; flappy_W(23, 561) <= 0; flappy_W(23, 562) <= 0; flappy_W(23, 563) <= 0; flappy_W(23, 564) <= 1; flappy_W(23, 565) <= 1; flappy_W(23, 566) <= 1; flappy_W(23, 567) <= 1; flappy_W(23, 568) <= 1; flappy_W(23, 569) <= 1; flappy_W(23, 570) <= 1; flappy_W(23, 571) <= 1; flappy_W(23, 572) <= 1; flappy_W(23, 573) <= 1; flappy_W(23, 574) <= 1; flappy_W(23, 575) <= 1; flappy_W(23, 576) <= 0; flappy_W(23, 577) <= 0; flappy_W(23, 578) <= 0; flappy_W(23, 579) <= 0; flappy_W(23, 580) <= 0; flappy_W(23, 581) <= 0; flappy_W(23, 582) <= 0; flappy_W(23, 583) <= 0; flappy_W(23, 584) <= 0; flappy_W(23, 585) <= 0; flappy_W(23, 586) <= 0; flappy_W(23, 587) <= 0; flappy_W(23, 588) <= 1; flappy_W(23, 589) <= 1; flappy_W(23, 590) <= 1; flappy_W(23, 591) <= 1; flappy_W(23, 592) <= 1; flappy_W(23, 593) <= 1; 
flappy_W(24, 0) <= 0; flappy_W(24, 1) <= 0; flappy_W(24, 2) <= 0; flappy_W(24, 3) <= 0; flappy_W(24, 4) <= 0; flappy_W(24, 5) <= 0; flappy_W(24, 6) <= 1; flappy_W(24, 7) <= 1; flappy_W(24, 8) <= 1; flappy_W(24, 9) <= 1; flappy_W(24, 10) <= 1; flappy_W(24, 11) <= 1; flappy_W(24, 12) <= 1; flappy_W(24, 13) <= 1; flappy_W(24, 14) <= 1; flappy_W(24, 15) <= 1; flappy_W(24, 16) <= 1; flappy_W(24, 17) <= 1; flappy_W(24, 18) <= 1; flappy_W(24, 19) <= 1; flappy_W(24, 20) <= 1; flappy_W(24, 21) <= 1; flappy_W(24, 22) <= 1; flappy_W(24, 23) <= 1; flappy_W(24, 24) <= 1; flappy_W(24, 25) <= 1; flappy_W(24, 26) <= 1; flappy_W(24, 27) <= 1; flappy_W(24, 28) <= 1; flappy_W(24, 29) <= 1; flappy_W(24, 30) <= 0; flappy_W(24, 31) <= 0; flappy_W(24, 32) <= 0; flappy_W(24, 33) <= 0; flappy_W(24, 34) <= 0; flappy_W(24, 35) <= 0; flappy_W(24, 36) <= 0; flappy_W(24, 37) <= 0; flappy_W(24, 38) <= 0; flappy_W(24, 39) <= 0; flappy_W(24, 40) <= 0; flappy_W(24, 41) <= 0; flappy_W(24, 42) <= 0; flappy_W(24, 43) <= 0; flappy_W(24, 44) <= 0; flappy_W(24, 45) <= 0; flappy_W(24, 46) <= 0; flappy_W(24, 47) <= 0; flappy_W(24, 48) <= 0; flappy_W(24, 49) <= 0; flappy_W(24, 50) <= 0; flappy_W(24, 51) <= 0; flappy_W(24, 52) <= 0; flappy_W(24, 53) <= 0; flappy_W(24, 54) <= 0; flappy_W(24, 55) <= 0; flappy_W(24, 56) <= 0; flappy_W(24, 57) <= 0; flappy_W(24, 58) <= 0; flappy_W(24, 59) <= 0; flappy_W(24, 60) <= 1; flappy_W(24, 61) <= 1; flappy_W(24, 62) <= 1; flappy_W(24, 63) <= 1; flappy_W(24, 64) <= 1; flappy_W(24, 65) <= 1; flappy_W(24, 66) <= 1; flappy_W(24, 67) <= 1; flappy_W(24, 68) <= 1; flappy_W(24, 69) <= 1; flappy_W(24, 70) <= 1; flappy_W(24, 71) <= 1; flappy_W(24, 72) <= 0; flappy_W(24, 73) <= 0; flappy_W(24, 74) <= 0; flappy_W(24, 75) <= 0; flappy_W(24, 76) <= 0; flappy_W(24, 77) <= 0; flappy_W(24, 78) <= 0; flappy_W(24, 79) <= 0; flappy_W(24, 80) <= 0; flappy_W(24, 81) <= 0; flappy_W(24, 82) <= 0; flappy_W(24, 83) <= 0; flappy_W(24, 84) <= 0; flappy_W(24, 85) <= 0; flappy_W(24, 86) <= 0; flappy_W(24, 87) <= 0; flappy_W(24, 88) <= 0; flappy_W(24, 89) <= 0; flappy_W(24, 90) <= 0; flappy_W(24, 91) <= 0; flappy_W(24, 92) <= 0; flappy_W(24, 93) <= 0; flappy_W(24, 94) <= 0; flappy_W(24, 95) <= 0; flappy_W(24, 96) <= 0; flappy_W(24, 97) <= 0; flappy_W(24, 98) <= 0; flappy_W(24, 99) <= 0; flappy_W(24, 100) <= 0; flappy_W(24, 101) <= 0; flappy_W(24, 102) <= 0; flappy_W(24, 103) <= 0; flappy_W(24, 104) <= 0; flappy_W(24, 105) <= 0; flappy_W(24, 106) <= 0; flappy_W(24, 107) <= 0; flappy_W(24, 108) <= 1; flappy_W(24, 109) <= 1; flappy_W(24, 110) <= 1; flappy_W(24, 111) <= 1; flappy_W(24, 112) <= 1; flappy_W(24, 113) <= 1; flappy_W(24, 114) <= 1; flappy_W(24, 115) <= 1; flappy_W(24, 116) <= 1; flappy_W(24, 117) <= 1; flappy_W(24, 118) <= 1; flappy_W(24, 119) <= 1; flappy_W(24, 120) <= 0; flappy_W(24, 121) <= 0; flappy_W(24, 122) <= 0; flappy_W(24, 123) <= 0; flappy_W(24, 124) <= 0; flappy_W(24, 125) <= 0; flappy_W(24, 126) <= 0; flappy_W(24, 127) <= 0; flappy_W(24, 128) <= 0; flappy_W(24, 129) <= 0; flappy_W(24, 130) <= 0; flappy_W(24, 131) <= 0; flappy_W(24, 132) <= 0; flappy_W(24, 133) <= 0; flappy_W(24, 134) <= 0; flappy_W(24, 135) <= 0; flappy_W(24, 136) <= 0; flappy_W(24, 137) <= 0; flappy_W(24, 138) <= 1; flappy_W(24, 139) <= 1; flappy_W(24, 140) <= 1; flappy_W(24, 141) <= 1; flappy_W(24, 142) <= 1; flappy_W(24, 143) <= 1; flappy_W(24, 144) <= 1; flappy_W(24, 145) <= 1; flappy_W(24, 146) <= 1; flappy_W(24, 147) <= 1; flappy_W(24, 148) <= 1; flappy_W(24, 149) <= 1; flappy_W(24, 150) <= 0; flappy_W(24, 151) <= 0; flappy_W(24, 152) <= 0; flappy_W(24, 153) <= 0; flappy_W(24, 154) <= 0; flappy_W(24, 155) <= 0; flappy_W(24, 156) <= 0; flappy_W(24, 157) <= 0; flappy_W(24, 158) <= 0; flappy_W(24, 159) <= 0; flappy_W(24, 160) <= 0; flappy_W(24, 161) <= 0; flappy_W(24, 162) <= 0; flappy_W(24, 163) <= 0; flappy_W(24, 164) <= 0; flappy_W(24, 165) <= 0; flappy_W(24, 166) <= 0; flappy_W(24, 167) <= 0; flappy_W(24, 168) <= 1; flappy_W(24, 169) <= 1; flappy_W(24, 170) <= 1; flappy_W(24, 171) <= 1; flappy_W(24, 172) <= 1; flappy_W(24, 173) <= 1; flappy_W(24, 174) <= 1; flappy_W(24, 175) <= 1; flappy_W(24, 176) <= 1; flappy_W(24, 177) <= 1; flappy_W(24, 178) <= 1; flappy_W(24, 179) <= 1; flappy_W(24, 180) <= 1; flappy_W(24, 181) <= 1; flappy_W(24, 182) <= 1; flappy_W(24, 183) <= 1; flappy_W(24, 184) <= 1; flappy_W(24, 185) <= 1; flappy_W(24, 186) <= 1; flappy_W(24, 187) <= 1; flappy_W(24, 188) <= 1; flappy_W(24, 189) <= 1; flappy_W(24, 190) <= 1; flappy_W(24, 191) <= 1; flappy_W(24, 192) <= 1; flappy_W(24, 193) <= 1; flappy_W(24, 194) <= 1; flappy_W(24, 195) <= 1; flappy_W(24, 196) <= 1; flappy_W(24, 197) <= 1; flappy_W(24, 198) <= 0; flappy_W(24, 199) <= 0; flappy_W(24, 200) <= 0; flappy_W(24, 201) <= 0; flappy_W(24, 202) <= 0; flappy_W(24, 203) <= 0; flappy_W(24, 204) <= 0; flappy_W(24, 205) <= 0; flappy_W(24, 206) <= 0; flappy_W(24, 207) <= 0; flappy_W(24, 208) <= 0; flappy_W(24, 209) <= 0; flappy_W(24, 210) <= 0; flappy_W(24, 211) <= 0; flappy_W(24, 212) <= 0; flappy_W(24, 213) <= 0; flappy_W(24, 214) <= 0; flappy_W(24, 215) <= 0; flappy_W(24, 216) <= 0; flappy_W(24, 217) <= 0; flappy_W(24, 218) <= 0; flappy_W(24, 219) <= 0; flappy_W(24, 220) <= 0; flappy_W(24, 221) <= 0; flappy_W(24, 222) <= 1; flappy_W(24, 223) <= 1; flappy_W(24, 224) <= 1; flappy_W(24, 225) <= 1; flappy_W(24, 226) <= 1; flappy_W(24, 227) <= 1; flappy_W(24, 228) <= 1; flappy_W(24, 229) <= 1; flappy_W(24, 230) <= 1; flappy_W(24, 231) <= 1; flappy_W(24, 232) <= 1; flappy_W(24, 233) <= 1; flappy_W(24, 234) <= 1; flappy_W(24, 235) <= 1; flappy_W(24, 236) <= 1; flappy_W(24, 237) <= 1; flappy_W(24, 238) <= 1; flappy_W(24, 239) <= 1; flappy_W(24, 240) <= 1; flappy_W(24, 241) <= 1; flappy_W(24, 242) <= 1; flappy_W(24, 243) <= 1; flappy_W(24, 244) <= 1; flappy_W(24, 245) <= 1; flappy_W(24, 246) <= 1; flappy_W(24, 247) <= 1; flappy_W(24, 248) <= 1; flappy_W(24, 249) <= 1; flappy_W(24, 250) <= 1; flappy_W(24, 251) <= 1; flappy_W(24, 252) <= 0; flappy_W(24, 253) <= 0; flappy_W(24, 254) <= 0; flappy_W(24, 255) <= 0; flappy_W(24, 256) <= 0; flappy_W(24, 257) <= 0; flappy_W(24, 258) <= 0; flappy_W(24, 259) <= 0; flappy_W(24, 260) <= 0; flappy_W(24, 261) <= 0; flappy_W(24, 262) <= 0; flappy_W(24, 263) <= 0; flappy_W(24, 264) <= 0; flappy_W(24, 265) <= 0; flappy_W(24, 266) <= 0; flappy_W(24, 267) <= 0; flappy_W(24, 268) <= 0; flappy_W(24, 269) <= 0; flappy_W(24, 270) <= 0; flappy_W(24, 271) <= 0; flappy_W(24, 272) <= 0; flappy_W(24, 273) <= 0; flappy_W(24, 274) <= 0; flappy_W(24, 275) <= 0; flappy_W(24, 276) <= 0; flappy_W(24, 277) <= 0; flappy_W(24, 278) <= 0; flappy_W(24, 279) <= 0; flappy_W(24, 280) <= 0; flappy_W(24, 281) <= 0; flappy_W(24, 282) <= 1; flappy_W(24, 283) <= 1; flappy_W(24, 284) <= 1; flappy_W(24, 285) <= 1; flappy_W(24, 286) <= 1; flappy_W(24, 287) <= 1; flappy_W(24, 288) <= 1; flappy_W(24, 289) <= 1; flappy_W(24, 290) <= 1; flappy_W(24, 291) <= 1; flappy_W(24, 292) <= 1; flappy_W(24, 293) <= 1; flappy_W(24, 294) <= 1; flappy_W(24, 295) <= 1; flappy_W(24, 296) <= 1; flappy_W(24, 297) <= 1; flappy_W(24, 298) <= 1; flappy_W(24, 299) <= 1; flappy_W(24, 300) <= 1; flappy_W(24, 301) <= 1; flappy_W(24, 302) <= 1; flappy_W(24, 303) <= 1; flappy_W(24, 304) <= 1; flappy_W(24, 305) <= 1; flappy_W(24, 306) <= 0; flappy_W(24, 307) <= 0; flappy_W(24, 308) <= 0; flappy_W(24, 309) <= 0; flappy_W(24, 310) <= 0; flappy_W(24, 311) <= 0; flappy_W(24, 312) <= 0; flappy_W(24, 313) <= 0; flappy_W(24, 314) <= 0; flappy_W(24, 315) <= 0; flappy_W(24, 316) <= 0; flappy_W(24, 317) <= 0; flappy_W(24, 318) <= 0; flappy_W(24, 319) <= 0; flappy_W(24, 320) <= 0; flappy_W(24, 321) <= 0; flappy_W(24, 322) <= 0; flappy_W(24, 323) <= 0; flappy_W(24, 324) <= 0; flappy_W(24, 325) <= 0; flappy_W(24, 326) <= 0; flappy_W(24, 327) <= 0; flappy_W(24, 328) <= 0; flappy_W(24, 329) <= 0; flappy_W(24, 330) <= 0; flappy_W(24, 331) <= 0; flappy_W(24, 332) <= 0; flappy_W(24, 333) <= 0; flappy_W(24, 334) <= 0; flappy_W(24, 335) <= 0; flappy_W(24, 336) <= 0; flappy_W(24, 337) <= 0; flappy_W(24, 338) <= 0; flappy_W(24, 339) <= 0; flappy_W(24, 340) <= 0; flappy_W(24, 341) <= 0; flappy_W(24, 342) <= 0; flappy_W(24, 343) <= 0; flappy_W(24, 344) <= 0; flappy_W(24, 345) <= 0; flappy_W(24, 346) <= 0; flappy_W(24, 347) <= 0; flappy_W(24, 348) <= 0; flappy_W(24, 349) <= 0; flappy_W(24, 350) <= 0; flappy_W(24, 351) <= 0; flappy_W(24, 352) <= 0; flappy_W(24, 353) <= 0; flappy_W(24, 354) <= 0; flappy_W(24, 355) <= 0; flappy_W(24, 356) <= 0; flappy_W(24, 357) <= 0; flappy_W(24, 358) <= 0; flappy_W(24, 359) <= 0; flappy_W(24, 360) <= 0; flappy_W(24, 361) <= 0; flappy_W(24, 362) <= 0; flappy_W(24, 363) <= 0; flappy_W(24, 364) <= 0; flappy_W(24, 365) <= 0; flappy_W(24, 366) <= 0; flappy_W(24, 367) <= 0; flappy_W(24, 368) <= 0; flappy_W(24, 369) <= 0; flappy_W(24, 370) <= 0; flappy_W(24, 371) <= 0; flappy_W(24, 372) <= 0; flappy_W(24, 373) <= 0; flappy_W(24, 374) <= 0; flappy_W(24, 375) <= 0; flappy_W(24, 376) <= 0; flappy_W(24, 377) <= 0; flappy_W(24, 378) <= 0; flappy_W(24, 379) <= 0; flappy_W(24, 380) <= 0; flappy_W(24, 381) <= 0; flappy_W(24, 382) <= 0; flappy_W(24, 383) <= 0; flappy_W(24, 384) <= 0; flappy_W(24, 385) <= 0; flappy_W(24, 386) <= 0; flappy_W(24, 387) <= 0; flappy_W(24, 388) <= 0; flappy_W(24, 389) <= 0; flappy_W(24, 390) <= 0; flappy_W(24, 391) <= 0; flappy_W(24, 392) <= 0; flappy_W(24, 393) <= 0; flappy_W(24, 394) <= 0; flappy_W(24, 395) <= 0; flappy_W(24, 396) <= 0; flappy_W(24, 397) <= 0; flappy_W(24, 398) <= 0; flappy_W(24, 399) <= 0; flappy_W(24, 400) <= 0; flappy_W(24, 401) <= 0; flappy_W(24, 402) <= 1; flappy_W(24, 403) <= 1; flappy_W(24, 404) <= 1; flappy_W(24, 405) <= 1; flappy_W(24, 406) <= 1; flappy_W(24, 407) <= 1; flappy_W(24, 408) <= 1; flappy_W(24, 409) <= 1; flappy_W(24, 410) <= 1; flappy_W(24, 411) <= 1; flappy_W(24, 412) <= 1; flappy_W(24, 413) <= 1; flappy_W(24, 414) <= 1; flappy_W(24, 415) <= 1; flappy_W(24, 416) <= 1; flappy_W(24, 417) <= 1; flappy_W(24, 418) <= 1; flappy_W(24, 419) <= 1; flappy_W(24, 420) <= 1; flappy_W(24, 421) <= 1; flappy_W(24, 422) <= 1; flappy_W(24, 423) <= 1; flappy_W(24, 424) <= 1; flappy_W(24, 425) <= 1; flappy_W(24, 426) <= 1; flappy_W(24, 427) <= 1; flappy_W(24, 428) <= 1; flappy_W(24, 429) <= 1; flappy_W(24, 430) <= 1; flappy_W(24, 431) <= 1; flappy_W(24, 432) <= 0; flappy_W(24, 433) <= 0; flappy_W(24, 434) <= 0; flappy_W(24, 435) <= 0; flappy_W(24, 436) <= 0; flappy_W(24, 437) <= 0; flappy_W(24, 438) <= 0; flappy_W(24, 439) <= 0; flappy_W(24, 440) <= 0; flappy_W(24, 441) <= 0; flappy_W(24, 442) <= 0; flappy_W(24, 443) <= 0; flappy_W(24, 444) <= 0; flappy_W(24, 445) <= 0; flappy_W(24, 446) <= 0; flappy_W(24, 447) <= 0; flappy_W(24, 448) <= 0; flappy_W(24, 449) <= 0; flappy_W(24, 450) <= 0; flappy_W(24, 451) <= 0; flappy_W(24, 452) <= 0; flappy_W(24, 453) <= 0; flappy_W(24, 454) <= 0; flappy_W(24, 455) <= 0; flappy_W(24, 456) <= 0; flappy_W(24, 457) <= 0; flappy_W(24, 458) <= 0; flappy_W(24, 459) <= 0; flappy_W(24, 460) <= 0; flappy_W(24, 461) <= 0; flappy_W(24, 462) <= 0; flappy_W(24, 463) <= 0; flappy_W(24, 464) <= 0; flappy_W(24, 465) <= 0; flappy_W(24, 466) <= 0; flappy_W(24, 467) <= 0; flappy_W(24, 468) <= 1; flappy_W(24, 469) <= 1; flappy_W(24, 470) <= 1; flappy_W(24, 471) <= 1; flappy_W(24, 472) <= 1; flappy_W(24, 473) <= 1; flappy_W(24, 474) <= 1; flappy_W(24, 475) <= 1; flappy_W(24, 476) <= 1; flappy_W(24, 477) <= 1; flappy_W(24, 478) <= 1; flappy_W(24, 479) <= 1; flappy_W(24, 480) <= 0; flappy_W(24, 481) <= 0; flappy_W(24, 482) <= 0; flappy_W(24, 483) <= 0; flappy_W(24, 484) <= 0; flappy_W(24, 485) <= 0; flappy_W(24, 486) <= 0; flappy_W(24, 487) <= 0; flappy_W(24, 488) <= 0; flappy_W(24, 489) <= 0; flappy_W(24, 490) <= 0; flappy_W(24, 491) <= 0; flappy_W(24, 492) <= 0; flappy_W(24, 493) <= 0; flappy_W(24, 494) <= 0; flappy_W(24, 495) <= 0; flappy_W(24, 496) <= 0; flappy_W(24, 497) <= 0; flappy_W(24, 498) <= 0; flappy_W(24, 499) <= 0; flappy_W(24, 500) <= 0; flappy_W(24, 501) <= 0; flappy_W(24, 502) <= 0; flappy_W(24, 503) <= 0; flappy_W(24, 504) <= 0; flappy_W(24, 505) <= 0; flappy_W(24, 506) <= 0; flappy_W(24, 507) <= 0; flappy_W(24, 508) <= 0; flappy_W(24, 509) <= 0; flappy_W(24, 510) <= 1; flappy_W(24, 511) <= 1; flappy_W(24, 512) <= 1; flappy_W(24, 513) <= 1; flappy_W(24, 514) <= 1; flappy_W(24, 515) <= 1; flappy_W(24, 516) <= 1; flappy_W(24, 517) <= 1; flappy_W(24, 518) <= 1; flappy_W(24, 519) <= 1; flappy_W(24, 520) <= 1; flappy_W(24, 521) <= 1; flappy_W(24, 522) <= 1; flappy_W(24, 523) <= 1; flappy_W(24, 524) <= 1; flappy_W(24, 525) <= 1; flappy_W(24, 526) <= 1; flappy_W(24, 527) <= 1; flappy_W(24, 528) <= 1; flappy_W(24, 529) <= 1; flappy_W(24, 530) <= 1; flappy_W(24, 531) <= 1; flappy_W(24, 532) <= 1; flappy_W(24, 533) <= 1; flappy_W(24, 534) <= 1; flappy_W(24, 535) <= 1; flappy_W(24, 536) <= 1; flappy_W(24, 537) <= 1; flappy_W(24, 538) <= 1; flappy_W(24, 539) <= 1; flappy_W(24, 540) <= 0; flappy_W(24, 541) <= 0; flappy_W(24, 542) <= 0; flappy_W(24, 543) <= 0; flappy_W(24, 544) <= 0; flappy_W(24, 545) <= 0; flappy_W(24, 546) <= 0; flappy_W(24, 547) <= 0; flappy_W(24, 548) <= 0; flappy_W(24, 549) <= 0; flappy_W(24, 550) <= 0; flappy_W(24, 551) <= 0; flappy_W(24, 552) <= 0; flappy_W(24, 553) <= 0; flappy_W(24, 554) <= 0; flappy_W(24, 555) <= 0; flappy_W(24, 556) <= 0; flappy_W(24, 557) <= 0; flappy_W(24, 558) <= 0; flappy_W(24, 559) <= 0; flappy_W(24, 560) <= 0; flappy_W(24, 561) <= 0; flappy_W(24, 562) <= 0; flappy_W(24, 563) <= 0; flappy_W(24, 564) <= 1; flappy_W(24, 565) <= 1; flappy_W(24, 566) <= 1; flappy_W(24, 567) <= 1; flappy_W(24, 568) <= 1; flappy_W(24, 569) <= 1; flappy_W(24, 570) <= 1; flappy_W(24, 571) <= 1; flappy_W(24, 572) <= 1; flappy_W(24, 573) <= 1; flappy_W(24, 574) <= 1; flappy_W(24, 575) <= 1; flappy_W(24, 576) <= 0; flappy_W(24, 577) <= 0; flappy_W(24, 578) <= 0; flappy_W(24, 579) <= 0; flappy_W(24, 580) <= 0; flappy_W(24, 581) <= 0; flappy_W(24, 582) <= 0; flappy_W(24, 583) <= 0; flappy_W(24, 584) <= 0; flappy_W(24, 585) <= 0; flappy_W(24, 586) <= 0; flappy_W(24, 587) <= 0; flappy_W(24, 588) <= 1; flappy_W(24, 589) <= 1; flappy_W(24, 590) <= 1; flappy_W(24, 591) <= 1; flappy_W(24, 592) <= 1; flappy_W(24, 593) <= 1; 
flappy_W(25, 0) <= 0; flappy_W(25, 1) <= 0; flappy_W(25, 2) <= 0; flappy_W(25, 3) <= 0; flappy_W(25, 4) <= 0; flappy_W(25, 5) <= 0; flappy_W(25, 6) <= 1; flappy_W(25, 7) <= 1; flappy_W(25, 8) <= 1; flappy_W(25, 9) <= 1; flappy_W(25, 10) <= 1; flappy_W(25, 11) <= 1; flappy_W(25, 12) <= 1; flappy_W(25, 13) <= 1; flappy_W(25, 14) <= 1; flappy_W(25, 15) <= 1; flappy_W(25, 16) <= 1; flappy_W(25, 17) <= 1; flappy_W(25, 18) <= 1; flappy_W(25, 19) <= 1; flappy_W(25, 20) <= 1; flappy_W(25, 21) <= 1; flappy_W(25, 22) <= 1; flappy_W(25, 23) <= 1; flappy_W(25, 24) <= 1; flappy_W(25, 25) <= 1; flappy_W(25, 26) <= 1; flappy_W(25, 27) <= 1; flappy_W(25, 28) <= 1; flappy_W(25, 29) <= 1; flappy_W(25, 30) <= 0; flappy_W(25, 31) <= 0; flappy_W(25, 32) <= 0; flappy_W(25, 33) <= 0; flappy_W(25, 34) <= 0; flappy_W(25, 35) <= 0; flappy_W(25, 36) <= 0; flappy_W(25, 37) <= 0; flappy_W(25, 38) <= 0; flappy_W(25, 39) <= 0; flappy_W(25, 40) <= 0; flappy_W(25, 41) <= 0; flappy_W(25, 42) <= 0; flappy_W(25, 43) <= 0; flappy_W(25, 44) <= 0; flappy_W(25, 45) <= 0; flappy_W(25, 46) <= 0; flappy_W(25, 47) <= 0; flappy_W(25, 48) <= 0; flappy_W(25, 49) <= 0; flappy_W(25, 50) <= 0; flappy_W(25, 51) <= 0; flappy_W(25, 52) <= 0; flappy_W(25, 53) <= 0; flappy_W(25, 54) <= 0; flappy_W(25, 55) <= 0; flappy_W(25, 56) <= 0; flappy_W(25, 57) <= 0; flappy_W(25, 58) <= 0; flappy_W(25, 59) <= 0; flappy_W(25, 60) <= 1; flappy_W(25, 61) <= 1; flappy_W(25, 62) <= 1; flappy_W(25, 63) <= 1; flappy_W(25, 64) <= 1; flappy_W(25, 65) <= 1; flappy_W(25, 66) <= 1; flappy_W(25, 67) <= 1; flappy_W(25, 68) <= 1; flappy_W(25, 69) <= 1; flappy_W(25, 70) <= 1; flappy_W(25, 71) <= 1; flappy_W(25, 72) <= 0; flappy_W(25, 73) <= 0; flappy_W(25, 74) <= 0; flappy_W(25, 75) <= 0; flappy_W(25, 76) <= 0; flappy_W(25, 77) <= 0; flappy_W(25, 78) <= 0; flappy_W(25, 79) <= 0; flappy_W(25, 80) <= 0; flappy_W(25, 81) <= 0; flappy_W(25, 82) <= 0; flappy_W(25, 83) <= 0; flappy_W(25, 84) <= 0; flappy_W(25, 85) <= 0; flappy_W(25, 86) <= 0; flappy_W(25, 87) <= 0; flappy_W(25, 88) <= 0; flappy_W(25, 89) <= 0; flappy_W(25, 90) <= 0; flappy_W(25, 91) <= 0; flappy_W(25, 92) <= 0; flappy_W(25, 93) <= 0; flappy_W(25, 94) <= 0; flappy_W(25, 95) <= 0; flappy_W(25, 96) <= 0; flappy_W(25, 97) <= 0; flappy_W(25, 98) <= 0; flappy_W(25, 99) <= 0; flappy_W(25, 100) <= 0; flappy_W(25, 101) <= 0; flappy_W(25, 102) <= 0; flappy_W(25, 103) <= 0; flappy_W(25, 104) <= 0; flappy_W(25, 105) <= 0; flappy_W(25, 106) <= 0; flappy_W(25, 107) <= 0; flappy_W(25, 108) <= 1; flappy_W(25, 109) <= 1; flappy_W(25, 110) <= 1; flappy_W(25, 111) <= 1; flappy_W(25, 112) <= 1; flappy_W(25, 113) <= 1; flappy_W(25, 114) <= 1; flappy_W(25, 115) <= 1; flappy_W(25, 116) <= 1; flappy_W(25, 117) <= 1; flappy_W(25, 118) <= 1; flappy_W(25, 119) <= 1; flappy_W(25, 120) <= 0; flappy_W(25, 121) <= 0; flappy_W(25, 122) <= 0; flappy_W(25, 123) <= 0; flappy_W(25, 124) <= 0; flappy_W(25, 125) <= 0; flappy_W(25, 126) <= 0; flappy_W(25, 127) <= 0; flappy_W(25, 128) <= 0; flappy_W(25, 129) <= 0; flappy_W(25, 130) <= 0; flappy_W(25, 131) <= 0; flappy_W(25, 132) <= 0; flappy_W(25, 133) <= 0; flappy_W(25, 134) <= 0; flappy_W(25, 135) <= 0; flappy_W(25, 136) <= 0; flappy_W(25, 137) <= 0; flappy_W(25, 138) <= 1; flappy_W(25, 139) <= 1; flappy_W(25, 140) <= 1; flappy_W(25, 141) <= 1; flappy_W(25, 142) <= 1; flappy_W(25, 143) <= 1; flappy_W(25, 144) <= 1; flappy_W(25, 145) <= 1; flappy_W(25, 146) <= 1; flappy_W(25, 147) <= 1; flappy_W(25, 148) <= 1; flappy_W(25, 149) <= 1; flappy_W(25, 150) <= 0; flappy_W(25, 151) <= 0; flappy_W(25, 152) <= 0; flappy_W(25, 153) <= 0; flappy_W(25, 154) <= 0; flappy_W(25, 155) <= 0; flappy_W(25, 156) <= 0; flappy_W(25, 157) <= 0; flappy_W(25, 158) <= 0; flappy_W(25, 159) <= 0; flappy_W(25, 160) <= 0; flappy_W(25, 161) <= 0; flappy_W(25, 162) <= 0; flappy_W(25, 163) <= 0; flappy_W(25, 164) <= 0; flappy_W(25, 165) <= 0; flappy_W(25, 166) <= 0; flappy_W(25, 167) <= 0; flappy_W(25, 168) <= 1; flappy_W(25, 169) <= 1; flappy_W(25, 170) <= 1; flappy_W(25, 171) <= 1; flappy_W(25, 172) <= 1; flappy_W(25, 173) <= 1; flappy_W(25, 174) <= 1; flappy_W(25, 175) <= 1; flappy_W(25, 176) <= 1; flappy_W(25, 177) <= 1; flappy_W(25, 178) <= 1; flappy_W(25, 179) <= 1; flappy_W(25, 180) <= 1; flappy_W(25, 181) <= 1; flappy_W(25, 182) <= 1; flappy_W(25, 183) <= 1; flappy_W(25, 184) <= 1; flappy_W(25, 185) <= 1; flappy_W(25, 186) <= 1; flappy_W(25, 187) <= 1; flappy_W(25, 188) <= 1; flappy_W(25, 189) <= 1; flappy_W(25, 190) <= 1; flappy_W(25, 191) <= 1; flappy_W(25, 192) <= 1; flappy_W(25, 193) <= 1; flappy_W(25, 194) <= 1; flappy_W(25, 195) <= 1; flappy_W(25, 196) <= 1; flappy_W(25, 197) <= 1; flappy_W(25, 198) <= 0; flappy_W(25, 199) <= 0; flappy_W(25, 200) <= 0; flappy_W(25, 201) <= 0; flappy_W(25, 202) <= 0; flappy_W(25, 203) <= 0; flappy_W(25, 204) <= 0; flappy_W(25, 205) <= 0; flappy_W(25, 206) <= 0; flappy_W(25, 207) <= 0; flappy_W(25, 208) <= 0; flappy_W(25, 209) <= 0; flappy_W(25, 210) <= 0; flappy_W(25, 211) <= 0; flappy_W(25, 212) <= 0; flappy_W(25, 213) <= 0; flappy_W(25, 214) <= 0; flappy_W(25, 215) <= 0; flappy_W(25, 216) <= 0; flappy_W(25, 217) <= 0; flappy_W(25, 218) <= 0; flappy_W(25, 219) <= 0; flappy_W(25, 220) <= 0; flappy_W(25, 221) <= 0; flappy_W(25, 222) <= 1; flappy_W(25, 223) <= 1; flappy_W(25, 224) <= 1; flappy_W(25, 225) <= 1; flappy_W(25, 226) <= 1; flappy_W(25, 227) <= 1; flappy_W(25, 228) <= 1; flappy_W(25, 229) <= 1; flappy_W(25, 230) <= 1; flappy_W(25, 231) <= 1; flappy_W(25, 232) <= 1; flappy_W(25, 233) <= 1; flappy_W(25, 234) <= 1; flappy_W(25, 235) <= 1; flappy_W(25, 236) <= 1; flappy_W(25, 237) <= 1; flappy_W(25, 238) <= 1; flappy_W(25, 239) <= 1; flappy_W(25, 240) <= 1; flappy_W(25, 241) <= 1; flappy_W(25, 242) <= 1; flappy_W(25, 243) <= 1; flappy_W(25, 244) <= 1; flappy_W(25, 245) <= 1; flappy_W(25, 246) <= 1; flappy_W(25, 247) <= 1; flappy_W(25, 248) <= 1; flappy_W(25, 249) <= 1; flappy_W(25, 250) <= 1; flappy_W(25, 251) <= 1; flappy_W(25, 252) <= 0; flappy_W(25, 253) <= 0; flappy_W(25, 254) <= 0; flappy_W(25, 255) <= 0; flappy_W(25, 256) <= 0; flappy_W(25, 257) <= 0; flappy_W(25, 258) <= 0; flappy_W(25, 259) <= 0; flappy_W(25, 260) <= 0; flappy_W(25, 261) <= 0; flappy_W(25, 262) <= 0; flappy_W(25, 263) <= 0; flappy_W(25, 264) <= 0; flappy_W(25, 265) <= 0; flappy_W(25, 266) <= 0; flappy_W(25, 267) <= 0; flappy_W(25, 268) <= 0; flappy_W(25, 269) <= 0; flappy_W(25, 270) <= 0; flappy_W(25, 271) <= 0; flappy_W(25, 272) <= 0; flappy_W(25, 273) <= 0; flappy_W(25, 274) <= 0; flappy_W(25, 275) <= 0; flappy_W(25, 276) <= 0; flappy_W(25, 277) <= 0; flappy_W(25, 278) <= 0; flappy_W(25, 279) <= 0; flappy_W(25, 280) <= 0; flappy_W(25, 281) <= 0; flappy_W(25, 282) <= 1; flappy_W(25, 283) <= 1; flappy_W(25, 284) <= 1; flappy_W(25, 285) <= 1; flappy_W(25, 286) <= 1; flappy_W(25, 287) <= 1; flappy_W(25, 288) <= 1; flappy_W(25, 289) <= 1; flappy_W(25, 290) <= 1; flappy_W(25, 291) <= 1; flappy_W(25, 292) <= 1; flappy_W(25, 293) <= 1; flappy_W(25, 294) <= 1; flappy_W(25, 295) <= 1; flappy_W(25, 296) <= 1; flappy_W(25, 297) <= 1; flappy_W(25, 298) <= 1; flappy_W(25, 299) <= 1; flappy_W(25, 300) <= 1; flappy_W(25, 301) <= 1; flappy_W(25, 302) <= 1; flappy_W(25, 303) <= 1; flappy_W(25, 304) <= 1; flappy_W(25, 305) <= 1; flappy_W(25, 306) <= 0; flappy_W(25, 307) <= 0; flappy_W(25, 308) <= 0; flappy_W(25, 309) <= 0; flappy_W(25, 310) <= 0; flappy_W(25, 311) <= 0; flappy_W(25, 312) <= 0; flappy_W(25, 313) <= 0; flappy_W(25, 314) <= 0; flappy_W(25, 315) <= 0; flappy_W(25, 316) <= 0; flappy_W(25, 317) <= 0; flappy_W(25, 318) <= 0; flappy_W(25, 319) <= 0; flappy_W(25, 320) <= 0; flappy_W(25, 321) <= 0; flappy_W(25, 322) <= 0; flappy_W(25, 323) <= 0; flappy_W(25, 324) <= 0; flappy_W(25, 325) <= 0; flappy_W(25, 326) <= 0; flappy_W(25, 327) <= 0; flappy_W(25, 328) <= 0; flappy_W(25, 329) <= 0; flappy_W(25, 330) <= 0; flappy_W(25, 331) <= 0; flappy_W(25, 332) <= 0; flappy_W(25, 333) <= 0; flappy_W(25, 334) <= 0; flappy_W(25, 335) <= 0; flappy_W(25, 336) <= 0; flappy_W(25, 337) <= 0; flappy_W(25, 338) <= 0; flappy_W(25, 339) <= 0; flappy_W(25, 340) <= 0; flappy_W(25, 341) <= 0; flappy_W(25, 342) <= 0; flappy_W(25, 343) <= 0; flappy_W(25, 344) <= 0; flappy_W(25, 345) <= 0; flappy_W(25, 346) <= 0; flappy_W(25, 347) <= 0; flappy_W(25, 348) <= 0; flappy_W(25, 349) <= 0; flappy_W(25, 350) <= 0; flappy_W(25, 351) <= 0; flappy_W(25, 352) <= 0; flappy_W(25, 353) <= 0; flappy_W(25, 354) <= 0; flappy_W(25, 355) <= 0; flappy_W(25, 356) <= 0; flappy_W(25, 357) <= 0; flappy_W(25, 358) <= 0; flappy_W(25, 359) <= 0; flappy_W(25, 360) <= 0; flappy_W(25, 361) <= 0; flappy_W(25, 362) <= 0; flappy_W(25, 363) <= 0; flappy_W(25, 364) <= 0; flappy_W(25, 365) <= 0; flappy_W(25, 366) <= 0; flappy_W(25, 367) <= 0; flappy_W(25, 368) <= 0; flappy_W(25, 369) <= 0; flappy_W(25, 370) <= 0; flappy_W(25, 371) <= 0; flappy_W(25, 372) <= 0; flappy_W(25, 373) <= 0; flappy_W(25, 374) <= 0; flappy_W(25, 375) <= 0; flappy_W(25, 376) <= 0; flappy_W(25, 377) <= 0; flappy_W(25, 378) <= 0; flappy_W(25, 379) <= 0; flappy_W(25, 380) <= 0; flappy_W(25, 381) <= 0; flappy_W(25, 382) <= 0; flappy_W(25, 383) <= 0; flappy_W(25, 384) <= 0; flappy_W(25, 385) <= 0; flappy_W(25, 386) <= 0; flappy_W(25, 387) <= 0; flappy_W(25, 388) <= 0; flappy_W(25, 389) <= 0; flappy_W(25, 390) <= 0; flappy_W(25, 391) <= 0; flappy_W(25, 392) <= 0; flappy_W(25, 393) <= 0; flappy_W(25, 394) <= 0; flappy_W(25, 395) <= 0; flappy_W(25, 396) <= 0; flappy_W(25, 397) <= 0; flappy_W(25, 398) <= 0; flappy_W(25, 399) <= 0; flappy_W(25, 400) <= 0; flappy_W(25, 401) <= 0; flappy_W(25, 402) <= 1; flappy_W(25, 403) <= 1; flappy_W(25, 404) <= 1; flappy_W(25, 405) <= 1; flappy_W(25, 406) <= 1; flappy_W(25, 407) <= 1; flappy_W(25, 408) <= 1; flappy_W(25, 409) <= 1; flappy_W(25, 410) <= 1; flappy_W(25, 411) <= 1; flappy_W(25, 412) <= 1; flappy_W(25, 413) <= 1; flappy_W(25, 414) <= 1; flappy_W(25, 415) <= 1; flappy_W(25, 416) <= 1; flappy_W(25, 417) <= 1; flappy_W(25, 418) <= 1; flappy_W(25, 419) <= 1; flappy_W(25, 420) <= 1; flappy_W(25, 421) <= 1; flappy_W(25, 422) <= 1; flappy_W(25, 423) <= 1; flappy_W(25, 424) <= 1; flappy_W(25, 425) <= 1; flappy_W(25, 426) <= 1; flappy_W(25, 427) <= 1; flappy_W(25, 428) <= 1; flappy_W(25, 429) <= 1; flappy_W(25, 430) <= 1; flappy_W(25, 431) <= 1; flappy_W(25, 432) <= 0; flappy_W(25, 433) <= 0; flappy_W(25, 434) <= 0; flappy_W(25, 435) <= 0; flappy_W(25, 436) <= 0; flappy_W(25, 437) <= 0; flappy_W(25, 438) <= 0; flappy_W(25, 439) <= 0; flappy_W(25, 440) <= 0; flappy_W(25, 441) <= 0; flappy_W(25, 442) <= 0; flappy_W(25, 443) <= 0; flappy_W(25, 444) <= 0; flappy_W(25, 445) <= 0; flappy_W(25, 446) <= 0; flappy_W(25, 447) <= 0; flappy_W(25, 448) <= 0; flappy_W(25, 449) <= 0; flappy_W(25, 450) <= 0; flappy_W(25, 451) <= 0; flappy_W(25, 452) <= 0; flappy_W(25, 453) <= 0; flappy_W(25, 454) <= 0; flappy_W(25, 455) <= 0; flappy_W(25, 456) <= 0; flappy_W(25, 457) <= 0; flappy_W(25, 458) <= 0; flappy_W(25, 459) <= 0; flappy_W(25, 460) <= 0; flappy_W(25, 461) <= 0; flappy_W(25, 462) <= 0; flappy_W(25, 463) <= 0; flappy_W(25, 464) <= 0; flappy_W(25, 465) <= 0; flappy_W(25, 466) <= 0; flappy_W(25, 467) <= 0; flappy_W(25, 468) <= 1; flappy_W(25, 469) <= 1; flappy_W(25, 470) <= 1; flappy_W(25, 471) <= 1; flappy_W(25, 472) <= 1; flappy_W(25, 473) <= 1; flappy_W(25, 474) <= 1; flappy_W(25, 475) <= 1; flappy_W(25, 476) <= 1; flappy_W(25, 477) <= 1; flappy_W(25, 478) <= 1; flappy_W(25, 479) <= 1; flappy_W(25, 480) <= 0; flappy_W(25, 481) <= 0; flappy_W(25, 482) <= 0; flappy_W(25, 483) <= 0; flappy_W(25, 484) <= 0; flappy_W(25, 485) <= 0; flappy_W(25, 486) <= 0; flappy_W(25, 487) <= 0; flappy_W(25, 488) <= 0; flappy_W(25, 489) <= 0; flappy_W(25, 490) <= 0; flappy_W(25, 491) <= 0; flappy_W(25, 492) <= 0; flappy_W(25, 493) <= 0; flappy_W(25, 494) <= 0; flappy_W(25, 495) <= 0; flappy_W(25, 496) <= 0; flappy_W(25, 497) <= 0; flappy_W(25, 498) <= 0; flappy_W(25, 499) <= 0; flappy_W(25, 500) <= 0; flappy_W(25, 501) <= 0; flappy_W(25, 502) <= 0; flappy_W(25, 503) <= 0; flappy_W(25, 504) <= 0; flappy_W(25, 505) <= 0; flappy_W(25, 506) <= 0; flappy_W(25, 507) <= 0; flappy_W(25, 508) <= 0; flappy_W(25, 509) <= 0; flappy_W(25, 510) <= 1; flappy_W(25, 511) <= 1; flappy_W(25, 512) <= 1; flappy_W(25, 513) <= 1; flappy_W(25, 514) <= 1; flappy_W(25, 515) <= 1; flappy_W(25, 516) <= 1; flappy_W(25, 517) <= 1; flappy_W(25, 518) <= 1; flappy_W(25, 519) <= 1; flappy_W(25, 520) <= 1; flappy_W(25, 521) <= 1; flappy_W(25, 522) <= 1; flappy_W(25, 523) <= 1; flappy_W(25, 524) <= 1; flappy_W(25, 525) <= 1; flappy_W(25, 526) <= 1; flappy_W(25, 527) <= 1; flappy_W(25, 528) <= 1; flappy_W(25, 529) <= 1; flappy_W(25, 530) <= 1; flappy_W(25, 531) <= 1; flappy_W(25, 532) <= 1; flappy_W(25, 533) <= 1; flappy_W(25, 534) <= 1; flappy_W(25, 535) <= 1; flappy_W(25, 536) <= 1; flappy_W(25, 537) <= 1; flappy_W(25, 538) <= 1; flappy_W(25, 539) <= 1; flappy_W(25, 540) <= 0; flappy_W(25, 541) <= 0; flappy_W(25, 542) <= 0; flappy_W(25, 543) <= 0; flappy_W(25, 544) <= 0; flappy_W(25, 545) <= 0; flappy_W(25, 546) <= 0; flappy_W(25, 547) <= 0; flappy_W(25, 548) <= 0; flappy_W(25, 549) <= 0; flappy_W(25, 550) <= 0; flappy_W(25, 551) <= 0; flappy_W(25, 552) <= 0; flappy_W(25, 553) <= 0; flappy_W(25, 554) <= 0; flappy_W(25, 555) <= 0; flappy_W(25, 556) <= 0; flappy_W(25, 557) <= 0; flappy_W(25, 558) <= 0; flappy_W(25, 559) <= 0; flappy_W(25, 560) <= 0; flappy_W(25, 561) <= 0; flappy_W(25, 562) <= 0; flappy_W(25, 563) <= 0; flappy_W(25, 564) <= 1; flappy_W(25, 565) <= 1; flappy_W(25, 566) <= 1; flappy_W(25, 567) <= 1; flappy_W(25, 568) <= 1; flappy_W(25, 569) <= 1; flappy_W(25, 570) <= 1; flappy_W(25, 571) <= 1; flappy_W(25, 572) <= 1; flappy_W(25, 573) <= 1; flappy_W(25, 574) <= 1; flappy_W(25, 575) <= 1; flappy_W(25, 576) <= 0; flappy_W(25, 577) <= 0; flappy_W(25, 578) <= 0; flappy_W(25, 579) <= 0; flappy_W(25, 580) <= 0; flappy_W(25, 581) <= 0; flappy_W(25, 582) <= 0; flappy_W(25, 583) <= 0; flappy_W(25, 584) <= 0; flappy_W(25, 585) <= 0; flappy_W(25, 586) <= 0; flappy_W(25, 587) <= 0; flappy_W(25, 588) <= 1; flappy_W(25, 589) <= 1; flappy_W(25, 590) <= 1; flappy_W(25, 591) <= 1; flappy_W(25, 592) <= 1; flappy_W(25, 593) <= 1; 
flappy_W(26, 0) <= 0; flappy_W(26, 1) <= 0; flappy_W(26, 2) <= 0; flappy_W(26, 3) <= 0; flappy_W(26, 4) <= 0; flappy_W(26, 5) <= 0; flappy_W(26, 6) <= 1; flappy_W(26, 7) <= 1; flappy_W(26, 8) <= 1; flappy_W(26, 9) <= 1; flappy_W(26, 10) <= 1; flappy_W(26, 11) <= 1; flappy_W(26, 12) <= 1; flappy_W(26, 13) <= 1; flappy_W(26, 14) <= 1; flappy_W(26, 15) <= 1; flappy_W(26, 16) <= 1; flappy_W(26, 17) <= 1; flappy_W(26, 18) <= 1; flappy_W(26, 19) <= 1; flappy_W(26, 20) <= 1; flappy_W(26, 21) <= 1; flappy_W(26, 22) <= 1; flappy_W(26, 23) <= 1; flappy_W(26, 24) <= 1; flappy_W(26, 25) <= 1; flappy_W(26, 26) <= 1; flappy_W(26, 27) <= 1; flappy_W(26, 28) <= 1; flappy_W(26, 29) <= 1; flappy_W(26, 30) <= 0; flappy_W(26, 31) <= 0; flappy_W(26, 32) <= 0; flappy_W(26, 33) <= 0; flappy_W(26, 34) <= 0; flappy_W(26, 35) <= 0; flappy_W(26, 36) <= 0; flappy_W(26, 37) <= 0; flappy_W(26, 38) <= 0; flappy_W(26, 39) <= 0; flappy_W(26, 40) <= 0; flappy_W(26, 41) <= 0; flappy_W(26, 42) <= 0; flappy_W(26, 43) <= 0; flappy_W(26, 44) <= 0; flappy_W(26, 45) <= 0; flappy_W(26, 46) <= 0; flappy_W(26, 47) <= 0; flappy_W(26, 48) <= 0; flappy_W(26, 49) <= 0; flappy_W(26, 50) <= 0; flappy_W(26, 51) <= 0; flappy_W(26, 52) <= 0; flappy_W(26, 53) <= 0; flappy_W(26, 54) <= 0; flappy_W(26, 55) <= 0; flappy_W(26, 56) <= 0; flappy_W(26, 57) <= 0; flappy_W(26, 58) <= 0; flappy_W(26, 59) <= 0; flappy_W(26, 60) <= 1; flappy_W(26, 61) <= 1; flappy_W(26, 62) <= 1; flappy_W(26, 63) <= 1; flappy_W(26, 64) <= 1; flappy_W(26, 65) <= 1; flappy_W(26, 66) <= 1; flappy_W(26, 67) <= 1; flappy_W(26, 68) <= 1; flappy_W(26, 69) <= 1; flappy_W(26, 70) <= 1; flappy_W(26, 71) <= 1; flappy_W(26, 72) <= 0; flappy_W(26, 73) <= 0; flappy_W(26, 74) <= 0; flappy_W(26, 75) <= 0; flappy_W(26, 76) <= 0; flappy_W(26, 77) <= 0; flappy_W(26, 78) <= 0; flappy_W(26, 79) <= 0; flappy_W(26, 80) <= 0; flappy_W(26, 81) <= 0; flappy_W(26, 82) <= 0; flappy_W(26, 83) <= 0; flappy_W(26, 84) <= 0; flappy_W(26, 85) <= 0; flappy_W(26, 86) <= 0; flappy_W(26, 87) <= 0; flappy_W(26, 88) <= 0; flappy_W(26, 89) <= 0; flappy_W(26, 90) <= 0; flappy_W(26, 91) <= 0; flappy_W(26, 92) <= 0; flappy_W(26, 93) <= 0; flappy_W(26, 94) <= 0; flappy_W(26, 95) <= 0; flappy_W(26, 96) <= 0; flappy_W(26, 97) <= 0; flappy_W(26, 98) <= 0; flappy_W(26, 99) <= 0; flappy_W(26, 100) <= 0; flappy_W(26, 101) <= 0; flappy_W(26, 102) <= 0; flappy_W(26, 103) <= 0; flappy_W(26, 104) <= 0; flappy_W(26, 105) <= 0; flappy_W(26, 106) <= 0; flappy_W(26, 107) <= 0; flappy_W(26, 108) <= 1; flappy_W(26, 109) <= 1; flappy_W(26, 110) <= 1; flappy_W(26, 111) <= 1; flappy_W(26, 112) <= 1; flappy_W(26, 113) <= 1; flappy_W(26, 114) <= 1; flappy_W(26, 115) <= 1; flappy_W(26, 116) <= 1; flappy_W(26, 117) <= 1; flappy_W(26, 118) <= 1; flappy_W(26, 119) <= 1; flappy_W(26, 120) <= 0; flappy_W(26, 121) <= 0; flappy_W(26, 122) <= 0; flappy_W(26, 123) <= 0; flappy_W(26, 124) <= 0; flappy_W(26, 125) <= 0; flappy_W(26, 126) <= 0; flappy_W(26, 127) <= 0; flappy_W(26, 128) <= 0; flappy_W(26, 129) <= 0; flappy_W(26, 130) <= 0; flappy_W(26, 131) <= 0; flappy_W(26, 132) <= 0; flappy_W(26, 133) <= 0; flappy_W(26, 134) <= 0; flappy_W(26, 135) <= 0; flappy_W(26, 136) <= 0; flappy_W(26, 137) <= 0; flappy_W(26, 138) <= 1; flappy_W(26, 139) <= 1; flappy_W(26, 140) <= 1; flappy_W(26, 141) <= 1; flappy_W(26, 142) <= 1; flappy_W(26, 143) <= 1; flappy_W(26, 144) <= 1; flappy_W(26, 145) <= 1; flappy_W(26, 146) <= 1; flappy_W(26, 147) <= 1; flappy_W(26, 148) <= 1; flappy_W(26, 149) <= 1; flappy_W(26, 150) <= 0; flappy_W(26, 151) <= 0; flappy_W(26, 152) <= 0; flappy_W(26, 153) <= 0; flappy_W(26, 154) <= 0; flappy_W(26, 155) <= 0; flappy_W(26, 156) <= 0; flappy_W(26, 157) <= 0; flappy_W(26, 158) <= 0; flappy_W(26, 159) <= 0; flappy_W(26, 160) <= 0; flappy_W(26, 161) <= 0; flappy_W(26, 162) <= 0; flappy_W(26, 163) <= 0; flappy_W(26, 164) <= 0; flappy_W(26, 165) <= 0; flappy_W(26, 166) <= 0; flappy_W(26, 167) <= 0; flappy_W(26, 168) <= 1; flappy_W(26, 169) <= 1; flappy_W(26, 170) <= 1; flappy_W(26, 171) <= 1; flappy_W(26, 172) <= 1; flappy_W(26, 173) <= 1; flappy_W(26, 174) <= 1; flappy_W(26, 175) <= 1; flappy_W(26, 176) <= 1; flappy_W(26, 177) <= 1; flappy_W(26, 178) <= 1; flappy_W(26, 179) <= 1; flappy_W(26, 180) <= 1; flappy_W(26, 181) <= 1; flappy_W(26, 182) <= 1; flappy_W(26, 183) <= 1; flappy_W(26, 184) <= 1; flappy_W(26, 185) <= 1; flappy_W(26, 186) <= 1; flappy_W(26, 187) <= 1; flappy_W(26, 188) <= 1; flappy_W(26, 189) <= 1; flappy_W(26, 190) <= 1; flappy_W(26, 191) <= 1; flappy_W(26, 192) <= 1; flappy_W(26, 193) <= 1; flappy_W(26, 194) <= 1; flappy_W(26, 195) <= 1; flappy_W(26, 196) <= 1; flappy_W(26, 197) <= 1; flappy_W(26, 198) <= 0; flappy_W(26, 199) <= 0; flappy_W(26, 200) <= 0; flappy_W(26, 201) <= 0; flappy_W(26, 202) <= 0; flappy_W(26, 203) <= 0; flappy_W(26, 204) <= 0; flappy_W(26, 205) <= 0; flappy_W(26, 206) <= 0; flappy_W(26, 207) <= 0; flappy_W(26, 208) <= 0; flappy_W(26, 209) <= 0; flappy_W(26, 210) <= 0; flappy_W(26, 211) <= 0; flappy_W(26, 212) <= 0; flappy_W(26, 213) <= 0; flappy_W(26, 214) <= 0; flappy_W(26, 215) <= 0; flappy_W(26, 216) <= 0; flappy_W(26, 217) <= 0; flappy_W(26, 218) <= 0; flappy_W(26, 219) <= 0; flappy_W(26, 220) <= 0; flappy_W(26, 221) <= 0; flappy_W(26, 222) <= 1; flappy_W(26, 223) <= 1; flappy_W(26, 224) <= 1; flappy_W(26, 225) <= 1; flappy_W(26, 226) <= 1; flappy_W(26, 227) <= 1; flappy_W(26, 228) <= 1; flappy_W(26, 229) <= 1; flappy_W(26, 230) <= 1; flappy_W(26, 231) <= 1; flappy_W(26, 232) <= 1; flappy_W(26, 233) <= 1; flappy_W(26, 234) <= 1; flappy_W(26, 235) <= 1; flappy_W(26, 236) <= 1; flappy_W(26, 237) <= 1; flappy_W(26, 238) <= 1; flappy_W(26, 239) <= 1; flappy_W(26, 240) <= 1; flappy_W(26, 241) <= 1; flappy_W(26, 242) <= 1; flappy_W(26, 243) <= 1; flappy_W(26, 244) <= 1; flappy_W(26, 245) <= 1; flappy_W(26, 246) <= 1; flappy_W(26, 247) <= 1; flappy_W(26, 248) <= 1; flappy_W(26, 249) <= 1; flappy_W(26, 250) <= 1; flappy_W(26, 251) <= 1; flappy_W(26, 252) <= 0; flappy_W(26, 253) <= 0; flappy_W(26, 254) <= 0; flappy_W(26, 255) <= 0; flappy_W(26, 256) <= 0; flappy_W(26, 257) <= 0; flappy_W(26, 258) <= 0; flappy_W(26, 259) <= 0; flappy_W(26, 260) <= 0; flappy_W(26, 261) <= 0; flappy_W(26, 262) <= 0; flappy_W(26, 263) <= 0; flappy_W(26, 264) <= 0; flappy_W(26, 265) <= 0; flappy_W(26, 266) <= 0; flappy_W(26, 267) <= 0; flappy_W(26, 268) <= 0; flappy_W(26, 269) <= 0; flappy_W(26, 270) <= 0; flappy_W(26, 271) <= 0; flappy_W(26, 272) <= 0; flappy_W(26, 273) <= 0; flappy_W(26, 274) <= 0; flappy_W(26, 275) <= 0; flappy_W(26, 276) <= 0; flappy_W(26, 277) <= 0; flappy_W(26, 278) <= 0; flappy_W(26, 279) <= 0; flappy_W(26, 280) <= 0; flappy_W(26, 281) <= 0; flappy_W(26, 282) <= 1; flappy_W(26, 283) <= 1; flappy_W(26, 284) <= 1; flappy_W(26, 285) <= 1; flappy_W(26, 286) <= 1; flappy_W(26, 287) <= 1; flappy_W(26, 288) <= 1; flappy_W(26, 289) <= 1; flappy_W(26, 290) <= 1; flappy_W(26, 291) <= 1; flappy_W(26, 292) <= 1; flappy_W(26, 293) <= 1; flappy_W(26, 294) <= 1; flappy_W(26, 295) <= 1; flappy_W(26, 296) <= 1; flappy_W(26, 297) <= 1; flappy_W(26, 298) <= 1; flappy_W(26, 299) <= 1; flappy_W(26, 300) <= 1; flappy_W(26, 301) <= 1; flappy_W(26, 302) <= 1; flappy_W(26, 303) <= 1; flappy_W(26, 304) <= 1; flappy_W(26, 305) <= 1; flappy_W(26, 306) <= 0; flappy_W(26, 307) <= 0; flappy_W(26, 308) <= 0; flappy_W(26, 309) <= 0; flappy_W(26, 310) <= 0; flappy_W(26, 311) <= 0; flappy_W(26, 312) <= 0; flappy_W(26, 313) <= 0; flappy_W(26, 314) <= 0; flappy_W(26, 315) <= 0; flappy_W(26, 316) <= 0; flappy_W(26, 317) <= 0; flappy_W(26, 318) <= 0; flappy_W(26, 319) <= 0; flappy_W(26, 320) <= 0; flappy_W(26, 321) <= 0; flappy_W(26, 322) <= 0; flappy_W(26, 323) <= 0; flappy_W(26, 324) <= 0; flappy_W(26, 325) <= 0; flappy_W(26, 326) <= 0; flappy_W(26, 327) <= 0; flappy_W(26, 328) <= 0; flappy_W(26, 329) <= 0; flappy_W(26, 330) <= 0; flappy_W(26, 331) <= 0; flappy_W(26, 332) <= 0; flappy_W(26, 333) <= 0; flappy_W(26, 334) <= 0; flappy_W(26, 335) <= 0; flappy_W(26, 336) <= 0; flappy_W(26, 337) <= 0; flappy_W(26, 338) <= 0; flappy_W(26, 339) <= 0; flappy_W(26, 340) <= 0; flappy_W(26, 341) <= 0; flappy_W(26, 342) <= 0; flappy_W(26, 343) <= 0; flappy_W(26, 344) <= 0; flappy_W(26, 345) <= 0; flappy_W(26, 346) <= 0; flappy_W(26, 347) <= 0; flappy_W(26, 348) <= 0; flappy_W(26, 349) <= 0; flappy_W(26, 350) <= 0; flappy_W(26, 351) <= 0; flappy_W(26, 352) <= 0; flappy_W(26, 353) <= 0; flappy_W(26, 354) <= 0; flappy_W(26, 355) <= 0; flappy_W(26, 356) <= 0; flappy_W(26, 357) <= 0; flappy_W(26, 358) <= 0; flappy_W(26, 359) <= 0; flappy_W(26, 360) <= 0; flappy_W(26, 361) <= 0; flappy_W(26, 362) <= 0; flappy_W(26, 363) <= 0; flappy_W(26, 364) <= 0; flappy_W(26, 365) <= 0; flappy_W(26, 366) <= 0; flappy_W(26, 367) <= 0; flappy_W(26, 368) <= 0; flappy_W(26, 369) <= 0; flappy_W(26, 370) <= 0; flappy_W(26, 371) <= 0; flappy_W(26, 372) <= 0; flappy_W(26, 373) <= 0; flappy_W(26, 374) <= 0; flappy_W(26, 375) <= 0; flappy_W(26, 376) <= 0; flappy_W(26, 377) <= 0; flappy_W(26, 378) <= 0; flappy_W(26, 379) <= 0; flappy_W(26, 380) <= 0; flappy_W(26, 381) <= 0; flappy_W(26, 382) <= 0; flappy_W(26, 383) <= 0; flappy_W(26, 384) <= 0; flappy_W(26, 385) <= 0; flappy_W(26, 386) <= 0; flappy_W(26, 387) <= 0; flappy_W(26, 388) <= 0; flappy_W(26, 389) <= 0; flappy_W(26, 390) <= 0; flappy_W(26, 391) <= 0; flappy_W(26, 392) <= 0; flappy_W(26, 393) <= 0; flappy_W(26, 394) <= 0; flappy_W(26, 395) <= 0; flappy_W(26, 396) <= 0; flappy_W(26, 397) <= 0; flappy_W(26, 398) <= 0; flappy_W(26, 399) <= 0; flappy_W(26, 400) <= 0; flappy_W(26, 401) <= 0; flappy_W(26, 402) <= 1; flappy_W(26, 403) <= 1; flappy_W(26, 404) <= 1; flappy_W(26, 405) <= 1; flappy_W(26, 406) <= 1; flappy_W(26, 407) <= 1; flappy_W(26, 408) <= 1; flappy_W(26, 409) <= 1; flappy_W(26, 410) <= 1; flappy_W(26, 411) <= 1; flappy_W(26, 412) <= 1; flappy_W(26, 413) <= 1; flappy_W(26, 414) <= 1; flappy_W(26, 415) <= 1; flappy_W(26, 416) <= 1; flappy_W(26, 417) <= 1; flappy_W(26, 418) <= 1; flappy_W(26, 419) <= 1; flappy_W(26, 420) <= 1; flappy_W(26, 421) <= 1; flappy_W(26, 422) <= 1; flappy_W(26, 423) <= 1; flappy_W(26, 424) <= 1; flappy_W(26, 425) <= 1; flappy_W(26, 426) <= 1; flappy_W(26, 427) <= 1; flappy_W(26, 428) <= 1; flappy_W(26, 429) <= 1; flappy_W(26, 430) <= 1; flappy_W(26, 431) <= 1; flappy_W(26, 432) <= 0; flappy_W(26, 433) <= 0; flappy_W(26, 434) <= 0; flappy_W(26, 435) <= 0; flappy_W(26, 436) <= 0; flappy_W(26, 437) <= 0; flappy_W(26, 438) <= 0; flappy_W(26, 439) <= 0; flappy_W(26, 440) <= 0; flappy_W(26, 441) <= 0; flappy_W(26, 442) <= 0; flappy_W(26, 443) <= 0; flappy_W(26, 444) <= 0; flappy_W(26, 445) <= 0; flappy_W(26, 446) <= 0; flappy_W(26, 447) <= 0; flappy_W(26, 448) <= 0; flappy_W(26, 449) <= 0; flappy_W(26, 450) <= 0; flappy_W(26, 451) <= 0; flappy_W(26, 452) <= 0; flappy_W(26, 453) <= 0; flappy_W(26, 454) <= 0; flappy_W(26, 455) <= 0; flappy_W(26, 456) <= 0; flappy_W(26, 457) <= 0; flappy_W(26, 458) <= 0; flappy_W(26, 459) <= 0; flappy_W(26, 460) <= 0; flappy_W(26, 461) <= 0; flappy_W(26, 462) <= 0; flappy_W(26, 463) <= 0; flappy_W(26, 464) <= 0; flappy_W(26, 465) <= 0; flappy_W(26, 466) <= 0; flappy_W(26, 467) <= 0; flappy_W(26, 468) <= 1; flappy_W(26, 469) <= 1; flappy_W(26, 470) <= 1; flappy_W(26, 471) <= 1; flappy_W(26, 472) <= 1; flappy_W(26, 473) <= 1; flappy_W(26, 474) <= 1; flappy_W(26, 475) <= 1; flappy_W(26, 476) <= 1; flappy_W(26, 477) <= 1; flappy_W(26, 478) <= 1; flappy_W(26, 479) <= 1; flappy_W(26, 480) <= 0; flappy_W(26, 481) <= 0; flappy_W(26, 482) <= 0; flappy_W(26, 483) <= 0; flappy_W(26, 484) <= 0; flappy_W(26, 485) <= 0; flappy_W(26, 486) <= 0; flappy_W(26, 487) <= 0; flappy_W(26, 488) <= 0; flappy_W(26, 489) <= 0; flappy_W(26, 490) <= 0; flappy_W(26, 491) <= 0; flappy_W(26, 492) <= 0; flappy_W(26, 493) <= 0; flappy_W(26, 494) <= 0; flappy_W(26, 495) <= 0; flappy_W(26, 496) <= 0; flappy_W(26, 497) <= 0; flappy_W(26, 498) <= 0; flappy_W(26, 499) <= 0; flappy_W(26, 500) <= 0; flappy_W(26, 501) <= 0; flappy_W(26, 502) <= 0; flappy_W(26, 503) <= 0; flappy_W(26, 504) <= 0; flappy_W(26, 505) <= 0; flappy_W(26, 506) <= 0; flappy_W(26, 507) <= 0; flappy_W(26, 508) <= 0; flappy_W(26, 509) <= 0; flappy_W(26, 510) <= 1; flappy_W(26, 511) <= 1; flappy_W(26, 512) <= 1; flappy_W(26, 513) <= 1; flappy_W(26, 514) <= 1; flappy_W(26, 515) <= 1; flappy_W(26, 516) <= 1; flappy_W(26, 517) <= 1; flappy_W(26, 518) <= 1; flappy_W(26, 519) <= 1; flappy_W(26, 520) <= 1; flappy_W(26, 521) <= 1; flappy_W(26, 522) <= 1; flappy_W(26, 523) <= 1; flappy_W(26, 524) <= 1; flappy_W(26, 525) <= 1; flappy_W(26, 526) <= 1; flappy_W(26, 527) <= 1; flappy_W(26, 528) <= 1; flappy_W(26, 529) <= 1; flappy_W(26, 530) <= 1; flappy_W(26, 531) <= 1; flappy_W(26, 532) <= 1; flappy_W(26, 533) <= 1; flappy_W(26, 534) <= 1; flappy_W(26, 535) <= 1; flappy_W(26, 536) <= 1; flappy_W(26, 537) <= 1; flappy_W(26, 538) <= 1; flappy_W(26, 539) <= 1; flappy_W(26, 540) <= 0; flappy_W(26, 541) <= 0; flappy_W(26, 542) <= 0; flappy_W(26, 543) <= 0; flappy_W(26, 544) <= 0; flappy_W(26, 545) <= 0; flappy_W(26, 546) <= 0; flappy_W(26, 547) <= 0; flappy_W(26, 548) <= 0; flappy_W(26, 549) <= 0; flappy_W(26, 550) <= 0; flappy_W(26, 551) <= 0; flappy_W(26, 552) <= 0; flappy_W(26, 553) <= 0; flappy_W(26, 554) <= 0; flappy_W(26, 555) <= 0; flappy_W(26, 556) <= 0; flappy_W(26, 557) <= 0; flappy_W(26, 558) <= 0; flappy_W(26, 559) <= 0; flappy_W(26, 560) <= 0; flappy_W(26, 561) <= 0; flappy_W(26, 562) <= 0; flappy_W(26, 563) <= 0; flappy_W(26, 564) <= 1; flappy_W(26, 565) <= 1; flappy_W(26, 566) <= 1; flappy_W(26, 567) <= 1; flappy_W(26, 568) <= 1; flappy_W(26, 569) <= 1; flappy_W(26, 570) <= 1; flappy_W(26, 571) <= 1; flappy_W(26, 572) <= 1; flappy_W(26, 573) <= 1; flappy_W(26, 574) <= 1; flappy_W(26, 575) <= 1; flappy_W(26, 576) <= 0; flappy_W(26, 577) <= 0; flappy_W(26, 578) <= 0; flappy_W(26, 579) <= 0; flappy_W(26, 580) <= 0; flappy_W(26, 581) <= 0; flappy_W(26, 582) <= 0; flappy_W(26, 583) <= 0; flappy_W(26, 584) <= 0; flappy_W(26, 585) <= 0; flappy_W(26, 586) <= 0; flappy_W(26, 587) <= 0; flappy_W(26, 588) <= 1; flappy_W(26, 589) <= 1; flappy_W(26, 590) <= 1; flappy_W(26, 591) <= 1; flappy_W(26, 592) <= 1; flappy_W(26, 593) <= 1; 
flappy_W(27, 0) <= 0; flappy_W(27, 1) <= 0; flappy_W(27, 2) <= 0; flappy_W(27, 3) <= 0; flappy_W(27, 4) <= 0; flappy_W(27, 5) <= 0; flappy_W(27, 6) <= 1; flappy_W(27, 7) <= 1; flappy_W(27, 8) <= 1; flappy_W(27, 9) <= 1; flappy_W(27, 10) <= 1; flappy_W(27, 11) <= 1; flappy_W(27, 12) <= 1; flappy_W(27, 13) <= 1; flappy_W(27, 14) <= 1; flappy_W(27, 15) <= 1; flappy_W(27, 16) <= 1; flappy_W(27, 17) <= 1; flappy_W(27, 18) <= 1; flappy_W(27, 19) <= 1; flappy_W(27, 20) <= 1; flappy_W(27, 21) <= 1; flappy_W(27, 22) <= 1; flappy_W(27, 23) <= 1; flappy_W(27, 24) <= 1; flappy_W(27, 25) <= 1; flappy_W(27, 26) <= 1; flappy_W(27, 27) <= 1; flappy_W(27, 28) <= 1; flappy_W(27, 29) <= 1; flappy_W(27, 30) <= 0; flappy_W(27, 31) <= 0; flappy_W(27, 32) <= 0; flappy_W(27, 33) <= 0; flappy_W(27, 34) <= 0; flappy_W(27, 35) <= 0; flappy_W(27, 36) <= 0; flappy_W(27, 37) <= 0; flappy_W(27, 38) <= 0; flappy_W(27, 39) <= 0; flappy_W(27, 40) <= 0; flappy_W(27, 41) <= 0; flappy_W(27, 42) <= 0; flappy_W(27, 43) <= 0; flappy_W(27, 44) <= 0; flappy_W(27, 45) <= 0; flappy_W(27, 46) <= 0; flappy_W(27, 47) <= 0; flappy_W(27, 48) <= 0; flappy_W(27, 49) <= 0; flappy_W(27, 50) <= 0; flappy_W(27, 51) <= 0; flappy_W(27, 52) <= 0; flappy_W(27, 53) <= 0; flappy_W(27, 54) <= 0; flappy_W(27, 55) <= 0; flappy_W(27, 56) <= 0; flappy_W(27, 57) <= 0; flappy_W(27, 58) <= 0; flappy_W(27, 59) <= 0; flappy_W(27, 60) <= 1; flappy_W(27, 61) <= 1; flappy_W(27, 62) <= 1; flappy_W(27, 63) <= 1; flappy_W(27, 64) <= 1; flappy_W(27, 65) <= 1; flappy_W(27, 66) <= 1; flappy_W(27, 67) <= 1; flappy_W(27, 68) <= 1; flappy_W(27, 69) <= 1; flappy_W(27, 70) <= 1; flappy_W(27, 71) <= 1; flappy_W(27, 72) <= 0; flappy_W(27, 73) <= 0; flappy_W(27, 74) <= 0; flappy_W(27, 75) <= 0; flappy_W(27, 76) <= 0; flappy_W(27, 77) <= 0; flappy_W(27, 78) <= 0; flappy_W(27, 79) <= 0; flappy_W(27, 80) <= 0; flappy_W(27, 81) <= 0; flappy_W(27, 82) <= 0; flappy_W(27, 83) <= 0; flappy_W(27, 84) <= 0; flappy_W(27, 85) <= 0; flappy_W(27, 86) <= 0; flappy_W(27, 87) <= 0; flappy_W(27, 88) <= 0; flappy_W(27, 89) <= 0; flappy_W(27, 90) <= 0; flappy_W(27, 91) <= 0; flappy_W(27, 92) <= 0; flappy_W(27, 93) <= 0; flappy_W(27, 94) <= 0; flappy_W(27, 95) <= 0; flappy_W(27, 96) <= 0; flappy_W(27, 97) <= 0; flappy_W(27, 98) <= 0; flappy_W(27, 99) <= 0; flappy_W(27, 100) <= 0; flappy_W(27, 101) <= 0; flappy_W(27, 102) <= 0; flappy_W(27, 103) <= 0; flappy_W(27, 104) <= 0; flappy_W(27, 105) <= 0; flappy_W(27, 106) <= 0; flappy_W(27, 107) <= 0; flappy_W(27, 108) <= 1; flappy_W(27, 109) <= 1; flappy_W(27, 110) <= 1; flappy_W(27, 111) <= 1; flappy_W(27, 112) <= 1; flappy_W(27, 113) <= 1; flappy_W(27, 114) <= 1; flappy_W(27, 115) <= 1; flappy_W(27, 116) <= 1; flappy_W(27, 117) <= 1; flappy_W(27, 118) <= 1; flappy_W(27, 119) <= 1; flappy_W(27, 120) <= 0; flappy_W(27, 121) <= 0; flappy_W(27, 122) <= 0; flappy_W(27, 123) <= 0; flappy_W(27, 124) <= 0; flappy_W(27, 125) <= 0; flappy_W(27, 126) <= 0; flappy_W(27, 127) <= 0; flappy_W(27, 128) <= 0; flappy_W(27, 129) <= 0; flappy_W(27, 130) <= 0; flappy_W(27, 131) <= 0; flappy_W(27, 132) <= 0; flappy_W(27, 133) <= 0; flappy_W(27, 134) <= 0; flappy_W(27, 135) <= 0; flappy_W(27, 136) <= 0; flappy_W(27, 137) <= 0; flappy_W(27, 138) <= 1; flappy_W(27, 139) <= 1; flappy_W(27, 140) <= 1; flappy_W(27, 141) <= 1; flappy_W(27, 142) <= 1; flappy_W(27, 143) <= 1; flappy_W(27, 144) <= 1; flappy_W(27, 145) <= 1; flappy_W(27, 146) <= 1; flappy_W(27, 147) <= 1; flappy_W(27, 148) <= 1; flappy_W(27, 149) <= 1; flappy_W(27, 150) <= 0; flappy_W(27, 151) <= 0; flappy_W(27, 152) <= 0; flappy_W(27, 153) <= 0; flappy_W(27, 154) <= 0; flappy_W(27, 155) <= 0; flappy_W(27, 156) <= 0; flappy_W(27, 157) <= 0; flappy_W(27, 158) <= 0; flappy_W(27, 159) <= 0; flappy_W(27, 160) <= 0; flappy_W(27, 161) <= 0; flappy_W(27, 162) <= 0; flappy_W(27, 163) <= 0; flappy_W(27, 164) <= 0; flappy_W(27, 165) <= 0; flappy_W(27, 166) <= 0; flappy_W(27, 167) <= 0; flappy_W(27, 168) <= 1; flappy_W(27, 169) <= 1; flappy_W(27, 170) <= 1; flappy_W(27, 171) <= 1; flappy_W(27, 172) <= 1; flappy_W(27, 173) <= 1; flappy_W(27, 174) <= 1; flappy_W(27, 175) <= 1; flappy_W(27, 176) <= 1; flappy_W(27, 177) <= 1; flappy_W(27, 178) <= 1; flappy_W(27, 179) <= 1; flappy_W(27, 180) <= 1; flappy_W(27, 181) <= 1; flappy_W(27, 182) <= 1; flappy_W(27, 183) <= 1; flappy_W(27, 184) <= 1; flappy_W(27, 185) <= 1; flappy_W(27, 186) <= 1; flappy_W(27, 187) <= 1; flappy_W(27, 188) <= 1; flappy_W(27, 189) <= 1; flappy_W(27, 190) <= 1; flappy_W(27, 191) <= 1; flappy_W(27, 192) <= 1; flappy_W(27, 193) <= 1; flappy_W(27, 194) <= 1; flappy_W(27, 195) <= 1; flappy_W(27, 196) <= 1; flappy_W(27, 197) <= 1; flappy_W(27, 198) <= 0; flappy_W(27, 199) <= 0; flappy_W(27, 200) <= 0; flappy_W(27, 201) <= 0; flappy_W(27, 202) <= 0; flappy_W(27, 203) <= 0; flappy_W(27, 204) <= 0; flappy_W(27, 205) <= 0; flappy_W(27, 206) <= 0; flappy_W(27, 207) <= 0; flappy_W(27, 208) <= 0; flappy_W(27, 209) <= 0; flappy_W(27, 210) <= 0; flappy_W(27, 211) <= 0; flappy_W(27, 212) <= 0; flappy_W(27, 213) <= 0; flappy_W(27, 214) <= 0; flappy_W(27, 215) <= 0; flappy_W(27, 216) <= 0; flappy_W(27, 217) <= 0; flappy_W(27, 218) <= 0; flappy_W(27, 219) <= 0; flappy_W(27, 220) <= 0; flappy_W(27, 221) <= 0; flappy_W(27, 222) <= 1; flappy_W(27, 223) <= 1; flappy_W(27, 224) <= 1; flappy_W(27, 225) <= 1; flappy_W(27, 226) <= 1; flappy_W(27, 227) <= 1; flappy_W(27, 228) <= 1; flappy_W(27, 229) <= 1; flappy_W(27, 230) <= 1; flappy_W(27, 231) <= 1; flappy_W(27, 232) <= 1; flappy_W(27, 233) <= 1; flappy_W(27, 234) <= 1; flappy_W(27, 235) <= 1; flappy_W(27, 236) <= 1; flappy_W(27, 237) <= 1; flappy_W(27, 238) <= 1; flappy_W(27, 239) <= 1; flappy_W(27, 240) <= 1; flappy_W(27, 241) <= 1; flappy_W(27, 242) <= 1; flappy_W(27, 243) <= 1; flappy_W(27, 244) <= 1; flappy_W(27, 245) <= 1; flappy_W(27, 246) <= 1; flappy_W(27, 247) <= 1; flappy_W(27, 248) <= 1; flappy_W(27, 249) <= 1; flappy_W(27, 250) <= 1; flappy_W(27, 251) <= 1; flappy_W(27, 252) <= 0; flappy_W(27, 253) <= 0; flappy_W(27, 254) <= 0; flappy_W(27, 255) <= 0; flappy_W(27, 256) <= 0; flappy_W(27, 257) <= 0; flappy_W(27, 258) <= 0; flappy_W(27, 259) <= 0; flappy_W(27, 260) <= 0; flappy_W(27, 261) <= 0; flappy_W(27, 262) <= 0; flappy_W(27, 263) <= 0; flappy_W(27, 264) <= 0; flappy_W(27, 265) <= 0; flappy_W(27, 266) <= 0; flappy_W(27, 267) <= 0; flappy_W(27, 268) <= 0; flappy_W(27, 269) <= 0; flappy_W(27, 270) <= 0; flappy_W(27, 271) <= 0; flappy_W(27, 272) <= 0; flappy_W(27, 273) <= 0; flappy_W(27, 274) <= 0; flappy_W(27, 275) <= 0; flappy_W(27, 276) <= 0; flappy_W(27, 277) <= 0; flappy_W(27, 278) <= 0; flappy_W(27, 279) <= 0; flappy_W(27, 280) <= 0; flappy_W(27, 281) <= 0; flappy_W(27, 282) <= 1; flappy_W(27, 283) <= 1; flappy_W(27, 284) <= 1; flappy_W(27, 285) <= 1; flappy_W(27, 286) <= 1; flappy_W(27, 287) <= 1; flappy_W(27, 288) <= 1; flappy_W(27, 289) <= 1; flappy_W(27, 290) <= 1; flappy_W(27, 291) <= 1; flappy_W(27, 292) <= 1; flappy_W(27, 293) <= 1; flappy_W(27, 294) <= 1; flappy_W(27, 295) <= 1; flappy_W(27, 296) <= 1; flappy_W(27, 297) <= 1; flappy_W(27, 298) <= 1; flappy_W(27, 299) <= 1; flappy_W(27, 300) <= 1; flappy_W(27, 301) <= 1; flappy_W(27, 302) <= 1; flappy_W(27, 303) <= 1; flappy_W(27, 304) <= 1; flappy_W(27, 305) <= 1; flappy_W(27, 306) <= 0; flappy_W(27, 307) <= 0; flappy_W(27, 308) <= 0; flappy_W(27, 309) <= 0; flappy_W(27, 310) <= 0; flappy_W(27, 311) <= 0; flappy_W(27, 312) <= 0; flappy_W(27, 313) <= 0; flappy_W(27, 314) <= 0; flappy_W(27, 315) <= 0; flappy_W(27, 316) <= 0; flappy_W(27, 317) <= 0; flappy_W(27, 318) <= 0; flappy_W(27, 319) <= 0; flappy_W(27, 320) <= 0; flappy_W(27, 321) <= 0; flappy_W(27, 322) <= 0; flappy_W(27, 323) <= 0; flappy_W(27, 324) <= 0; flappy_W(27, 325) <= 0; flappy_W(27, 326) <= 0; flappy_W(27, 327) <= 0; flappy_W(27, 328) <= 0; flappy_W(27, 329) <= 0; flappy_W(27, 330) <= 0; flappy_W(27, 331) <= 0; flappy_W(27, 332) <= 0; flappy_W(27, 333) <= 0; flappy_W(27, 334) <= 0; flappy_W(27, 335) <= 0; flappy_W(27, 336) <= 0; flappy_W(27, 337) <= 0; flappy_W(27, 338) <= 0; flappy_W(27, 339) <= 0; flappy_W(27, 340) <= 0; flappy_W(27, 341) <= 0; flappy_W(27, 342) <= 0; flappy_W(27, 343) <= 0; flappy_W(27, 344) <= 0; flappy_W(27, 345) <= 0; flappy_W(27, 346) <= 0; flappy_W(27, 347) <= 0; flappy_W(27, 348) <= 0; flappy_W(27, 349) <= 0; flappy_W(27, 350) <= 0; flappy_W(27, 351) <= 0; flappy_W(27, 352) <= 0; flappy_W(27, 353) <= 0; flappy_W(27, 354) <= 0; flappy_W(27, 355) <= 0; flappy_W(27, 356) <= 0; flappy_W(27, 357) <= 0; flappy_W(27, 358) <= 0; flappy_W(27, 359) <= 0; flappy_W(27, 360) <= 0; flappy_W(27, 361) <= 0; flappy_W(27, 362) <= 0; flappy_W(27, 363) <= 0; flappy_W(27, 364) <= 0; flappy_W(27, 365) <= 0; flappy_W(27, 366) <= 0; flappy_W(27, 367) <= 0; flappy_W(27, 368) <= 0; flappy_W(27, 369) <= 0; flappy_W(27, 370) <= 0; flappy_W(27, 371) <= 0; flappy_W(27, 372) <= 0; flappy_W(27, 373) <= 0; flappy_W(27, 374) <= 0; flappy_W(27, 375) <= 0; flappy_W(27, 376) <= 0; flappy_W(27, 377) <= 0; flappy_W(27, 378) <= 0; flappy_W(27, 379) <= 0; flappy_W(27, 380) <= 0; flappy_W(27, 381) <= 0; flappy_W(27, 382) <= 0; flappy_W(27, 383) <= 0; flappy_W(27, 384) <= 0; flappy_W(27, 385) <= 0; flappy_W(27, 386) <= 0; flappy_W(27, 387) <= 0; flappy_W(27, 388) <= 0; flappy_W(27, 389) <= 0; flappy_W(27, 390) <= 0; flappy_W(27, 391) <= 0; flappy_W(27, 392) <= 0; flappy_W(27, 393) <= 0; flappy_W(27, 394) <= 0; flappy_W(27, 395) <= 0; flappy_W(27, 396) <= 0; flappy_W(27, 397) <= 0; flappy_W(27, 398) <= 0; flappy_W(27, 399) <= 0; flappy_W(27, 400) <= 0; flappy_W(27, 401) <= 0; flappy_W(27, 402) <= 1; flappy_W(27, 403) <= 1; flappy_W(27, 404) <= 1; flappy_W(27, 405) <= 1; flappy_W(27, 406) <= 1; flappy_W(27, 407) <= 1; flappy_W(27, 408) <= 1; flappy_W(27, 409) <= 1; flappy_W(27, 410) <= 1; flappy_W(27, 411) <= 1; flappy_W(27, 412) <= 1; flappy_W(27, 413) <= 1; flappy_W(27, 414) <= 1; flappy_W(27, 415) <= 1; flappy_W(27, 416) <= 1; flappy_W(27, 417) <= 1; flappy_W(27, 418) <= 1; flappy_W(27, 419) <= 1; flappy_W(27, 420) <= 1; flappy_W(27, 421) <= 1; flappy_W(27, 422) <= 1; flappy_W(27, 423) <= 1; flappy_W(27, 424) <= 1; flappy_W(27, 425) <= 1; flappy_W(27, 426) <= 1; flappy_W(27, 427) <= 1; flappy_W(27, 428) <= 1; flappy_W(27, 429) <= 1; flappy_W(27, 430) <= 1; flappy_W(27, 431) <= 1; flappy_W(27, 432) <= 0; flappy_W(27, 433) <= 0; flappy_W(27, 434) <= 0; flappy_W(27, 435) <= 0; flappy_W(27, 436) <= 0; flappy_W(27, 437) <= 0; flappy_W(27, 438) <= 0; flappy_W(27, 439) <= 0; flappy_W(27, 440) <= 0; flappy_W(27, 441) <= 0; flappy_W(27, 442) <= 0; flappy_W(27, 443) <= 0; flappy_W(27, 444) <= 0; flappy_W(27, 445) <= 0; flappy_W(27, 446) <= 0; flappy_W(27, 447) <= 0; flappy_W(27, 448) <= 0; flappy_W(27, 449) <= 0; flappy_W(27, 450) <= 0; flappy_W(27, 451) <= 0; flappy_W(27, 452) <= 0; flappy_W(27, 453) <= 0; flappy_W(27, 454) <= 0; flappy_W(27, 455) <= 0; flappy_W(27, 456) <= 0; flappy_W(27, 457) <= 0; flappy_W(27, 458) <= 0; flappy_W(27, 459) <= 0; flappy_W(27, 460) <= 0; flappy_W(27, 461) <= 0; flappy_W(27, 462) <= 0; flappy_W(27, 463) <= 0; flappy_W(27, 464) <= 0; flappy_W(27, 465) <= 0; flappy_W(27, 466) <= 0; flappy_W(27, 467) <= 0; flappy_W(27, 468) <= 1; flappy_W(27, 469) <= 1; flappy_W(27, 470) <= 1; flappy_W(27, 471) <= 1; flappy_W(27, 472) <= 1; flappy_W(27, 473) <= 1; flappy_W(27, 474) <= 1; flappy_W(27, 475) <= 1; flappy_W(27, 476) <= 1; flappy_W(27, 477) <= 1; flappy_W(27, 478) <= 1; flappy_W(27, 479) <= 1; flappy_W(27, 480) <= 0; flappy_W(27, 481) <= 0; flappy_W(27, 482) <= 0; flappy_W(27, 483) <= 0; flappy_W(27, 484) <= 0; flappy_W(27, 485) <= 0; flappy_W(27, 486) <= 0; flappy_W(27, 487) <= 0; flappy_W(27, 488) <= 0; flappy_W(27, 489) <= 0; flappy_W(27, 490) <= 0; flappy_W(27, 491) <= 0; flappy_W(27, 492) <= 0; flappy_W(27, 493) <= 0; flappy_W(27, 494) <= 0; flappy_W(27, 495) <= 0; flappy_W(27, 496) <= 0; flappy_W(27, 497) <= 0; flappy_W(27, 498) <= 0; flappy_W(27, 499) <= 0; flappy_W(27, 500) <= 0; flappy_W(27, 501) <= 0; flappy_W(27, 502) <= 0; flappy_W(27, 503) <= 0; flappy_W(27, 504) <= 0; flappy_W(27, 505) <= 0; flappy_W(27, 506) <= 0; flappy_W(27, 507) <= 0; flappy_W(27, 508) <= 0; flappy_W(27, 509) <= 0; flappy_W(27, 510) <= 1; flappy_W(27, 511) <= 1; flappy_W(27, 512) <= 1; flappy_W(27, 513) <= 1; flappy_W(27, 514) <= 1; flappy_W(27, 515) <= 1; flappy_W(27, 516) <= 1; flappy_W(27, 517) <= 1; flappy_W(27, 518) <= 1; flappy_W(27, 519) <= 1; flappy_W(27, 520) <= 1; flappy_W(27, 521) <= 1; flappy_W(27, 522) <= 1; flappy_W(27, 523) <= 1; flappy_W(27, 524) <= 1; flappy_W(27, 525) <= 1; flappy_W(27, 526) <= 1; flappy_W(27, 527) <= 1; flappy_W(27, 528) <= 1; flappy_W(27, 529) <= 1; flappy_W(27, 530) <= 1; flappy_W(27, 531) <= 1; flappy_W(27, 532) <= 1; flappy_W(27, 533) <= 1; flappy_W(27, 534) <= 1; flappy_W(27, 535) <= 1; flappy_W(27, 536) <= 1; flappy_W(27, 537) <= 1; flappy_W(27, 538) <= 1; flappy_W(27, 539) <= 1; flappy_W(27, 540) <= 0; flappy_W(27, 541) <= 0; flappy_W(27, 542) <= 0; flappy_W(27, 543) <= 0; flappy_W(27, 544) <= 0; flappy_W(27, 545) <= 0; flappy_W(27, 546) <= 0; flappy_W(27, 547) <= 0; flappy_W(27, 548) <= 0; flappy_W(27, 549) <= 0; flappy_W(27, 550) <= 0; flappy_W(27, 551) <= 0; flappy_W(27, 552) <= 0; flappy_W(27, 553) <= 0; flappy_W(27, 554) <= 0; flappy_W(27, 555) <= 0; flappy_W(27, 556) <= 0; flappy_W(27, 557) <= 0; flappy_W(27, 558) <= 0; flappy_W(27, 559) <= 0; flappy_W(27, 560) <= 0; flappy_W(27, 561) <= 0; flappy_W(27, 562) <= 0; flappy_W(27, 563) <= 0; flappy_W(27, 564) <= 1; flappy_W(27, 565) <= 1; flappy_W(27, 566) <= 1; flappy_W(27, 567) <= 1; flappy_W(27, 568) <= 1; flappy_W(27, 569) <= 1; flappy_W(27, 570) <= 1; flappy_W(27, 571) <= 1; flappy_W(27, 572) <= 1; flappy_W(27, 573) <= 1; flappy_W(27, 574) <= 1; flappy_W(27, 575) <= 1; flappy_W(27, 576) <= 0; flappy_W(27, 577) <= 0; flappy_W(27, 578) <= 0; flappy_W(27, 579) <= 0; flappy_W(27, 580) <= 0; flappy_W(27, 581) <= 0; flappy_W(27, 582) <= 0; flappy_W(27, 583) <= 0; flappy_W(27, 584) <= 0; flappy_W(27, 585) <= 0; flappy_W(27, 586) <= 0; flappy_W(27, 587) <= 0; flappy_W(27, 588) <= 1; flappy_W(27, 589) <= 1; flappy_W(27, 590) <= 1; flappy_W(27, 591) <= 1; flappy_W(27, 592) <= 1; flappy_W(27, 593) <= 1; 
flappy_W(28, 0) <= 0; flappy_W(28, 1) <= 0; flappy_W(28, 2) <= 0; flappy_W(28, 3) <= 0; flappy_W(28, 4) <= 0; flappy_W(28, 5) <= 0; flappy_W(28, 6) <= 1; flappy_W(28, 7) <= 1; flappy_W(28, 8) <= 1; flappy_W(28, 9) <= 1; flappy_W(28, 10) <= 1; flappy_W(28, 11) <= 1; flappy_W(28, 12) <= 1; flappy_W(28, 13) <= 1; flappy_W(28, 14) <= 1; flappy_W(28, 15) <= 1; flappy_W(28, 16) <= 1; flappy_W(28, 17) <= 1; flappy_W(28, 18) <= 1; flappy_W(28, 19) <= 1; flappy_W(28, 20) <= 1; flappy_W(28, 21) <= 1; flappy_W(28, 22) <= 1; flappy_W(28, 23) <= 1; flappy_W(28, 24) <= 1; flappy_W(28, 25) <= 1; flappy_W(28, 26) <= 1; flappy_W(28, 27) <= 1; flappy_W(28, 28) <= 1; flappy_W(28, 29) <= 1; flappy_W(28, 30) <= 0; flappy_W(28, 31) <= 0; flappy_W(28, 32) <= 0; flappy_W(28, 33) <= 0; flappy_W(28, 34) <= 0; flappy_W(28, 35) <= 0; flappy_W(28, 36) <= 0; flappy_W(28, 37) <= 0; flappy_W(28, 38) <= 0; flappy_W(28, 39) <= 0; flappy_W(28, 40) <= 0; flappy_W(28, 41) <= 0; flappy_W(28, 42) <= 0; flappy_W(28, 43) <= 0; flappy_W(28, 44) <= 0; flappy_W(28, 45) <= 0; flappy_W(28, 46) <= 0; flappy_W(28, 47) <= 0; flappy_W(28, 48) <= 0; flappy_W(28, 49) <= 0; flappy_W(28, 50) <= 0; flappy_W(28, 51) <= 0; flappy_W(28, 52) <= 0; flappy_W(28, 53) <= 0; flappy_W(28, 54) <= 0; flappy_W(28, 55) <= 0; flappy_W(28, 56) <= 0; flappy_W(28, 57) <= 0; flappy_W(28, 58) <= 0; flappy_W(28, 59) <= 0; flappy_W(28, 60) <= 1; flappy_W(28, 61) <= 1; flappy_W(28, 62) <= 1; flappy_W(28, 63) <= 1; flappy_W(28, 64) <= 1; flappy_W(28, 65) <= 1; flappy_W(28, 66) <= 1; flappy_W(28, 67) <= 1; flappy_W(28, 68) <= 1; flappy_W(28, 69) <= 1; flappy_W(28, 70) <= 1; flappy_W(28, 71) <= 1; flappy_W(28, 72) <= 0; flappy_W(28, 73) <= 0; flappy_W(28, 74) <= 0; flappy_W(28, 75) <= 0; flappy_W(28, 76) <= 0; flappy_W(28, 77) <= 0; flappy_W(28, 78) <= 0; flappy_W(28, 79) <= 0; flappy_W(28, 80) <= 0; flappy_W(28, 81) <= 0; flappy_W(28, 82) <= 0; flappy_W(28, 83) <= 0; flappy_W(28, 84) <= 0; flappy_W(28, 85) <= 0; flappy_W(28, 86) <= 0; flappy_W(28, 87) <= 0; flappy_W(28, 88) <= 0; flappy_W(28, 89) <= 0; flappy_W(28, 90) <= 0; flappy_W(28, 91) <= 0; flappy_W(28, 92) <= 0; flappy_W(28, 93) <= 0; flappy_W(28, 94) <= 0; flappy_W(28, 95) <= 0; flappy_W(28, 96) <= 0; flappy_W(28, 97) <= 0; flappy_W(28, 98) <= 0; flappy_W(28, 99) <= 0; flappy_W(28, 100) <= 0; flappy_W(28, 101) <= 0; flappy_W(28, 102) <= 0; flappy_W(28, 103) <= 0; flappy_W(28, 104) <= 0; flappy_W(28, 105) <= 0; flappy_W(28, 106) <= 0; flappy_W(28, 107) <= 0; flappy_W(28, 108) <= 1; flappy_W(28, 109) <= 1; flappy_W(28, 110) <= 1; flappy_W(28, 111) <= 1; flappy_W(28, 112) <= 1; flappy_W(28, 113) <= 1; flappy_W(28, 114) <= 1; flappy_W(28, 115) <= 1; flappy_W(28, 116) <= 1; flappy_W(28, 117) <= 1; flappy_W(28, 118) <= 1; flappy_W(28, 119) <= 1; flappy_W(28, 120) <= 0; flappy_W(28, 121) <= 0; flappy_W(28, 122) <= 0; flappy_W(28, 123) <= 0; flappy_W(28, 124) <= 0; flappy_W(28, 125) <= 0; flappy_W(28, 126) <= 0; flappy_W(28, 127) <= 0; flappy_W(28, 128) <= 0; flappy_W(28, 129) <= 0; flappy_W(28, 130) <= 0; flappy_W(28, 131) <= 0; flappy_W(28, 132) <= 0; flappy_W(28, 133) <= 0; flappy_W(28, 134) <= 0; flappy_W(28, 135) <= 0; flappy_W(28, 136) <= 0; flappy_W(28, 137) <= 0; flappy_W(28, 138) <= 1; flappy_W(28, 139) <= 1; flappy_W(28, 140) <= 1; flappy_W(28, 141) <= 1; flappy_W(28, 142) <= 1; flappy_W(28, 143) <= 1; flappy_W(28, 144) <= 1; flappy_W(28, 145) <= 1; flappy_W(28, 146) <= 1; flappy_W(28, 147) <= 1; flappy_W(28, 148) <= 1; flappy_W(28, 149) <= 1; flappy_W(28, 150) <= 0; flappy_W(28, 151) <= 0; flappy_W(28, 152) <= 0; flappy_W(28, 153) <= 0; flappy_W(28, 154) <= 0; flappy_W(28, 155) <= 0; flappy_W(28, 156) <= 0; flappy_W(28, 157) <= 0; flappy_W(28, 158) <= 0; flappy_W(28, 159) <= 0; flappy_W(28, 160) <= 0; flappy_W(28, 161) <= 0; flappy_W(28, 162) <= 0; flappy_W(28, 163) <= 0; flappy_W(28, 164) <= 0; flappy_W(28, 165) <= 0; flappy_W(28, 166) <= 0; flappy_W(28, 167) <= 0; flappy_W(28, 168) <= 1; flappy_W(28, 169) <= 1; flappy_W(28, 170) <= 1; flappy_W(28, 171) <= 1; flappy_W(28, 172) <= 1; flappy_W(28, 173) <= 1; flappy_W(28, 174) <= 1; flappy_W(28, 175) <= 1; flappy_W(28, 176) <= 1; flappy_W(28, 177) <= 1; flappy_W(28, 178) <= 1; flappy_W(28, 179) <= 1; flappy_W(28, 180) <= 1; flappy_W(28, 181) <= 1; flappy_W(28, 182) <= 1; flappy_W(28, 183) <= 1; flappy_W(28, 184) <= 1; flappy_W(28, 185) <= 1; flappy_W(28, 186) <= 1; flappy_W(28, 187) <= 1; flappy_W(28, 188) <= 1; flappy_W(28, 189) <= 1; flappy_W(28, 190) <= 1; flappy_W(28, 191) <= 1; flappy_W(28, 192) <= 1; flappy_W(28, 193) <= 1; flappy_W(28, 194) <= 1; flappy_W(28, 195) <= 1; flappy_W(28, 196) <= 1; flappy_W(28, 197) <= 1; flappy_W(28, 198) <= 0; flappy_W(28, 199) <= 0; flappy_W(28, 200) <= 0; flappy_W(28, 201) <= 0; flappy_W(28, 202) <= 0; flappy_W(28, 203) <= 0; flappy_W(28, 204) <= 0; flappy_W(28, 205) <= 0; flappy_W(28, 206) <= 0; flappy_W(28, 207) <= 0; flappy_W(28, 208) <= 0; flappy_W(28, 209) <= 0; flappy_W(28, 210) <= 0; flappy_W(28, 211) <= 0; flappy_W(28, 212) <= 0; flappy_W(28, 213) <= 0; flappy_W(28, 214) <= 0; flappy_W(28, 215) <= 0; flappy_W(28, 216) <= 0; flappy_W(28, 217) <= 0; flappy_W(28, 218) <= 0; flappy_W(28, 219) <= 0; flappy_W(28, 220) <= 0; flappy_W(28, 221) <= 0; flappy_W(28, 222) <= 1; flappy_W(28, 223) <= 1; flappy_W(28, 224) <= 1; flappy_W(28, 225) <= 1; flappy_W(28, 226) <= 1; flappy_W(28, 227) <= 1; flappy_W(28, 228) <= 1; flappy_W(28, 229) <= 1; flappy_W(28, 230) <= 1; flappy_W(28, 231) <= 1; flappy_W(28, 232) <= 1; flappy_W(28, 233) <= 1; flappy_W(28, 234) <= 1; flappy_W(28, 235) <= 1; flappy_W(28, 236) <= 1; flappy_W(28, 237) <= 1; flappy_W(28, 238) <= 1; flappy_W(28, 239) <= 1; flappy_W(28, 240) <= 1; flappy_W(28, 241) <= 1; flappy_W(28, 242) <= 1; flappy_W(28, 243) <= 1; flappy_W(28, 244) <= 1; flappy_W(28, 245) <= 1; flappy_W(28, 246) <= 1; flappy_W(28, 247) <= 1; flappy_W(28, 248) <= 1; flappy_W(28, 249) <= 1; flappy_W(28, 250) <= 1; flappy_W(28, 251) <= 1; flappy_W(28, 252) <= 0; flappy_W(28, 253) <= 0; flappy_W(28, 254) <= 0; flappy_W(28, 255) <= 0; flappy_W(28, 256) <= 0; flappy_W(28, 257) <= 0; flappy_W(28, 258) <= 0; flappy_W(28, 259) <= 0; flappy_W(28, 260) <= 0; flappy_W(28, 261) <= 0; flappy_W(28, 262) <= 0; flappy_W(28, 263) <= 0; flappy_W(28, 264) <= 0; flappy_W(28, 265) <= 0; flappy_W(28, 266) <= 0; flappy_W(28, 267) <= 0; flappy_W(28, 268) <= 0; flappy_W(28, 269) <= 0; flappy_W(28, 270) <= 0; flappy_W(28, 271) <= 0; flappy_W(28, 272) <= 0; flappy_W(28, 273) <= 0; flappy_W(28, 274) <= 0; flappy_W(28, 275) <= 0; flappy_W(28, 276) <= 0; flappy_W(28, 277) <= 0; flappy_W(28, 278) <= 0; flappy_W(28, 279) <= 0; flappy_W(28, 280) <= 0; flappy_W(28, 281) <= 0; flappy_W(28, 282) <= 1; flappy_W(28, 283) <= 1; flappy_W(28, 284) <= 1; flappy_W(28, 285) <= 1; flappy_W(28, 286) <= 1; flappy_W(28, 287) <= 1; flappy_W(28, 288) <= 1; flappy_W(28, 289) <= 1; flappy_W(28, 290) <= 1; flappy_W(28, 291) <= 1; flappy_W(28, 292) <= 1; flappy_W(28, 293) <= 1; flappy_W(28, 294) <= 1; flappy_W(28, 295) <= 1; flappy_W(28, 296) <= 1; flappy_W(28, 297) <= 1; flappy_W(28, 298) <= 1; flappy_W(28, 299) <= 1; flappy_W(28, 300) <= 1; flappy_W(28, 301) <= 1; flappy_W(28, 302) <= 1; flappy_W(28, 303) <= 1; flappy_W(28, 304) <= 1; flappy_W(28, 305) <= 1; flappy_W(28, 306) <= 0; flappy_W(28, 307) <= 0; flappy_W(28, 308) <= 0; flappy_W(28, 309) <= 0; flappy_W(28, 310) <= 0; flappy_W(28, 311) <= 0; flappy_W(28, 312) <= 0; flappy_W(28, 313) <= 0; flappy_W(28, 314) <= 0; flappy_W(28, 315) <= 0; flappy_W(28, 316) <= 0; flappy_W(28, 317) <= 0; flappy_W(28, 318) <= 0; flappy_W(28, 319) <= 0; flappy_W(28, 320) <= 0; flappy_W(28, 321) <= 0; flappy_W(28, 322) <= 0; flappy_W(28, 323) <= 0; flappy_W(28, 324) <= 0; flappy_W(28, 325) <= 0; flappy_W(28, 326) <= 0; flappy_W(28, 327) <= 0; flappy_W(28, 328) <= 0; flappy_W(28, 329) <= 0; flappy_W(28, 330) <= 0; flappy_W(28, 331) <= 0; flappy_W(28, 332) <= 0; flappy_W(28, 333) <= 0; flappy_W(28, 334) <= 0; flappy_W(28, 335) <= 0; flappy_W(28, 336) <= 0; flappy_W(28, 337) <= 0; flappy_W(28, 338) <= 0; flappy_W(28, 339) <= 0; flappy_W(28, 340) <= 0; flappy_W(28, 341) <= 0; flappy_W(28, 342) <= 0; flappy_W(28, 343) <= 0; flappy_W(28, 344) <= 0; flappy_W(28, 345) <= 0; flappy_W(28, 346) <= 0; flappy_W(28, 347) <= 0; flappy_W(28, 348) <= 0; flappy_W(28, 349) <= 0; flappy_W(28, 350) <= 0; flappy_W(28, 351) <= 0; flappy_W(28, 352) <= 0; flappy_W(28, 353) <= 0; flappy_W(28, 354) <= 0; flappy_W(28, 355) <= 0; flappy_W(28, 356) <= 0; flappy_W(28, 357) <= 0; flappy_W(28, 358) <= 0; flappy_W(28, 359) <= 0; flappy_W(28, 360) <= 0; flappy_W(28, 361) <= 0; flappy_W(28, 362) <= 0; flappy_W(28, 363) <= 0; flappy_W(28, 364) <= 0; flappy_W(28, 365) <= 0; flappy_W(28, 366) <= 0; flappy_W(28, 367) <= 0; flappy_W(28, 368) <= 0; flappy_W(28, 369) <= 0; flappy_W(28, 370) <= 0; flappy_W(28, 371) <= 0; flappy_W(28, 372) <= 0; flappy_W(28, 373) <= 0; flappy_W(28, 374) <= 0; flappy_W(28, 375) <= 0; flappy_W(28, 376) <= 0; flappy_W(28, 377) <= 0; flappy_W(28, 378) <= 0; flappy_W(28, 379) <= 0; flappy_W(28, 380) <= 0; flappy_W(28, 381) <= 0; flappy_W(28, 382) <= 0; flappy_W(28, 383) <= 0; flappy_W(28, 384) <= 0; flappy_W(28, 385) <= 0; flappy_W(28, 386) <= 0; flappy_W(28, 387) <= 0; flappy_W(28, 388) <= 0; flappy_W(28, 389) <= 0; flappy_W(28, 390) <= 0; flappy_W(28, 391) <= 0; flappy_W(28, 392) <= 0; flappy_W(28, 393) <= 0; flappy_W(28, 394) <= 0; flappy_W(28, 395) <= 0; flappy_W(28, 396) <= 0; flappy_W(28, 397) <= 0; flappy_W(28, 398) <= 0; flappy_W(28, 399) <= 0; flappy_W(28, 400) <= 0; flappy_W(28, 401) <= 0; flappy_W(28, 402) <= 1; flappy_W(28, 403) <= 1; flappy_W(28, 404) <= 1; flappy_W(28, 405) <= 1; flappy_W(28, 406) <= 1; flappy_W(28, 407) <= 1; flappy_W(28, 408) <= 1; flappy_W(28, 409) <= 1; flappy_W(28, 410) <= 1; flappy_W(28, 411) <= 1; flappy_W(28, 412) <= 1; flappy_W(28, 413) <= 1; flappy_W(28, 414) <= 1; flappy_W(28, 415) <= 1; flappy_W(28, 416) <= 1; flappy_W(28, 417) <= 1; flappy_W(28, 418) <= 1; flappy_W(28, 419) <= 1; flappy_W(28, 420) <= 1; flappy_W(28, 421) <= 1; flappy_W(28, 422) <= 1; flappy_W(28, 423) <= 1; flappy_W(28, 424) <= 1; flappy_W(28, 425) <= 1; flappy_W(28, 426) <= 1; flappy_W(28, 427) <= 1; flappy_W(28, 428) <= 1; flappy_W(28, 429) <= 1; flappy_W(28, 430) <= 1; flappy_W(28, 431) <= 1; flappy_W(28, 432) <= 0; flappy_W(28, 433) <= 0; flappy_W(28, 434) <= 0; flappy_W(28, 435) <= 0; flappy_W(28, 436) <= 0; flappy_W(28, 437) <= 0; flappy_W(28, 438) <= 0; flappy_W(28, 439) <= 0; flappy_W(28, 440) <= 0; flappy_W(28, 441) <= 0; flappy_W(28, 442) <= 0; flappy_W(28, 443) <= 0; flappy_W(28, 444) <= 0; flappy_W(28, 445) <= 0; flappy_W(28, 446) <= 0; flappy_W(28, 447) <= 0; flappy_W(28, 448) <= 0; flappy_W(28, 449) <= 0; flappy_W(28, 450) <= 0; flappy_W(28, 451) <= 0; flappy_W(28, 452) <= 0; flappy_W(28, 453) <= 0; flappy_W(28, 454) <= 0; flappy_W(28, 455) <= 0; flappy_W(28, 456) <= 0; flappy_W(28, 457) <= 0; flappy_W(28, 458) <= 0; flappy_W(28, 459) <= 0; flappy_W(28, 460) <= 0; flappy_W(28, 461) <= 0; flappy_W(28, 462) <= 0; flappy_W(28, 463) <= 0; flappy_W(28, 464) <= 0; flappy_W(28, 465) <= 0; flappy_W(28, 466) <= 0; flappy_W(28, 467) <= 0; flappy_W(28, 468) <= 1; flappy_W(28, 469) <= 1; flappy_W(28, 470) <= 1; flappy_W(28, 471) <= 1; flappy_W(28, 472) <= 1; flappy_W(28, 473) <= 1; flappy_W(28, 474) <= 1; flappy_W(28, 475) <= 1; flappy_W(28, 476) <= 1; flappy_W(28, 477) <= 1; flappy_W(28, 478) <= 1; flappy_W(28, 479) <= 1; flappy_W(28, 480) <= 0; flappy_W(28, 481) <= 0; flappy_W(28, 482) <= 0; flappy_W(28, 483) <= 0; flappy_W(28, 484) <= 0; flappy_W(28, 485) <= 0; flappy_W(28, 486) <= 0; flappy_W(28, 487) <= 0; flappy_W(28, 488) <= 0; flappy_W(28, 489) <= 0; flappy_W(28, 490) <= 0; flappy_W(28, 491) <= 0; flappy_W(28, 492) <= 0; flappy_W(28, 493) <= 0; flappy_W(28, 494) <= 0; flappy_W(28, 495) <= 0; flappy_W(28, 496) <= 0; flappy_W(28, 497) <= 0; flappy_W(28, 498) <= 0; flappy_W(28, 499) <= 0; flappy_W(28, 500) <= 0; flappy_W(28, 501) <= 0; flappy_W(28, 502) <= 0; flappy_W(28, 503) <= 0; flappy_W(28, 504) <= 0; flappy_W(28, 505) <= 0; flappy_W(28, 506) <= 0; flappy_W(28, 507) <= 0; flappy_W(28, 508) <= 0; flappy_W(28, 509) <= 0; flappy_W(28, 510) <= 1; flappy_W(28, 511) <= 1; flappy_W(28, 512) <= 1; flappy_W(28, 513) <= 1; flappy_W(28, 514) <= 1; flappy_W(28, 515) <= 1; flappy_W(28, 516) <= 1; flappy_W(28, 517) <= 1; flappy_W(28, 518) <= 1; flappy_W(28, 519) <= 1; flappy_W(28, 520) <= 1; flappy_W(28, 521) <= 1; flappy_W(28, 522) <= 1; flappy_W(28, 523) <= 1; flappy_W(28, 524) <= 1; flappy_W(28, 525) <= 1; flappy_W(28, 526) <= 1; flappy_W(28, 527) <= 1; flappy_W(28, 528) <= 1; flappy_W(28, 529) <= 1; flappy_W(28, 530) <= 1; flappy_W(28, 531) <= 1; flappy_W(28, 532) <= 1; flappy_W(28, 533) <= 1; flappy_W(28, 534) <= 1; flappy_W(28, 535) <= 1; flappy_W(28, 536) <= 1; flappy_W(28, 537) <= 1; flappy_W(28, 538) <= 1; flappy_W(28, 539) <= 1; flappy_W(28, 540) <= 0; flappy_W(28, 541) <= 0; flappy_W(28, 542) <= 0; flappy_W(28, 543) <= 0; flappy_W(28, 544) <= 0; flappy_W(28, 545) <= 0; flappy_W(28, 546) <= 0; flappy_W(28, 547) <= 0; flappy_W(28, 548) <= 0; flappy_W(28, 549) <= 0; flappy_W(28, 550) <= 0; flappy_W(28, 551) <= 0; flappy_W(28, 552) <= 0; flappy_W(28, 553) <= 0; flappy_W(28, 554) <= 0; flappy_W(28, 555) <= 0; flappy_W(28, 556) <= 0; flappy_W(28, 557) <= 0; flappy_W(28, 558) <= 0; flappy_W(28, 559) <= 0; flappy_W(28, 560) <= 0; flappy_W(28, 561) <= 0; flappy_W(28, 562) <= 0; flappy_W(28, 563) <= 0; flappy_W(28, 564) <= 1; flappy_W(28, 565) <= 1; flappy_W(28, 566) <= 1; flappy_W(28, 567) <= 1; flappy_W(28, 568) <= 1; flappy_W(28, 569) <= 1; flappy_W(28, 570) <= 1; flappy_W(28, 571) <= 1; flappy_W(28, 572) <= 1; flappy_W(28, 573) <= 1; flappy_W(28, 574) <= 1; flappy_W(28, 575) <= 1; flappy_W(28, 576) <= 0; flappy_W(28, 577) <= 0; flappy_W(28, 578) <= 0; flappy_W(28, 579) <= 0; flappy_W(28, 580) <= 0; flappy_W(28, 581) <= 0; flappy_W(28, 582) <= 0; flappy_W(28, 583) <= 0; flappy_W(28, 584) <= 0; flappy_W(28, 585) <= 0; flappy_W(28, 586) <= 0; flappy_W(28, 587) <= 0; flappy_W(28, 588) <= 1; flappy_W(28, 589) <= 1; flappy_W(28, 590) <= 1; flappy_W(28, 591) <= 1; flappy_W(28, 592) <= 1; flappy_W(28, 593) <= 1; 
flappy_W(29, 0) <= 0; flappy_W(29, 1) <= 0; flappy_W(29, 2) <= 0; flappy_W(29, 3) <= 0; flappy_W(29, 4) <= 0; flappy_W(29, 5) <= 0; flappy_W(29, 6) <= 1; flappy_W(29, 7) <= 1; flappy_W(29, 8) <= 1; flappy_W(29, 9) <= 1; flappy_W(29, 10) <= 1; flappy_W(29, 11) <= 1; flappy_W(29, 12) <= 1; flappy_W(29, 13) <= 1; flappy_W(29, 14) <= 1; flappy_W(29, 15) <= 1; flappy_W(29, 16) <= 1; flappy_W(29, 17) <= 1; flappy_W(29, 18) <= 1; flappy_W(29, 19) <= 1; flappy_W(29, 20) <= 1; flappy_W(29, 21) <= 1; flappy_W(29, 22) <= 1; flappy_W(29, 23) <= 1; flappy_W(29, 24) <= 1; flappy_W(29, 25) <= 1; flappy_W(29, 26) <= 1; flappy_W(29, 27) <= 1; flappy_W(29, 28) <= 1; flappy_W(29, 29) <= 1; flappy_W(29, 30) <= 0; flappy_W(29, 31) <= 0; flappy_W(29, 32) <= 0; flappy_W(29, 33) <= 0; flappy_W(29, 34) <= 0; flappy_W(29, 35) <= 0; flappy_W(29, 36) <= 0; flappy_W(29, 37) <= 0; flappy_W(29, 38) <= 0; flappy_W(29, 39) <= 0; flappy_W(29, 40) <= 0; flappy_W(29, 41) <= 0; flappy_W(29, 42) <= 0; flappy_W(29, 43) <= 0; flappy_W(29, 44) <= 0; flappy_W(29, 45) <= 0; flappy_W(29, 46) <= 0; flappy_W(29, 47) <= 0; flappy_W(29, 48) <= 0; flappy_W(29, 49) <= 0; flappy_W(29, 50) <= 0; flappy_W(29, 51) <= 0; flappy_W(29, 52) <= 0; flappy_W(29, 53) <= 0; flappy_W(29, 54) <= 0; flappy_W(29, 55) <= 0; flappy_W(29, 56) <= 0; flappy_W(29, 57) <= 0; flappy_W(29, 58) <= 0; flappy_W(29, 59) <= 0; flappy_W(29, 60) <= 1; flappy_W(29, 61) <= 1; flappy_W(29, 62) <= 1; flappy_W(29, 63) <= 1; flappy_W(29, 64) <= 1; flappy_W(29, 65) <= 1; flappy_W(29, 66) <= 1; flappy_W(29, 67) <= 1; flappy_W(29, 68) <= 1; flappy_W(29, 69) <= 1; flappy_W(29, 70) <= 1; flappy_W(29, 71) <= 1; flappy_W(29, 72) <= 0; flappy_W(29, 73) <= 0; flappy_W(29, 74) <= 0; flappy_W(29, 75) <= 0; flappy_W(29, 76) <= 0; flappy_W(29, 77) <= 0; flappy_W(29, 78) <= 0; flappy_W(29, 79) <= 0; flappy_W(29, 80) <= 0; flappy_W(29, 81) <= 0; flappy_W(29, 82) <= 0; flappy_W(29, 83) <= 0; flappy_W(29, 84) <= 0; flappy_W(29, 85) <= 0; flappy_W(29, 86) <= 0; flappy_W(29, 87) <= 0; flappy_W(29, 88) <= 0; flappy_W(29, 89) <= 0; flappy_W(29, 90) <= 0; flappy_W(29, 91) <= 0; flappy_W(29, 92) <= 0; flappy_W(29, 93) <= 0; flappy_W(29, 94) <= 0; flappy_W(29, 95) <= 0; flappy_W(29, 96) <= 0; flappy_W(29, 97) <= 0; flappy_W(29, 98) <= 0; flappy_W(29, 99) <= 0; flappy_W(29, 100) <= 0; flappy_W(29, 101) <= 0; flappy_W(29, 102) <= 0; flappy_W(29, 103) <= 0; flappy_W(29, 104) <= 0; flappy_W(29, 105) <= 0; flappy_W(29, 106) <= 0; flappy_W(29, 107) <= 0; flappy_W(29, 108) <= 1; flappy_W(29, 109) <= 1; flappy_W(29, 110) <= 1; flappy_W(29, 111) <= 1; flappy_W(29, 112) <= 1; flappy_W(29, 113) <= 1; flappy_W(29, 114) <= 1; flappy_W(29, 115) <= 1; flappy_W(29, 116) <= 1; flappy_W(29, 117) <= 1; flappy_W(29, 118) <= 1; flappy_W(29, 119) <= 1; flappy_W(29, 120) <= 0; flappy_W(29, 121) <= 0; flappy_W(29, 122) <= 0; flappy_W(29, 123) <= 0; flappy_W(29, 124) <= 0; flappy_W(29, 125) <= 0; flappy_W(29, 126) <= 0; flappy_W(29, 127) <= 0; flappy_W(29, 128) <= 0; flappy_W(29, 129) <= 0; flappy_W(29, 130) <= 0; flappy_W(29, 131) <= 0; flappy_W(29, 132) <= 0; flappy_W(29, 133) <= 0; flappy_W(29, 134) <= 0; flappy_W(29, 135) <= 0; flappy_W(29, 136) <= 0; flappy_W(29, 137) <= 0; flappy_W(29, 138) <= 1; flappy_W(29, 139) <= 1; flappy_W(29, 140) <= 1; flappy_W(29, 141) <= 1; flappy_W(29, 142) <= 1; flappy_W(29, 143) <= 1; flappy_W(29, 144) <= 1; flappy_W(29, 145) <= 1; flappy_W(29, 146) <= 1; flappy_W(29, 147) <= 1; flappy_W(29, 148) <= 1; flappy_W(29, 149) <= 1; flappy_W(29, 150) <= 0; flappy_W(29, 151) <= 0; flappy_W(29, 152) <= 0; flappy_W(29, 153) <= 0; flappy_W(29, 154) <= 0; flappy_W(29, 155) <= 0; flappy_W(29, 156) <= 0; flappy_W(29, 157) <= 0; flappy_W(29, 158) <= 0; flappy_W(29, 159) <= 0; flappy_W(29, 160) <= 0; flappy_W(29, 161) <= 0; flappy_W(29, 162) <= 0; flappy_W(29, 163) <= 0; flappy_W(29, 164) <= 0; flappy_W(29, 165) <= 0; flappy_W(29, 166) <= 0; flappy_W(29, 167) <= 0; flappy_W(29, 168) <= 1; flappy_W(29, 169) <= 1; flappy_W(29, 170) <= 1; flappy_W(29, 171) <= 1; flappy_W(29, 172) <= 1; flappy_W(29, 173) <= 1; flappy_W(29, 174) <= 1; flappy_W(29, 175) <= 1; flappy_W(29, 176) <= 1; flappy_W(29, 177) <= 1; flappy_W(29, 178) <= 1; flappy_W(29, 179) <= 1; flappy_W(29, 180) <= 1; flappy_W(29, 181) <= 1; flappy_W(29, 182) <= 1; flappy_W(29, 183) <= 1; flappy_W(29, 184) <= 1; flappy_W(29, 185) <= 1; flappy_W(29, 186) <= 1; flappy_W(29, 187) <= 1; flappy_W(29, 188) <= 1; flappy_W(29, 189) <= 1; flappy_W(29, 190) <= 1; flappy_W(29, 191) <= 1; flappy_W(29, 192) <= 1; flappy_W(29, 193) <= 1; flappy_W(29, 194) <= 1; flappy_W(29, 195) <= 1; flappy_W(29, 196) <= 1; flappy_W(29, 197) <= 1; flappy_W(29, 198) <= 0; flappy_W(29, 199) <= 0; flappy_W(29, 200) <= 0; flappy_W(29, 201) <= 0; flappy_W(29, 202) <= 0; flappy_W(29, 203) <= 0; flappy_W(29, 204) <= 0; flappy_W(29, 205) <= 0; flappy_W(29, 206) <= 0; flappy_W(29, 207) <= 0; flappy_W(29, 208) <= 0; flappy_W(29, 209) <= 0; flappy_W(29, 210) <= 0; flappy_W(29, 211) <= 0; flappy_W(29, 212) <= 0; flappy_W(29, 213) <= 0; flappy_W(29, 214) <= 0; flappy_W(29, 215) <= 0; flappy_W(29, 216) <= 0; flappy_W(29, 217) <= 0; flappy_W(29, 218) <= 0; flappy_W(29, 219) <= 0; flappy_W(29, 220) <= 0; flappy_W(29, 221) <= 0; flappy_W(29, 222) <= 1; flappy_W(29, 223) <= 1; flappy_W(29, 224) <= 1; flappy_W(29, 225) <= 1; flappy_W(29, 226) <= 1; flappy_W(29, 227) <= 1; flappy_W(29, 228) <= 1; flappy_W(29, 229) <= 1; flappy_W(29, 230) <= 1; flappy_W(29, 231) <= 1; flappy_W(29, 232) <= 1; flappy_W(29, 233) <= 1; flappy_W(29, 234) <= 1; flappy_W(29, 235) <= 1; flappy_W(29, 236) <= 1; flappy_W(29, 237) <= 1; flappy_W(29, 238) <= 1; flappy_W(29, 239) <= 1; flappy_W(29, 240) <= 1; flappy_W(29, 241) <= 1; flappy_W(29, 242) <= 1; flappy_W(29, 243) <= 1; flappy_W(29, 244) <= 1; flappy_W(29, 245) <= 1; flappy_W(29, 246) <= 1; flappy_W(29, 247) <= 1; flappy_W(29, 248) <= 1; flappy_W(29, 249) <= 1; flappy_W(29, 250) <= 1; flappy_W(29, 251) <= 1; flappy_W(29, 252) <= 0; flappy_W(29, 253) <= 0; flappy_W(29, 254) <= 0; flappy_W(29, 255) <= 0; flappy_W(29, 256) <= 0; flappy_W(29, 257) <= 0; flappy_W(29, 258) <= 0; flappy_W(29, 259) <= 0; flappy_W(29, 260) <= 0; flappy_W(29, 261) <= 0; flappy_W(29, 262) <= 0; flappy_W(29, 263) <= 0; flappy_W(29, 264) <= 0; flappy_W(29, 265) <= 0; flappy_W(29, 266) <= 0; flappy_W(29, 267) <= 0; flappy_W(29, 268) <= 0; flappy_W(29, 269) <= 0; flappy_W(29, 270) <= 0; flappy_W(29, 271) <= 0; flappy_W(29, 272) <= 0; flappy_W(29, 273) <= 0; flappy_W(29, 274) <= 0; flappy_W(29, 275) <= 0; flappy_W(29, 276) <= 0; flappy_W(29, 277) <= 0; flappy_W(29, 278) <= 0; flappy_W(29, 279) <= 0; flappy_W(29, 280) <= 0; flappy_W(29, 281) <= 0; flappy_W(29, 282) <= 1; flappy_W(29, 283) <= 1; flappy_W(29, 284) <= 1; flappy_W(29, 285) <= 1; flappy_W(29, 286) <= 1; flappy_W(29, 287) <= 1; flappy_W(29, 288) <= 1; flappy_W(29, 289) <= 1; flappy_W(29, 290) <= 1; flappy_W(29, 291) <= 1; flappy_W(29, 292) <= 1; flappy_W(29, 293) <= 1; flappy_W(29, 294) <= 1; flappy_W(29, 295) <= 1; flappy_W(29, 296) <= 1; flappy_W(29, 297) <= 1; flappy_W(29, 298) <= 1; flappy_W(29, 299) <= 1; flappy_W(29, 300) <= 1; flappy_W(29, 301) <= 1; flappy_W(29, 302) <= 1; flappy_W(29, 303) <= 1; flappy_W(29, 304) <= 1; flappy_W(29, 305) <= 1; flappy_W(29, 306) <= 0; flappy_W(29, 307) <= 0; flappy_W(29, 308) <= 0; flappy_W(29, 309) <= 0; flappy_W(29, 310) <= 0; flappy_W(29, 311) <= 0; flappy_W(29, 312) <= 0; flappy_W(29, 313) <= 0; flappy_W(29, 314) <= 0; flappy_W(29, 315) <= 0; flappy_W(29, 316) <= 0; flappy_W(29, 317) <= 0; flappy_W(29, 318) <= 0; flappy_W(29, 319) <= 0; flappy_W(29, 320) <= 0; flappy_W(29, 321) <= 0; flappy_W(29, 322) <= 0; flappy_W(29, 323) <= 0; flappy_W(29, 324) <= 0; flappy_W(29, 325) <= 0; flappy_W(29, 326) <= 0; flappy_W(29, 327) <= 0; flappy_W(29, 328) <= 0; flappy_W(29, 329) <= 0; flappy_W(29, 330) <= 0; flappy_W(29, 331) <= 0; flappy_W(29, 332) <= 0; flappy_W(29, 333) <= 0; flappy_W(29, 334) <= 0; flappy_W(29, 335) <= 0; flappy_W(29, 336) <= 0; flappy_W(29, 337) <= 0; flappy_W(29, 338) <= 0; flappy_W(29, 339) <= 0; flappy_W(29, 340) <= 0; flappy_W(29, 341) <= 0; flappy_W(29, 342) <= 0; flappy_W(29, 343) <= 0; flappy_W(29, 344) <= 0; flappy_W(29, 345) <= 0; flappy_W(29, 346) <= 0; flappy_W(29, 347) <= 0; flappy_W(29, 348) <= 0; flappy_W(29, 349) <= 0; flappy_W(29, 350) <= 0; flappy_W(29, 351) <= 0; flappy_W(29, 352) <= 0; flappy_W(29, 353) <= 0; flappy_W(29, 354) <= 0; flappy_W(29, 355) <= 0; flappy_W(29, 356) <= 0; flappy_W(29, 357) <= 0; flappy_W(29, 358) <= 0; flappy_W(29, 359) <= 0; flappy_W(29, 360) <= 0; flappy_W(29, 361) <= 0; flappy_W(29, 362) <= 0; flappy_W(29, 363) <= 0; flappy_W(29, 364) <= 0; flappy_W(29, 365) <= 0; flappy_W(29, 366) <= 0; flappy_W(29, 367) <= 0; flappy_W(29, 368) <= 0; flappy_W(29, 369) <= 0; flappy_W(29, 370) <= 0; flappy_W(29, 371) <= 0; flappy_W(29, 372) <= 0; flappy_W(29, 373) <= 0; flappy_W(29, 374) <= 0; flappy_W(29, 375) <= 0; flappy_W(29, 376) <= 0; flappy_W(29, 377) <= 0; flappy_W(29, 378) <= 0; flappy_W(29, 379) <= 0; flappy_W(29, 380) <= 0; flappy_W(29, 381) <= 0; flappy_W(29, 382) <= 0; flappy_W(29, 383) <= 0; flappy_W(29, 384) <= 0; flappy_W(29, 385) <= 0; flappy_W(29, 386) <= 0; flappy_W(29, 387) <= 0; flappy_W(29, 388) <= 0; flappy_W(29, 389) <= 0; flappy_W(29, 390) <= 0; flappy_W(29, 391) <= 0; flappy_W(29, 392) <= 0; flappy_W(29, 393) <= 0; flappy_W(29, 394) <= 0; flappy_W(29, 395) <= 0; flappy_W(29, 396) <= 0; flappy_W(29, 397) <= 0; flappy_W(29, 398) <= 0; flappy_W(29, 399) <= 0; flappy_W(29, 400) <= 0; flappy_W(29, 401) <= 0; flappy_W(29, 402) <= 1; flappy_W(29, 403) <= 1; flappy_W(29, 404) <= 1; flappy_W(29, 405) <= 1; flappy_W(29, 406) <= 1; flappy_W(29, 407) <= 1; flappy_W(29, 408) <= 1; flappy_W(29, 409) <= 1; flappy_W(29, 410) <= 1; flappy_W(29, 411) <= 1; flappy_W(29, 412) <= 1; flappy_W(29, 413) <= 1; flappy_W(29, 414) <= 1; flappy_W(29, 415) <= 1; flappy_W(29, 416) <= 1; flappy_W(29, 417) <= 1; flappy_W(29, 418) <= 1; flappy_W(29, 419) <= 1; flappy_W(29, 420) <= 1; flappy_W(29, 421) <= 1; flappy_W(29, 422) <= 1; flappy_W(29, 423) <= 1; flappy_W(29, 424) <= 1; flappy_W(29, 425) <= 1; flappy_W(29, 426) <= 1; flappy_W(29, 427) <= 1; flappy_W(29, 428) <= 1; flappy_W(29, 429) <= 1; flappy_W(29, 430) <= 1; flappy_W(29, 431) <= 1; flappy_W(29, 432) <= 0; flappy_W(29, 433) <= 0; flappy_W(29, 434) <= 0; flappy_W(29, 435) <= 0; flappy_W(29, 436) <= 0; flappy_W(29, 437) <= 0; flappy_W(29, 438) <= 0; flappy_W(29, 439) <= 0; flappy_W(29, 440) <= 0; flappy_W(29, 441) <= 0; flappy_W(29, 442) <= 0; flappy_W(29, 443) <= 0; flappy_W(29, 444) <= 0; flappy_W(29, 445) <= 0; flappy_W(29, 446) <= 0; flappy_W(29, 447) <= 0; flappy_W(29, 448) <= 0; flappy_W(29, 449) <= 0; flappy_W(29, 450) <= 0; flappy_W(29, 451) <= 0; flappy_W(29, 452) <= 0; flappy_W(29, 453) <= 0; flappy_W(29, 454) <= 0; flappy_W(29, 455) <= 0; flappy_W(29, 456) <= 0; flappy_W(29, 457) <= 0; flappy_W(29, 458) <= 0; flappy_W(29, 459) <= 0; flappy_W(29, 460) <= 0; flappy_W(29, 461) <= 0; flappy_W(29, 462) <= 0; flappy_W(29, 463) <= 0; flappy_W(29, 464) <= 0; flappy_W(29, 465) <= 0; flappy_W(29, 466) <= 0; flappy_W(29, 467) <= 0; flappy_W(29, 468) <= 1; flappy_W(29, 469) <= 1; flappy_W(29, 470) <= 1; flappy_W(29, 471) <= 1; flappy_W(29, 472) <= 1; flappy_W(29, 473) <= 1; flappy_W(29, 474) <= 1; flappy_W(29, 475) <= 1; flappy_W(29, 476) <= 1; flappy_W(29, 477) <= 1; flappy_W(29, 478) <= 1; flappy_W(29, 479) <= 1; flappy_W(29, 480) <= 0; flappy_W(29, 481) <= 0; flappy_W(29, 482) <= 0; flappy_W(29, 483) <= 0; flappy_W(29, 484) <= 0; flappy_W(29, 485) <= 0; flappy_W(29, 486) <= 0; flappy_W(29, 487) <= 0; flappy_W(29, 488) <= 0; flappy_W(29, 489) <= 0; flappy_W(29, 490) <= 0; flappy_W(29, 491) <= 0; flappy_W(29, 492) <= 0; flappy_W(29, 493) <= 0; flappy_W(29, 494) <= 0; flappy_W(29, 495) <= 0; flappy_W(29, 496) <= 0; flappy_W(29, 497) <= 0; flappy_W(29, 498) <= 0; flappy_W(29, 499) <= 0; flappy_W(29, 500) <= 0; flappy_W(29, 501) <= 0; flappy_W(29, 502) <= 0; flappy_W(29, 503) <= 0; flappy_W(29, 504) <= 0; flappy_W(29, 505) <= 0; flappy_W(29, 506) <= 0; flappy_W(29, 507) <= 0; flappy_W(29, 508) <= 0; flappy_W(29, 509) <= 0; flappy_W(29, 510) <= 1; flappy_W(29, 511) <= 1; flappy_W(29, 512) <= 1; flappy_W(29, 513) <= 1; flappy_W(29, 514) <= 1; flappy_W(29, 515) <= 1; flappy_W(29, 516) <= 1; flappy_W(29, 517) <= 1; flappy_W(29, 518) <= 1; flappy_W(29, 519) <= 1; flappy_W(29, 520) <= 1; flappy_W(29, 521) <= 1; flappy_W(29, 522) <= 1; flappy_W(29, 523) <= 1; flappy_W(29, 524) <= 1; flappy_W(29, 525) <= 1; flappy_W(29, 526) <= 1; flappy_W(29, 527) <= 1; flappy_W(29, 528) <= 1; flappy_W(29, 529) <= 1; flappy_W(29, 530) <= 1; flappy_W(29, 531) <= 1; flappy_W(29, 532) <= 1; flappy_W(29, 533) <= 1; flappy_W(29, 534) <= 1; flappy_W(29, 535) <= 1; flappy_W(29, 536) <= 1; flappy_W(29, 537) <= 1; flappy_W(29, 538) <= 1; flappy_W(29, 539) <= 1; flappy_W(29, 540) <= 0; flappy_W(29, 541) <= 0; flappy_W(29, 542) <= 0; flappy_W(29, 543) <= 0; flappy_W(29, 544) <= 0; flappy_W(29, 545) <= 0; flappy_W(29, 546) <= 0; flappy_W(29, 547) <= 0; flappy_W(29, 548) <= 0; flappy_W(29, 549) <= 0; flappy_W(29, 550) <= 0; flappy_W(29, 551) <= 0; flappy_W(29, 552) <= 0; flappy_W(29, 553) <= 0; flappy_W(29, 554) <= 0; flappy_W(29, 555) <= 0; flappy_W(29, 556) <= 0; flappy_W(29, 557) <= 0; flappy_W(29, 558) <= 0; flappy_W(29, 559) <= 0; flappy_W(29, 560) <= 0; flappy_W(29, 561) <= 0; flappy_W(29, 562) <= 0; flappy_W(29, 563) <= 0; flappy_W(29, 564) <= 1; flappy_W(29, 565) <= 1; flappy_W(29, 566) <= 1; flappy_W(29, 567) <= 1; flappy_W(29, 568) <= 1; flappy_W(29, 569) <= 1; flappy_W(29, 570) <= 1; flappy_W(29, 571) <= 1; flappy_W(29, 572) <= 1; flappy_W(29, 573) <= 1; flappy_W(29, 574) <= 1; flappy_W(29, 575) <= 1; flappy_W(29, 576) <= 0; flappy_W(29, 577) <= 0; flappy_W(29, 578) <= 0; flappy_W(29, 579) <= 0; flappy_W(29, 580) <= 0; flappy_W(29, 581) <= 0; flappy_W(29, 582) <= 0; flappy_W(29, 583) <= 0; flappy_W(29, 584) <= 0; flappy_W(29, 585) <= 0; flappy_W(29, 586) <= 0; flappy_W(29, 587) <= 0; flappy_W(29, 588) <= 1; flappy_W(29, 589) <= 1; flappy_W(29, 590) <= 1; flappy_W(29, 591) <= 1; flappy_W(29, 592) <= 1; flappy_W(29, 593) <= 1; 
flappy_W(30, 0) <= 0; flappy_W(30, 1) <= 0; flappy_W(30, 2) <= 0; flappy_W(30, 3) <= 0; flappy_W(30, 4) <= 0; flappy_W(30, 5) <= 0; flappy_W(30, 6) <= 1; flappy_W(30, 7) <= 1; flappy_W(30, 8) <= 1; flappy_W(30, 9) <= 1; flappy_W(30, 10) <= 1; flappy_W(30, 11) <= 1; flappy_W(30, 12) <= 1; flappy_W(30, 13) <= 1; flappy_W(30, 14) <= 1; flappy_W(30, 15) <= 1; flappy_W(30, 16) <= 1; flappy_W(30, 17) <= 1; flappy_W(30, 18) <= 0; flappy_W(30, 19) <= 0; flappy_W(30, 20) <= 0; flappy_W(30, 21) <= 0; flappy_W(30, 22) <= 0; flappy_W(30, 23) <= 0; flappy_W(30, 24) <= 1; flappy_W(30, 25) <= 1; flappy_W(30, 26) <= 1; flappy_W(30, 27) <= 1; flappy_W(30, 28) <= 1; flappy_W(30, 29) <= 1; flappy_W(30, 30) <= 0; flappy_W(30, 31) <= 0; flappy_W(30, 32) <= 0; flappy_W(30, 33) <= 0; flappy_W(30, 34) <= 0; flappy_W(30, 35) <= 0; flappy_W(30, 36) <= 0; flappy_W(30, 37) <= 0; flappy_W(30, 38) <= 0; flappy_W(30, 39) <= 0; flappy_W(30, 40) <= 0; flappy_W(30, 41) <= 0; flappy_W(30, 42) <= 0; flappy_W(30, 43) <= 0; flappy_W(30, 44) <= 0; flappy_W(30, 45) <= 0; flappy_W(30, 46) <= 0; flappy_W(30, 47) <= 0; flappy_W(30, 48) <= 0; flappy_W(30, 49) <= 0; flappy_W(30, 50) <= 0; flappy_W(30, 51) <= 0; flappy_W(30, 52) <= 0; flappy_W(30, 53) <= 0; flappy_W(30, 54) <= 0; flappy_W(30, 55) <= 0; flappy_W(30, 56) <= 0; flappy_W(30, 57) <= 0; flappy_W(30, 58) <= 0; flappy_W(30, 59) <= 0; flappy_W(30, 60) <= 1; flappy_W(30, 61) <= 1; flappy_W(30, 62) <= 1; flappy_W(30, 63) <= 1; flappy_W(30, 64) <= 1; flappy_W(30, 65) <= 1; flappy_W(30, 66) <= 1; flappy_W(30, 67) <= 1; flappy_W(30, 68) <= 1; flappy_W(30, 69) <= 1; flappy_W(30, 70) <= 1; flappy_W(30, 71) <= 1; flappy_W(30, 72) <= 0; flappy_W(30, 73) <= 0; flappy_W(30, 74) <= 0; flappy_W(30, 75) <= 0; flappy_W(30, 76) <= 0; flappy_W(30, 77) <= 0; flappy_W(30, 78) <= 0; flappy_W(30, 79) <= 0; flappy_W(30, 80) <= 0; flappy_W(30, 81) <= 0; flappy_W(30, 82) <= 0; flappy_W(30, 83) <= 0; flappy_W(30, 84) <= 0; flappy_W(30, 85) <= 0; flappy_W(30, 86) <= 0; flappy_W(30, 87) <= 0; flappy_W(30, 88) <= 0; flappy_W(30, 89) <= 0; flappy_W(30, 90) <= 0; flappy_W(30, 91) <= 0; flappy_W(30, 92) <= 0; flappy_W(30, 93) <= 0; flappy_W(30, 94) <= 0; flappy_W(30, 95) <= 0; flappy_W(30, 96) <= 0; flappy_W(30, 97) <= 0; flappy_W(30, 98) <= 0; flappy_W(30, 99) <= 0; flappy_W(30, 100) <= 0; flappy_W(30, 101) <= 0; flappy_W(30, 102) <= 0; flappy_W(30, 103) <= 0; flappy_W(30, 104) <= 0; flappy_W(30, 105) <= 0; flappy_W(30, 106) <= 0; flappy_W(30, 107) <= 0; flappy_W(30, 108) <= 1; flappy_W(30, 109) <= 1; flappy_W(30, 110) <= 1; flappy_W(30, 111) <= 1; flappy_W(30, 112) <= 1; flappy_W(30, 113) <= 1; flappy_W(30, 114) <= 1; flappy_W(30, 115) <= 1; flappy_W(30, 116) <= 1; flappy_W(30, 117) <= 1; flappy_W(30, 118) <= 1; flappy_W(30, 119) <= 1; flappy_W(30, 120) <= 1; flappy_W(30, 121) <= 1; flappy_W(30, 122) <= 1; flappy_W(30, 123) <= 1; flappy_W(30, 124) <= 1; flappy_W(30, 125) <= 1; flappy_W(30, 126) <= 1; flappy_W(30, 127) <= 1; flappy_W(30, 128) <= 1; flappy_W(30, 129) <= 1; flappy_W(30, 130) <= 1; flappy_W(30, 131) <= 1; flappy_W(30, 132) <= 1; flappy_W(30, 133) <= 1; flappy_W(30, 134) <= 1; flappy_W(30, 135) <= 1; flappy_W(30, 136) <= 1; flappy_W(30, 137) <= 1; flappy_W(30, 138) <= 1; flappy_W(30, 139) <= 1; flappy_W(30, 140) <= 1; flappy_W(30, 141) <= 1; flappy_W(30, 142) <= 1; flappy_W(30, 143) <= 1; flappy_W(30, 144) <= 1; flappy_W(30, 145) <= 1; flappy_W(30, 146) <= 1; flappy_W(30, 147) <= 1; flappy_W(30, 148) <= 1; flappy_W(30, 149) <= 1; flappy_W(30, 150) <= 0; flappy_W(30, 151) <= 0; flappy_W(30, 152) <= 0; flappy_W(30, 153) <= 0; flappy_W(30, 154) <= 0; flappy_W(30, 155) <= 0; flappy_W(30, 156) <= 0; flappy_W(30, 157) <= 0; flappy_W(30, 158) <= 0; flappy_W(30, 159) <= 0; flappy_W(30, 160) <= 0; flappy_W(30, 161) <= 0; flappy_W(30, 162) <= 0; flappy_W(30, 163) <= 0; flappy_W(30, 164) <= 0; flappy_W(30, 165) <= 0; flappy_W(30, 166) <= 0; flappy_W(30, 167) <= 0; flappy_W(30, 168) <= 1; flappy_W(30, 169) <= 1; flappy_W(30, 170) <= 1; flappy_W(30, 171) <= 1; flappy_W(30, 172) <= 1; flappy_W(30, 173) <= 1; flappy_W(30, 174) <= 1; flappy_W(30, 175) <= 1; flappy_W(30, 176) <= 1; flappy_W(30, 177) <= 1; flappy_W(30, 178) <= 1; flappy_W(30, 179) <= 1; flappy_W(30, 180) <= 0; flappy_W(30, 181) <= 0; flappy_W(30, 182) <= 0; flappy_W(30, 183) <= 0; flappy_W(30, 184) <= 0; flappy_W(30, 185) <= 0; flappy_W(30, 186) <= 0; flappy_W(30, 187) <= 0; flappy_W(30, 188) <= 0; flappy_W(30, 189) <= 0; flappy_W(30, 190) <= 0; flappy_W(30, 191) <= 0; flappy_W(30, 192) <= 0; flappy_W(30, 193) <= 0; flappy_W(30, 194) <= 0; flappy_W(30, 195) <= 0; flappy_W(30, 196) <= 0; flappy_W(30, 197) <= 0; flappy_W(30, 198) <= 0; flappy_W(30, 199) <= 0; flappy_W(30, 200) <= 0; flappy_W(30, 201) <= 0; flappy_W(30, 202) <= 0; flappy_W(30, 203) <= 0; flappy_W(30, 204) <= 0; flappy_W(30, 205) <= 0; flappy_W(30, 206) <= 0; flappy_W(30, 207) <= 0; flappy_W(30, 208) <= 0; flappy_W(30, 209) <= 0; flappy_W(30, 210) <= 0; flappy_W(30, 211) <= 0; flappy_W(30, 212) <= 0; flappy_W(30, 213) <= 0; flappy_W(30, 214) <= 0; flappy_W(30, 215) <= 0; flappy_W(30, 216) <= 0; flappy_W(30, 217) <= 0; flappy_W(30, 218) <= 0; flappy_W(30, 219) <= 0; flappy_W(30, 220) <= 0; flappy_W(30, 221) <= 0; flappy_W(30, 222) <= 1; flappy_W(30, 223) <= 1; flappy_W(30, 224) <= 1; flappy_W(30, 225) <= 1; flappy_W(30, 226) <= 1; flappy_W(30, 227) <= 1; flappy_W(30, 228) <= 1; flappy_W(30, 229) <= 1; flappy_W(30, 230) <= 1; flappy_W(30, 231) <= 1; flappy_W(30, 232) <= 1; flappy_W(30, 233) <= 1; flappy_W(30, 234) <= 0; flappy_W(30, 235) <= 0; flappy_W(30, 236) <= 0; flappy_W(30, 237) <= 0; flappy_W(30, 238) <= 0; flappy_W(30, 239) <= 0; flappy_W(30, 240) <= 0; flappy_W(30, 241) <= 0; flappy_W(30, 242) <= 0; flappy_W(30, 243) <= 0; flappy_W(30, 244) <= 0; flappy_W(30, 245) <= 0; flappy_W(30, 246) <= 0; flappy_W(30, 247) <= 0; flappy_W(30, 248) <= 0; flappy_W(30, 249) <= 0; flappy_W(30, 250) <= 0; flappy_W(30, 251) <= 0; flappy_W(30, 252) <= 0; flappy_W(30, 253) <= 0; flappy_W(30, 254) <= 0; flappy_W(30, 255) <= 0; flappy_W(30, 256) <= 0; flappy_W(30, 257) <= 0; flappy_W(30, 258) <= 0; flappy_W(30, 259) <= 0; flappy_W(30, 260) <= 0; flappy_W(30, 261) <= 0; flappy_W(30, 262) <= 0; flappy_W(30, 263) <= 0; flappy_W(30, 264) <= 0; flappy_W(30, 265) <= 0; flappy_W(30, 266) <= 0; flappy_W(30, 267) <= 0; flappy_W(30, 268) <= 0; flappy_W(30, 269) <= 0; flappy_W(30, 270) <= 0; flappy_W(30, 271) <= 0; flappy_W(30, 272) <= 0; flappy_W(30, 273) <= 0; flappy_W(30, 274) <= 0; flappy_W(30, 275) <= 0; flappy_W(30, 276) <= 0; flappy_W(30, 277) <= 0; flappy_W(30, 278) <= 0; flappy_W(30, 279) <= 0; flappy_W(30, 280) <= 0; flappy_W(30, 281) <= 0; flappy_W(30, 282) <= 0; flappy_W(30, 283) <= 0; flappy_W(30, 284) <= 0; flappy_W(30, 285) <= 0; flappy_W(30, 286) <= 0; flappy_W(30, 287) <= 0; flappy_W(30, 288) <= 1; flappy_W(30, 289) <= 1; flappy_W(30, 290) <= 1; flappy_W(30, 291) <= 1; flappy_W(30, 292) <= 1; flappy_W(30, 293) <= 1; flappy_W(30, 294) <= 1; flappy_W(30, 295) <= 1; flappy_W(30, 296) <= 1; flappy_W(30, 297) <= 1; flappy_W(30, 298) <= 1; flappy_W(30, 299) <= 1; flappy_W(30, 300) <= 0; flappy_W(30, 301) <= 0; flappy_W(30, 302) <= 0; flappy_W(30, 303) <= 0; flappy_W(30, 304) <= 0; flappy_W(30, 305) <= 0; flappy_W(30, 306) <= 0; flappy_W(30, 307) <= 0; flappy_W(30, 308) <= 0; flappy_W(30, 309) <= 0; flappy_W(30, 310) <= 0; flappy_W(30, 311) <= 0; flappy_W(30, 312) <= 0; flappy_W(30, 313) <= 0; flappy_W(30, 314) <= 0; flappy_W(30, 315) <= 0; flappy_W(30, 316) <= 0; flappy_W(30, 317) <= 0; flappy_W(30, 318) <= 0; flappy_W(30, 319) <= 0; flappy_W(30, 320) <= 0; flappy_W(30, 321) <= 0; flappy_W(30, 322) <= 0; flappy_W(30, 323) <= 0; flappy_W(30, 324) <= 0; flappy_W(30, 325) <= 0; flappy_W(30, 326) <= 0; flappy_W(30, 327) <= 0; flappy_W(30, 328) <= 0; flappy_W(30, 329) <= 0; flappy_W(30, 330) <= 0; flappy_W(30, 331) <= 0; flappy_W(30, 332) <= 0; flappy_W(30, 333) <= 0; flappy_W(30, 334) <= 0; flappy_W(30, 335) <= 0; flappy_W(30, 336) <= 0; flappy_W(30, 337) <= 0; flappy_W(30, 338) <= 0; flappy_W(30, 339) <= 0; flappy_W(30, 340) <= 0; flappy_W(30, 341) <= 0; flappy_W(30, 342) <= 0; flappy_W(30, 343) <= 0; flappy_W(30, 344) <= 0; flappy_W(30, 345) <= 0; flappy_W(30, 346) <= 0; flappy_W(30, 347) <= 0; flappy_W(30, 348) <= 0; flappy_W(30, 349) <= 0; flappy_W(30, 350) <= 0; flappy_W(30, 351) <= 0; flappy_W(30, 352) <= 0; flappy_W(30, 353) <= 0; flappy_W(30, 354) <= 0; flappy_W(30, 355) <= 0; flappy_W(30, 356) <= 0; flappy_W(30, 357) <= 0; flappy_W(30, 358) <= 0; flappy_W(30, 359) <= 0; flappy_W(30, 360) <= 0; flappy_W(30, 361) <= 0; flappy_W(30, 362) <= 0; flappy_W(30, 363) <= 0; flappy_W(30, 364) <= 0; flappy_W(30, 365) <= 0; flappy_W(30, 366) <= 0; flappy_W(30, 367) <= 0; flappy_W(30, 368) <= 0; flappy_W(30, 369) <= 0; flappy_W(30, 370) <= 0; flappy_W(30, 371) <= 0; flappy_W(30, 372) <= 0; flappy_W(30, 373) <= 0; flappy_W(30, 374) <= 0; flappy_W(30, 375) <= 0; flappy_W(30, 376) <= 0; flappy_W(30, 377) <= 0; flappy_W(30, 378) <= 0; flappy_W(30, 379) <= 0; flappy_W(30, 380) <= 0; flappy_W(30, 381) <= 0; flappy_W(30, 382) <= 0; flappy_W(30, 383) <= 0; flappy_W(30, 384) <= 0; flappy_W(30, 385) <= 0; flappy_W(30, 386) <= 0; flappy_W(30, 387) <= 0; flappy_W(30, 388) <= 0; flappy_W(30, 389) <= 0; flappy_W(30, 390) <= 0; flappy_W(30, 391) <= 0; flappy_W(30, 392) <= 0; flappy_W(30, 393) <= 0; flappy_W(30, 394) <= 0; flappy_W(30, 395) <= 0; flappy_W(30, 396) <= 0; flappy_W(30, 397) <= 0; flappy_W(30, 398) <= 0; flappy_W(30, 399) <= 0; flappy_W(30, 400) <= 0; flappy_W(30, 401) <= 0; flappy_W(30, 402) <= 1; flappy_W(30, 403) <= 1; flappy_W(30, 404) <= 1; flappy_W(30, 405) <= 1; flappy_W(30, 406) <= 1; flappy_W(30, 407) <= 1; flappy_W(30, 408) <= 1; flappy_W(30, 409) <= 1; flappy_W(30, 410) <= 1; flappy_W(30, 411) <= 1; flappy_W(30, 412) <= 1; flappy_W(30, 413) <= 1; flappy_W(30, 414) <= 0; flappy_W(30, 415) <= 0; flappy_W(30, 416) <= 0; flappy_W(30, 417) <= 0; flappy_W(30, 418) <= 0; flappy_W(30, 419) <= 0; flappy_W(30, 420) <= 0; flappy_W(30, 421) <= 0; flappy_W(30, 422) <= 0; flappy_W(30, 423) <= 0; flappy_W(30, 424) <= 0; flappy_W(30, 425) <= 0; flappy_W(30, 426) <= 1; flappy_W(30, 427) <= 1; flappy_W(30, 428) <= 1; flappy_W(30, 429) <= 1; flappy_W(30, 430) <= 1; flappy_W(30, 431) <= 1; flappy_W(30, 432) <= 1; flappy_W(30, 433) <= 1; flappy_W(30, 434) <= 1; flappy_W(30, 435) <= 1; flappy_W(30, 436) <= 1; flappy_W(30, 437) <= 1; flappy_W(30, 438) <= 0; flappy_W(30, 439) <= 0; flappy_W(30, 440) <= 0; flappy_W(30, 441) <= 0; flappy_W(30, 442) <= 0; flappy_W(30, 443) <= 0; flappy_W(30, 444) <= 0; flappy_W(30, 445) <= 0; flappy_W(30, 446) <= 0; flappy_W(30, 447) <= 0; flappy_W(30, 448) <= 0; flappy_W(30, 449) <= 0; flappy_W(30, 450) <= 0; flappy_W(30, 451) <= 0; flappy_W(30, 452) <= 0; flappy_W(30, 453) <= 0; flappy_W(30, 454) <= 0; flappy_W(30, 455) <= 0; flappy_W(30, 456) <= 0; flappy_W(30, 457) <= 0; flappy_W(30, 458) <= 0; flappy_W(30, 459) <= 0; flappy_W(30, 460) <= 0; flappy_W(30, 461) <= 0; flappy_W(30, 462) <= 0; flappy_W(30, 463) <= 0; flappy_W(30, 464) <= 0; flappy_W(30, 465) <= 0; flappy_W(30, 466) <= 0; flappy_W(30, 467) <= 0; flappy_W(30, 468) <= 1; flappy_W(30, 469) <= 1; flappy_W(30, 470) <= 1; flappy_W(30, 471) <= 1; flappy_W(30, 472) <= 1; flappy_W(30, 473) <= 1; flappy_W(30, 474) <= 1; flappy_W(30, 475) <= 1; flappy_W(30, 476) <= 1; flappy_W(30, 477) <= 1; flappy_W(30, 478) <= 1; flappy_W(30, 479) <= 1; flappy_W(30, 480) <= 0; flappy_W(30, 481) <= 0; flappy_W(30, 482) <= 0; flappy_W(30, 483) <= 0; flappy_W(30, 484) <= 0; flappy_W(30, 485) <= 0; flappy_W(30, 486) <= 0; flappy_W(30, 487) <= 0; flappy_W(30, 488) <= 0; flappy_W(30, 489) <= 0; flappy_W(30, 490) <= 0; flappy_W(30, 491) <= 0; flappy_W(30, 492) <= 0; flappy_W(30, 493) <= 0; flappy_W(30, 494) <= 0; flappy_W(30, 495) <= 0; flappy_W(30, 496) <= 0; flappy_W(30, 497) <= 0; flappy_W(30, 498) <= 0; flappy_W(30, 499) <= 0; flappy_W(30, 500) <= 0; flappy_W(30, 501) <= 0; flappy_W(30, 502) <= 0; flappy_W(30, 503) <= 0; flappy_W(30, 504) <= 0; flappy_W(30, 505) <= 0; flappy_W(30, 506) <= 0; flappy_W(30, 507) <= 0; flappy_W(30, 508) <= 0; flappy_W(30, 509) <= 0; flappy_W(30, 510) <= 1; flappy_W(30, 511) <= 1; flappy_W(30, 512) <= 1; flappy_W(30, 513) <= 1; flappy_W(30, 514) <= 1; flappy_W(30, 515) <= 1; flappy_W(30, 516) <= 1; flappy_W(30, 517) <= 1; flappy_W(30, 518) <= 1; flappy_W(30, 519) <= 1; flappy_W(30, 520) <= 1; flappy_W(30, 521) <= 1; flappy_W(30, 522) <= 0; flappy_W(30, 523) <= 0; flappy_W(30, 524) <= 0; flappy_W(30, 525) <= 0; flappy_W(30, 526) <= 0; flappy_W(30, 527) <= 0; flappy_W(30, 528) <= 1; flappy_W(30, 529) <= 1; flappy_W(30, 530) <= 1; flappy_W(30, 531) <= 1; flappy_W(30, 532) <= 1; flappy_W(30, 533) <= 1; flappy_W(30, 534) <= 1; flappy_W(30, 535) <= 1; flappy_W(30, 536) <= 1; flappy_W(30, 537) <= 1; flappy_W(30, 538) <= 1; flappy_W(30, 539) <= 1; flappy_W(30, 540) <= 0; flappy_W(30, 541) <= 0; flappy_W(30, 542) <= 0; flappy_W(30, 543) <= 0; flappy_W(30, 544) <= 0; flappy_W(30, 545) <= 0; flappy_W(30, 546) <= 0; flappy_W(30, 547) <= 0; flappy_W(30, 548) <= 0; flappy_W(30, 549) <= 0; flappy_W(30, 550) <= 0; flappy_W(30, 551) <= 0; flappy_W(30, 552) <= 0; flappy_W(30, 553) <= 0; flappy_W(30, 554) <= 0; flappy_W(30, 555) <= 0; flappy_W(30, 556) <= 0; flappy_W(30, 557) <= 0; flappy_W(30, 558) <= 0; flappy_W(30, 559) <= 0; flappy_W(30, 560) <= 0; flappy_W(30, 561) <= 0; flappy_W(30, 562) <= 0; flappy_W(30, 563) <= 0; flappy_W(30, 564) <= 1; flappy_W(30, 565) <= 1; flappy_W(30, 566) <= 1; flappy_W(30, 567) <= 1; flappy_W(30, 568) <= 1; flappy_W(30, 569) <= 1; flappy_W(30, 570) <= 1; flappy_W(30, 571) <= 1; flappy_W(30, 572) <= 1; flappy_W(30, 573) <= 1; flappy_W(30, 574) <= 1; flappy_W(30, 575) <= 1; flappy_W(30, 576) <= 0; flappy_W(30, 577) <= 0; flappy_W(30, 578) <= 0; flappy_W(30, 579) <= 0; flappy_W(30, 580) <= 0; flappy_W(30, 581) <= 0; flappy_W(30, 582) <= 0; flappy_W(30, 583) <= 0; flappy_W(30, 584) <= 0; flappy_W(30, 585) <= 0; flappy_W(30, 586) <= 0; flappy_W(30, 587) <= 0; flappy_W(30, 588) <= 1; flappy_W(30, 589) <= 1; flappy_W(30, 590) <= 1; flappy_W(30, 591) <= 1; flappy_W(30, 592) <= 1; flappy_W(30, 593) <= 1; 
flappy_W(31, 0) <= 0; flappy_W(31, 1) <= 0; flappy_W(31, 2) <= 0; flappy_W(31, 3) <= 0; flappy_W(31, 4) <= 0; flappy_W(31, 5) <= 0; flappy_W(31, 6) <= 1; flappy_W(31, 7) <= 1; flappy_W(31, 8) <= 1; flappy_W(31, 9) <= 1; flappy_W(31, 10) <= 1; flappy_W(31, 11) <= 1; flappy_W(31, 12) <= 1; flappy_W(31, 13) <= 1; flappy_W(31, 14) <= 1; flappy_W(31, 15) <= 1; flappy_W(31, 16) <= 1; flappy_W(31, 17) <= 1; flappy_W(31, 18) <= 0; flappy_W(31, 19) <= 0; flappy_W(31, 20) <= 0; flappy_W(31, 21) <= 0; flappy_W(31, 22) <= 0; flappy_W(31, 23) <= 0; flappy_W(31, 24) <= 1; flappy_W(31, 25) <= 1; flappy_W(31, 26) <= 1; flappy_W(31, 27) <= 1; flappy_W(31, 28) <= 1; flappy_W(31, 29) <= 1; flappy_W(31, 30) <= 0; flappy_W(31, 31) <= 0; flappy_W(31, 32) <= 0; flappy_W(31, 33) <= 0; flappy_W(31, 34) <= 0; flappy_W(31, 35) <= 0; flappy_W(31, 36) <= 0; flappy_W(31, 37) <= 0; flappy_W(31, 38) <= 0; flappy_W(31, 39) <= 0; flappy_W(31, 40) <= 0; flappy_W(31, 41) <= 0; flappy_W(31, 42) <= 0; flappy_W(31, 43) <= 0; flappy_W(31, 44) <= 0; flappy_W(31, 45) <= 0; flappy_W(31, 46) <= 0; flappy_W(31, 47) <= 0; flappy_W(31, 48) <= 0; flappy_W(31, 49) <= 0; flappy_W(31, 50) <= 0; flappy_W(31, 51) <= 0; flappy_W(31, 52) <= 0; flappy_W(31, 53) <= 0; flappy_W(31, 54) <= 0; flappy_W(31, 55) <= 0; flappy_W(31, 56) <= 0; flappy_W(31, 57) <= 0; flappy_W(31, 58) <= 0; flappy_W(31, 59) <= 0; flappy_W(31, 60) <= 1; flappy_W(31, 61) <= 1; flappy_W(31, 62) <= 1; flappy_W(31, 63) <= 1; flappy_W(31, 64) <= 1; flappy_W(31, 65) <= 1; flappy_W(31, 66) <= 1; flappy_W(31, 67) <= 1; flappy_W(31, 68) <= 1; flappy_W(31, 69) <= 1; flappy_W(31, 70) <= 1; flappy_W(31, 71) <= 1; flappy_W(31, 72) <= 0; flappy_W(31, 73) <= 0; flappy_W(31, 74) <= 0; flappy_W(31, 75) <= 0; flappy_W(31, 76) <= 0; flappy_W(31, 77) <= 0; flappy_W(31, 78) <= 0; flappy_W(31, 79) <= 0; flappy_W(31, 80) <= 0; flappy_W(31, 81) <= 0; flappy_W(31, 82) <= 0; flappy_W(31, 83) <= 0; flappy_W(31, 84) <= 0; flappy_W(31, 85) <= 0; flappy_W(31, 86) <= 0; flappy_W(31, 87) <= 0; flappy_W(31, 88) <= 0; flappy_W(31, 89) <= 0; flappy_W(31, 90) <= 0; flappy_W(31, 91) <= 0; flappy_W(31, 92) <= 0; flappy_W(31, 93) <= 0; flappy_W(31, 94) <= 0; flappy_W(31, 95) <= 0; flappy_W(31, 96) <= 0; flappy_W(31, 97) <= 0; flappy_W(31, 98) <= 0; flappy_W(31, 99) <= 0; flappy_W(31, 100) <= 0; flappy_W(31, 101) <= 0; flappy_W(31, 102) <= 0; flappy_W(31, 103) <= 0; flappy_W(31, 104) <= 0; flappy_W(31, 105) <= 0; flappy_W(31, 106) <= 0; flappy_W(31, 107) <= 0; flappy_W(31, 108) <= 1; flappy_W(31, 109) <= 1; flappy_W(31, 110) <= 1; flappy_W(31, 111) <= 1; flappy_W(31, 112) <= 1; flappy_W(31, 113) <= 1; flappy_W(31, 114) <= 1; flappy_W(31, 115) <= 1; flappy_W(31, 116) <= 1; flappy_W(31, 117) <= 1; flappy_W(31, 118) <= 1; flappy_W(31, 119) <= 1; flappy_W(31, 120) <= 1; flappy_W(31, 121) <= 1; flappy_W(31, 122) <= 1; flappy_W(31, 123) <= 1; flappy_W(31, 124) <= 1; flappy_W(31, 125) <= 1; flappy_W(31, 126) <= 1; flappy_W(31, 127) <= 1; flappy_W(31, 128) <= 1; flappy_W(31, 129) <= 1; flappy_W(31, 130) <= 1; flappy_W(31, 131) <= 1; flappy_W(31, 132) <= 1; flappy_W(31, 133) <= 1; flappy_W(31, 134) <= 1; flappy_W(31, 135) <= 1; flappy_W(31, 136) <= 1; flappy_W(31, 137) <= 1; flappy_W(31, 138) <= 1; flappy_W(31, 139) <= 1; flappy_W(31, 140) <= 1; flappy_W(31, 141) <= 1; flappy_W(31, 142) <= 1; flappy_W(31, 143) <= 1; flappy_W(31, 144) <= 1; flappy_W(31, 145) <= 1; flappy_W(31, 146) <= 1; flappy_W(31, 147) <= 1; flappy_W(31, 148) <= 1; flappy_W(31, 149) <= 1; flappy_W(31, 150) <= 0; flappy_W(31, 151) <= 0; flappy_W(31, 152) <= 0; flappy_W(31, 153) <= 0; flappy_W(31, 154) <= 0; flappy_W(31, 155) <= 0; flappy_W(31, 156) <= 0; flappy_W(31, 157) <= 0; flappy_W(31, 158) <= 0; flappy_W(31, 159) <= 0; flappy_W(31, 160) <= 0; flappy_W(31, 161) <= 0; flappy_W(31, 162) <= 0; flappy_W(31, 163) <= 0; flappy_W(31, 164) <= 0; flappy_W(31, 165) <= 0; flappy_W(31, 166) <= 0; flappy_W(31, 167) <= 0; flappy_W(31, 168) <= 1; flappy_W(31, 169) <= 1; flappy_W(31, 170) <= 1; flappy_W(31, 171) <= 1; flappy_W(31, 172) <= 1; flappy_W(31, 173) <= 1; flappy_W(31, 174) <= 1; flappy_W(31, 175) <= 1; flappy_W(31, 176) <= 1; flappy_W(31, 177) <= 1; flappy_W(31, 178) <= 1; flappy_W(31, 179) <= 1; flappy_W(31, 180) <= 0; flappy_W(31, 181) <= 0; flappy_W(31, 182) <= 0; flappy_W(31, 183) <= 0; flappy_W(31, 184) <= 0; flappy_W(31, 185) <= 0; flappy_W(31, 186) <= 0; flappy_W(31, 187) <= 0; flappy_W(31, 188) <= 0; flappy_W(31, 189) <= 0; flappy_W(31, 190) <= 0; flappy_W(31, 191) <= 0; flappy_W(31, 192) <= 0; flappy_W(31, 193) <= 0; flappy_W(31, 194) <= 0; flappy_W(31, 195) <= 0; flappy_W(31, 196) <= 0; flappy_W(31, 197) <= 0; flappy_W(31, 198) <= 0; flappy_W(31, 199) <= 0; flappy_W(31, 200) <= 0; flappy_W(31, 201) <= 0; flappy_W(31, 202) <= 0; flappy_W(31, 203) <= 0; flappy_W(31, 204) <= 0; flappy_W(31, 205) <= 0; flappy_W(31, 206) <= 0; flappy_W(31, 207) <= 0; flappy_W(31, 208) <= 0; flappy_W(31, 209) <= 0; flappy_W(31, 210) <= 0; flappy_W(31, 211) <= 0; flappy_W(31, 212) <= 0; flappy_W(31, 213) <= 0; flappy_W(31, 214) <= 0; flappy_W(31, 215) <= 0; flappy_W(31, 216) <= 0; flappy_W(31, 217) <= 0; flappy_W(31, 218) <= 0; flappy_W(31, 219) <= 0; flappy_W(31, 220) <= 0; flappy_W(31, 221) <= 0; flappy_W(31, 222) <= 1; flappy_W(31, 223) <= 1; flappy_W(31, 224) <= 1; flappy_W(31, 225) <= 1; flappy_W(31, 226) <= 1; flappy_W(31, 227) <= 1; flappy_W(31, 228) <= 1; flappy_W(31, 229) <= 1; flappy_W(31, 230) <= 1; flappy_W(31, 231) <= 1; flappy_W(31, 232) <= 1; flappy_W(31, 233) <= 1; flappy_W(31, 234) <= 0; flappy_W(31, 235) <= 0; flappy_W(31, 236) <= 0; flappy_W(31, 237) <= 0; flappy_W(31, 238) <= 0; flappy_W(31, 239) <= 0; flappy_W(31, 240) <= 0; flappy_W(31, 241) <= 0; flappy_W(31, 242) <= 0; flappy_W(31, 243) <= 0; flappy_W(31, 244) <= 0; flappy_W(31, 245) <= 0; flappy_W(31, 246) <= 0; flappy_W(31, 247) <= 0; flappy_W(31, 248) <= 0; flappy_W(31, 249) <= 0; flappy_W(31, 250) <= 0; flappy_W(31, 251) <= 0; flappy_W(31, 252) <= 0; flappy_W(31, 253) <= 0; flappy_W(31, 254) <= 0; flappy_W(31, 255) <= 0; flappy_W(31, 256) <= 0; flappy_W(31, 257) <= 0; flappy_W(31, 258) <= 0; flappy_W(31, 259) <= 0; flappy_W(31, 260) <= 0; flappy_W(31, 261) <= 0; flappy_W(31, 262) <= 0; flappy_W(31, 263) <= 0; flappy_W(31, 264) <= 0; flappy_W(31, 265) <= 0; flappy_W(31, 266) <= 0; flappy_W(31, 267) <= 0; flappy_W(31, 268) <= 0; flappy_W(31, 269) <= 0; flappy_W(31, 270) <= 0; flappy_W(31, 271) <= 0; flappy_W(31, 272) <= 0; flappy_W(31, 273) <= 0; flappy_W(31, 274) <= 0; flappy_W(31, 275) <= 0; flappy_W(31, 276) <= 0; flappy_W(31, 277) <= 0; flappy_W(31, 278) <= 0; flappy_W(31, 279) <= 0; flappy_W(31, 280) <= 0; flappy_W(31, 281) <= 0; flappy_W(31, 282) <= 0; flappy_W(31, 283) <= 0; flappy_W(31, 284) <= 0; flappy_W(31, 285) <= 0; flappy_W(31, 286) <= 0; flappy_W(31, 287) <= 0; flappy_W(31, 288) <= 1; flappy_W(31, 289) <= 1; flappy_W(31, 290) <= 1; flappy_W(31, 291) <= 1; flappy_W(31, 292) <= 1; flappy_W(31, 293) <= 1; flappy_W(31, 294) <= 1; flappy_W(31, 295) <= 1; flappy_W(31, 296) <= 1; flappy_W(31, 297) <= 1; flappy_W(31, 298) <= 1; flappy_W(31, 299) <= 1; flappy_W(31, 300) <= 0; flappy_W(31, 301) <= 0; flappy_W(31, 302) <= 0; flappy_W(31, 303) <= 0; flappy_W(31, 304) <= 0; flappy_W(31, 305) <= 0; flappy_W(31, 306) <= 0; flappy_W(31, 307) <= 0; flappy_W(31, 308) <= 0; flappy_W(31, 309) <= 0; flappy_W(31, 310) <= 0; flappy_W(31, 311) <= 0; flappy_W(31, 312) <= 0; flappy_W(31, 313) <= 0; flappy_W(31, 314) <= 0; flappy_W(31, 315) <= 0; flappy_W(31, 316) <= 0; flappy_W(31, 317) <= 0; flappy_W(31, 318) <= 0; flappy_W(31, 319) <= 0; flappy_W(31, 320) <= 0; flappy_W(31, 321) <= 0; flappy_W(31, 322) <= 0; flappy_W(31, 323) <= 0; flappy_W(31, 324) <= 0; flappy_W(31, 325) <= 0; flappy_W(31, 326) <= 0; flappy_W(31, 327) <= 0; flappy_W(31, 328) <= 0; flappy_W(31, 329) <= 0; flappy_W(31, 330) <= 0; flappy_W(31, 331) <= 0; flappy_W(31, 332) <= 0; flappy_W(31, 333) <= 0; flappy_W(31, 334) <= 0; flappy_W(31, 335) <= 0; flappy_W(31, 336) <= 0; flappy_W(31, 337) <= 0; flappy_W(31, 338) <= 0; flappy_W(31, 339) <= 0; flappy_W(31, 340) <= 0; flappy_W(31, 341) <= 0; flappy_W(31, 342) <= 0; flappy_W(31, 343) <= 0; flappy_W(31, 344) <= 0; flappy_W(31, 345) <= 0; flappy_W(31, 346) <= 0; flappy_W(31, 347) <= 0; flappy_W(31, 348) <= 0; flappy_W(31, 349) <= 0; flappy_W(31, 350) <= 0; flappy_W(31, 351) <= 0; flappy_W(31, 352) <= 0; flappy_W(31, 353) <= 0; flappy_W(31, 354) <= 0; flappy_W(31, 355) <= 0; flappy_W(31, 356) <= 0; flappy_W(31, 357) <= 0; flappy_W(31, 358) <= 0; flappy_W(31, 359) <= 0; flappy_W(31, 360) <= 0; flappy_W(31, 361) <= 0; flappy_W(31, 362) <= 0; flappy_W(31, 363) <= 0; flappy_W(31, 364) <= 0; flappy_W(31, 365) <= 0; flappy_W(31, 366) <= 0; flappy_W(31, 367) <= 0; flappy_W(31, 368) <= 0; flappy_W(31, 369) <= 0; flappy_W(31, 370) <= 0; flappy_W(31, 371) <= 0; flappy_W(31, 372) <= 0; flappy_W(31, 373) <= 0; flappy_W(31, 374) <= 0; flappy_W(31, 375) <= 0; flappy_W(31, 376) <= 0; flappy_W(31, 377) <= 0; flappy_W(31, 378) <= 0; flappy_W(31, 379) <= 0; flappy_W(31, 380) <= 0; flappy_W(31, 381) <= 0; flappy_W(31, 382) <= 0; flappy_W(31, 383) <= 0; flappy_W(31, 384) <= 0; flappy_W(31, 385) <= 0; flappy_W(31, 386) <= 0; flappy_W(31, 387) <= 0; flappy_W(31, 388) <= 0; flappy_W(31, 389) <= 0; flappy_W(31, 390) <= 0; flappy_W(31, 391) <= 0; flappy_W(31, 392) <= 0; flappy_W(31, 393) <= 0; flappy_W(31, 394) <= 0; flappy_W(31, 395) <= 0; flappy_W(31, 396) <= 0; flappy_W(31, 397) <= 0; flappy_W(31, 398) <= 0; flappy_W(31, 399) <= 0; flappy_W(31, 400) <= 0; flappy_W(31, 401) <= 0; flappy_W(31, 402) <= 1; flappy_W(31, 403) <= 1; flappy_W(31, 404) <= 1; flappy_W(31, 405) <= 1; flappy_W(31, 406) <= 1; flappy_W(31, 407) <= 1; flappy_W(31, 408) <= 1; flappy_W(31, 409) <= 1; flappy_W(31, 410) <= 1; flappy_W(31, 411) <= 1; flappy_W(31, 412) <= 1; flappy_W(31, 413) <= 1; flappy_W(31, 414) <= 0; flappy_W(31, 415) <= 0; flappy_W(31, 416) <= 0; flappy_W(31, 417) <= 0; flappy_W(31, 418) <= 0; flappy_W(31, 419) <= 0; flappy_W(31, 420) <= 0; flappy_W(31, 421) <= 0; flappy_W(31, 422) <= 0; flappy_W(31, 423) <= 0; flappy_W(31, 424) <= 0; flappy_W(31, 425) <= 0; flappy_W(31, 426) <= 1; flappy_W(31, 427) <= 1; flappy_W(31, 428) <= 1; flappy_W(31, 429) <= 1; flappy_W(31, 430) <= 1; flappy_W(31, 431) <= 1; flappy_W(31, 432) <= 1; flappy_W(31, 433) <= 1; flappy_W(31, 434) <= 1; flappy_W(31, 435) <= 1; flappy_W(31, 436) <= 1; flappy_W(31, 437) <= 1; flappy_W(31, 438) <= 0; flappy_W(31, 439) <= 0; flappy_W(31, 440) <= 0; flappy_W(31, 441) <= 0; flappy_W(31, 442) <= 0; flappy_W(31, 443) <= 0; flappy_W(31, 444) <= 0; flappy_W(31, 445) <= 0; flappy_W(31, 446) <= 0; flappy_W(31, 447) <= 0; flappy_W(31, 448) <= 0; flappy_W(31, 449) <= 0; flappy_W(31, 450) <= 0; flappy_W(31, 451) <= 0; flappy_W(31, 452) <= 0; flappy_W(31, 453) <= 0; flappy_W(31, 454) <= 0; flappy_W(31, 455) <= 0; flappy_W(31, 456) <= 0; flappy_W(31, 457) <= 0; flappy_W(31, 458) <= 0; flappy_W(31, 459) <= 0; flappy_W(31, 460) <= 0; flappy_W(31, 461) <= 0; flappy_W(31, 462) <= 0; flappy_W(31, 463) <= 0; flappy_W(31, 464) <= 0; flappy_W(31, 465) <= 0; flappy_W(31, 466) <= 0; flappy_W(31, 467) <= 0; flappy_W(31, 468) <= 1; flappy_W(31, 469) <= 1; flappy_W(31, 470) <= 1; flappy_W(31, 471) <= 1; flappy_W(31, 472) <= 1; flappy_W(31, 473) <= 1; flappy_W(31, 474) <= 1; flappy_W(31, 475) <= 1; flappy_W(31, 476) <= 1; flappy_W(31, 477) <= 1; flappy_W(31, 478) <= 1; flappy_W(31, 479) <= 1; flappy_W(31, 480) <= 0; flappy_W(31, 481) <= 0; flappy_W(31, 482) <= 0; flappy_W(31, 483) <= 0; flappy_W(31, 484) <= 0; flappy_W(31, 485) <= 0; flappy_W(31, 486) <= 0; flappy_W(31, 487) <= 0; flappy_W(31, 488) <= 0; flappy_W(31, 489) <= 0; flappy_W(31, 490) <= 0; flappy_W(31, 491) <= 0; flappy_W(31, 492) <= 0; flappy_W(31, 493) <= 0; flappy_W(31, 494) <= 0; flappy_W(31, 495) <= 0; flappy_W(31, 496) <= 0; flappy_W(31, 497) <= 0; flappy_W(31, 498) <= 0; flappy_W(31, 499) <= 0; flappy_W(31, 500) <= 0; flappy_W(31, 501) <= 0; flappy_W(31, 502) <= 0; flappy_W(31, 503) <= 0; flappy_W(31, 504) <= 0; flappy_W(31, 505) <= 0; flappy_W(31, 506) <= 0; flappy_W(31, 507) <= 0; flappy_W(31, 508) <= 0; flappy_W(31, 509) <= 0; flappy_W(31, 510) <= 1; flappy_W(31, 511) <= 1; flappy_W(31, 512) <= 1; flappy_W(31, 513) <= 1; flappy_W(31, 514) <= 1; flappy_W(31, 515) <= 1; flappy_W(31, 516) <= 1; flappy_W(31, 517) <= 1; flappy_W(31, 518) <= 1; flappy_W(31, 519) <= 1; flappy_W(31, 520) <= 1; flappy_W(31, 521) <= 1; flappy_W(31, 522) <= 0; flappy_W(31, 523) <= 0; flappy_W(31, 524) <= 0; flappy_W(31, 525) <= 0; flappy_W(31, 526) <= 0; flappy_W(31, 527) <= 0; flappy_W(31, 528) <= 1; flappy_W(31, 529) <= 1; flappy_W(31, 530) <= 1; flappy_W(31, 531) <= 1; flappy_W(31, 532) <= 1; flappy_W(31, 533) <= 1; flappy_W(31, 534) <= 1; flappy_W(31, 535) <= 1; flappy_W(31, 536) <= 1; flappy_W(31, 537) <= 1; flappy_W(31, 538) <= 1; flappy_W(31, 539) <= 1; flappy_W(31, 540) <= 0; flappy_W(31, 541) <= 0; flappy_W(31, 542) <= 0; flappy_W(31, 543) <= 0; flappy_W(31, 544) <= 0; flappy_W(31, 545) <= 0; flappy_W(31, 546) <= 0; flappy_W(31, 547) <= 0; flappy_W(31, 548) <= 0; flappy_W(31, 549) <= 0; flappy_W(31, 550) <= 0; flappy_W(31, 551) <= 0; flappy_W(31, 552) <= 0; flappy_W(31, 553) <= 0; flappy_W(31, 554) <= 0; flappy_W(31, 555) <= 0; flappy_W(31, 556) <= 0; flappy_W(31, 557) <= 0; flappy_W(31, 558) <= 0; flappy_W(31, 559) <= 0; flappy_W(31, 560) <= 0; flappy_W(31, 561) <= 0; flappy_W(31, 562) <= 0; flappy_W(31, 563) <= 0; flappy_W(31, 564) <= 1; flappy_W(31, 565) <= 1; flappy_W(31, 566) <= 1; flappy_W(31, 567) <= 1; flappy_W(31, 568) <= 1; flappy_W(31, 569) <= 1; flappy_W(31, 570) <= 1; flappy_W(31, 571) <= 1; flappy_W(31, 572) <= 1; flappy_W(31, 573) <= 1; flappy_W(31, 574) <= 1; flappy_W(31, 575) <= 1; flappy_W(31, 576) <= 0; flappy_W(31, 577) <= 0; flappy_W(31, 578) <= 0; flappy_W(31, 579) <= 0; flappy_W(31, 580) <= 0; flappy_W(31, 581) <= 0; flappy_W(31, 582) <= 0; flappy_W(31, 583) <= 0; flappy_W(31, 584) <= 0; flappy_W(31, 585) <= 0; flappy_W(31, 586) <= 0; flappy_W(31, 587) <= 0; flappy_W(31, 588) <= 1; flappy_W(31, 589) <= 1; flappy_W(31, 590) <= 1; flappy_W(31, 591) <= 1; flappy_W(31, 592) <= 1; flappy_W(31, 593) <= 1; 
flappy_W(32, 0) <= 0; flappy_W(32, 1) <= 0; flappy_W(32, 2) <= 0; flappy_W(32, 3) <= 0; flappy_W(32, 4) <= 0; flappy_W(32, 5) <= 0; flappy_W(32, 6) <= 1; flappy_W(32, 7) <= 1; flappy_W(32, 8) <= 1; flappy_W(32, 9) <= 1; flappy_W(32, 10) <= 1; flappy_W(32, 11) <= 1; flappy_W(32, 12) <= 1; flappy_W(32, 13) <= 1; flappy_W(32, 14) <= 1; flappy_W(32, 15) <= 1; flappy_W(32, 16) <= 1; flappy_W(32, 17) <= 1; flappy_W(32, 18) <= 0; flappy_W(32, 19) <= 0; flappy_W(32, 20) <= 0; flappy_W(32, 21) <= 0; flappy_W(32, 22) <= 0; flappy_W(32, 23) <= 0; flappy_W(32, 24) <= 1; flappy_W(32, 25) <= 1; flappy_W(32, 26) <= 1; flappy_W(32, 27) <= 1; flappy_W(32, 28) <= 1; flappy_W(32, 29) <= 1; flappy_W(32, 30) <= 0; flappy_W(32, 31) <= 0; flappy_W(32, 32) <= 0; flappy_W(32, 33) <= 0; flappy_W(32, 34) <= 0; flappy_W(32, 35) <= 0; flappy_W(32, 36) <= 0; flappy_W(32, 37) <= 0; flappy_W(32, 38) <= 0; flappy_W(32, 39) <= 0; flappy_W(32, 40) <= 0; flappy_W(32, 41) <= 0; flappy_W(32, 42) <= 0; flappy_W(32, 43) <= 0; flappy_W(32, 44) <= 0; flappy_W(32, 45) <= 0; flappy_W(32, 46) <= 0; flappy_W(32, 47) <= 0; flappy_W(32, 48) <= 0; flappy_W(32, 49) <= 0; flappy_W(32, 50) <= 0; flappy_W(32, 51) <= 0; flappy_W(32, 52) <= 0; flappy_W(32, 53) <= 0; flappy_W(32, 54) <= 0; flappy_W(32, 55) <= 0; flappy_W(32, 56) <= 0; flappy_W(32, 57) <= 0; flappy_W(32, 58) <= 0; flappy_W(32, 59) <= 0; flappy_W(32, 60) <= 1; flappy_W(32, 61) <= 1; flappy_W(32, 62) <= 1; flappy_W(32, 63) <= 1; flappy_W(32, 64) <= 1; flappy_W(32, 65) <= 1; flappy_W(32, 66) <= 1; flappy_W(32, 67) <= 1; flappy_W(32, 68) <= 1; flappy_W(32, 69) <= 1; flappy_W(32, 70) <= 1; flappy_W(32, 71) <= 1; flappy_W(32, 72) <= 0; flappy_W(32, 73) <= 0; flappy_W(32, 74) <= 0; flappy_W(32, 75) <= 0; flappy_W(32, 76) <= 0; flappy_W(32, 77) <= 0; flappy_W(32, 78) <= 0; flappy_W(32, 79) <= 0; flappy_W(32, 80) <= 0; flappy_W(32, 81) <= 0; flappy_W(32, 82) <= 0; flappy_W(32, 83) <= 0; flappy_W(32, 84) <= 0; flappy_W(32, 85) <= 0; flappy_W(32, 86) <= 0; flappy_W(32, 87) <= 0; flappy_W(32, 88) <= 0; flappy_W(32, 89) <= 0; flappy_W(32, 90) <= 0; flappy_W(32, 91) <= 0; flappy_W(32, 92) <= 0; flappy_W(32, 93) <= 0; flappy_W(32, 94) <= 0; flappy_W(32, 95) <= 0; flappy_W(32, 96) <= 0; flappy_W(32, 97) <= 0; flappy_W(32, 98) <= 0; flappy_W(32, 99) <= 0; flappy_W(32, 100) <= 0; flappy_W(32, 101) <= 0; flappy_W(32, 102) <= 0; flappy_W(32, 103) <= 0; flappy_W(32, 104) <= 0; flappy_W(32, 105) <= 0; flappy_W(32, 106) <= 0; flappy_W(32, 107) <= 0; flappy_W(32, 108) <= 1; flappy_W(32, 109) <= 1; flappy_W(32, 110) <= 1; flappy_W(32, 111) <= 1; flappy_W(32, 112) <= 1; flappy_W(32, 113) <= 1; flappy_W(32, 114) <= 1; flappy_W(32, 115) <= 1; flappy_W(32, 116) <= 1; flappy_W(32, 117) <= 1; flappy_W(32, 118) <= 1; flappy_W(32, 119) <= 1; flappy_W(32, 120) <= 1; flappy_W(32, 121) <= 1; flappy_W(32, 122) <= 1; flappy_W(32, 123) <= 1; flappy_W(32, 124) <= 1; flappy_W(32, 125) <= 1; flappy_W(32, 126) <= 1; flappy_W(32, 127) <= 1; flappy_W(32, 128) <= 1; flappy_W(32, 129) <= 1; flappy_W(32, 130) <= 1; flappy_W(32, 131) <= 1; flappy_W(32, 132) <= 1; flappy_W(32, 133) <= 1; flappy_W(32, 134) <= 1; flappy_W(32, 135) <= 1; flappy_W(32, 136) <= 1; flappy_W(32, 137) <= 1; flappy_W(32, 138) <= 1; flappy_W(32, 139) <= 1; flappy_W(32, 140) <= 1; flappy_W(32, 141) <= 1; flappy_W(32, 142) <= 1; flappy_W(32, 143) <= 1; flappy_W(32, 144) <= 1; flappy_W(32, 145) <= 1; flappy_W(32, 146) <= 1; flappy_W(32, 147) <= 1; flappy_W(32, 148) <= 1; flappy_W(32, 149) <= 1; flappy_W(32, 150) <= 0; flappy_W(32, 151) <= 0; flappy_W(32, 152) <= 0; flappy_W(32, 153) <= 0; flappy_W(32, 154) <= 0; flappy_W(32, 155) <= 0; flappy_W(32, 156) <= 0; flappy_W(32, 157) <= 0; flappy_W(32, 158) <= 0; flappy_W(32, 159) <= 0; flappy_W(32, 160) <= 0; flappy_W(32, 161) <= 0; flappy_W(32, 162) <= 0; flappy_W(32, 163) <= 0; flappy_W(32, 164) <= 0; flappy_W(32, 165) <= 0; flappy_W(32, 166) <= 0; flappy_W(32, 167) <= 0; flappy_W(32, 168) <= 1; flappy_W(32, 169) <= 1; flappy_W(32, 170) <= 1; flappy_W(32, 171) <= 1; flappy_W(32, 172) <= 1; flappy_W(32, 173) <= 1; flappy_W(32, 174) <= 1; flappy_W(32, 175) <= 1; flappy_W(32, 176) <= 1; flappy_W(32, 177) <= 1; flappy_W(32, 178) <= 1; flappy_W(32, 179) <= 1; flappy_W(32, 180) <= 0; flappy_W(32, 181) <= 0; flappy_W(32, 182) <= 0; flappy_W(32, 183) <= 0; flappy_W(32, 184) <= 0; flappy_W(32, 185) <= 0; flappy_W(32, 186) <= 0; flappy_W(32, 187) <= 0; flappy_W(32, 188) <= 0; flappy_W(32, 189) <= 0; flappy_W(32, 190) <= 0; flappy_W(32, 191) <= 0; flappy_W(32, 192) <= 0; flappy_W(32, 193) <= 0; flappy_W(32, 194) <= 0; flappy_W(32, 195) <= 0; flappy_W(32, 196) <= 0; flappy_W(32, 197) <= 0; flappy_W(32, 198) <= 0; flappy_W(32, 199) <= 0; flappy_W(32, 200) <= 0; flappy_W(32, 201) <= 0; flappy_W(32, 202) <= 0; flappy_W(32, 203) <= 0; flappy_W(32, 204) <= 0; flappy_W(32, 205) <= 0; flappy_W(32, 206) <= 0; flappy_W(32, 207) <= 0; flappy_W(32, 208) <= 0; flappy_W(32, 209) <= 0; flappy_W(32, 210) <= 0; flappy_W(32, 211) <= 0; flappy_W(32, 212) <= 0; flappy_W(32, 213) <= 0; flappy_W(32, 214) <= 0; flappy_W(32, 215) <= 0; flappy_W(32, 216) <= 0; flappy_W(32, 217) <= 0; flappy_W(32, 218) <= 0; flappy_W(32, 219) <= 0; flappy_W(32, 220) <= 0; flappy_W(32, 221) <= 0; flappy_W(32, 222) <= 1; flappy_W(32, 223) <= 1; flappy_W(32, 224) <= 1; flappy_W(32, 225) <= 1; flappy_W(32, 226) <= 1; flappy_W(32, 227) <= 1; flappy_W(32, 228) <= 1; flappy_W(32, 229) <= 1; flappy_W(32, 230) <= 1; flappy_W(32, 231) <= 1; flappy_W(32, 232) <= 1; flappy_W(32, 233) <= 1; flappy_W(32, 234) <= 0; flappy_W(32, 235) <= 0; flappy_W(32, 236) <= 0; flappy_W(32, 237) <= 0; flappy_W(32, 238) <= 0; flappy_W(32, 239) <= 0; flappy_W(32, 240) <= 0; flappy_W(32, 241) <= 0; flappy_W(32, 242) <= 0; flappy_W(32, 243) <= 0; flappy_W(32, 244) <= 0; flappy_W(32, 245) <= 0; flappy_W(32, 246) <= 0; flappy_W(32, 247) <= 0; flappy_W(32, 248) <= 0; flappy_W(32, 249) <= 0; flappy_W(32, 250) <= 0; flappy_W(32, 251) <= 0; flappy_W(32, 252) <= 0; flappy_W(32, 253) <= 0; flappy_W(32, 254) <= 0; flappy_W(32, 255) <= 0; flappy_W(32, 256) <= 0; flappy_W(32, 257) <= 0; flappy_W(32, 258) <= 0; flappy_W(32, 259) <= 0; flappy_W(32, 260) <= 0; flappy_W(32, 261) <= 0; flappy_W(32, 262) <= 0; flappy_W(32, 263) <= 0; flappy_W(32, 264) <= 0; flappy_W(32, 265) <= 0; flappy_W(32, 266) <= 0; flappy_W(32, 267) <= 0; flappy_W(32, 268) <= 0; flappy_W(32, 269) <= 0; flappy_W(32, 270) <= 0; flappy_W(32, 271) <= 0; flappy_W(32, 272) <= 0; flappy_W(32, 273) <= 0; flappy_W(32, 274) <= 0; flappy_W(32, 275) <= 0; flappy_W(32, 276) <= 0; flappy_W(32, 277) <= 0; flappy_W(32, 278) <= 0; flappy_W(32, 279) <= 0; flappy_W(32, 280) <= 0; flappy_W(32, 281) <= 0; flappy_W(32, 282) <= 0; flappy_W(32, 283) <= 0; flappy_W(32, 284) <= 0; flappy_W(32, 285) <= 0; flappy_W(32, 286) <= 0; flappy_W(32, 287) <= 0; flappy_W(32, 288) <= 1; flappy_W(32, 289) <= 1; flappy_W(32, 290) <= 1; flappy_W(32, 291) <= 1; flappy_W(32, 292) <= 1; flappy_W(32, 293) <= 1; flappy_W(32, 294) <= 1; flappy_W(32, 295) <= 1; flappy_W(32, 296) <= 1; flappy_W(32, 297) <= 1; flappy_W(32, 298) <= 1; flappy_W(32, 299) <= 1; flappy_W(32, 300) <= 0; flappy_W(32, 301) <= 0; flappy_W(32, 302) <= 0; flappy_W(32, 303) <= 0; flappy_W(32, 304) <= 0; flappy_W(32, 305) <= 0; flappy_W(32, 306) <= 0; flappy_W(32, 307) <= 0; flappy_W(32, 308) <= 0; flappy_W(32, 309) <= 0; flappy_W(32, 310) <= 0; flappy_W(32, 311) <= 0; flappy_W(32, 312) <= 0; flappy_W(32, 313) <= 0; flappy_W(32, 314) <= 0; flappy_W(32, 315) <= 0; flappy_W(32, 316) <= 0; flappy_W(32, 317) <= 0; flappy_W(32, 318) <= 0; flappy_W(32, 319) <= 0; flappy_W(32, 320) <= 0; flappy_W(32, 321) <= 0; flappy_W(32, 322) <= 0; flappy_W(32, 323) <= 0; flappy_W(32, 324) <= 0; flappy_W(32, 325) <= 0; flappy_W(32, 326) <= 0; flappy_W(32, 327) <= 0; flappy_W(32, 328) <= 0; flappy_W(32, 329) <= 0; flappy_W(32, 330) <= 0; flappy_W(32, 331) <= 0; flappy_W(32, 332) <= 0; flappy_W(32, 333) <= 0; flappy_W(32, 334) <= 0; flappy_W(32, 335) <= 0; flappy_W(32, 336) <= 0; flappy_W(32, 337) <= 0; flappy_W(32, 338) <= 0; flappy_W(32, 339) <= 0; flappy_W(32, 340) <= 0; flappy_W(32, 341) <= 0; flappy_W(32, 342) <= 0; flappy_W(32, 343) <= 0; flappy_W(32, 344) <= 0; flappy_W(32, 345) <= 0; flappy_W(32, 346) <= 0; flappy_W(32, 347) <= 0; flappy_W(32, 348) <= 0; flappy_W(32, 349) <= 0; flappy_W(32, 350) <= 0; flappy_W(32, 351) <= 0; flappy_W(32, 352) <= 0; flappy_W(32, 353) <= 0; flappy_W(32, 354) <= 0; flappy_W(32, 355) <= 0; flappy_W(32, 356) <= 0; flappy_W(32, 357) <= 0; flappy_W(32, 358) <= 0; flappy_W(32, 359) <= 0; flappy_W(32, 360) <= 0; flappy_W(32, 361) <= 0; flappy_W(32, 362) <= 0; flappy_W(32, 363) <= 0; flappy_W(32, 364) <= 0; flappy_W(32, 365) <= 0; flappy_W(32, 366) <= 0; flappy_W(32, 367) <= 0; flappy_W(32, 368) <= 0; flappy_W(32, 369) <= 0; flappy_W(32, 370) <= 0; flappy_W(32, 371) <= 0; flappy_W(32, 372) <= 0; flappy_W(32, 373) <= 0; flappy_W(32, 374) <= 0; flappy_W(32, 375) <= 0; flappy_W(32, 376) <= 0; flappy_W(32, 377) <= 0; flappy_W(32, 378) <= 0; flappy_W(32, 379) <= 0; flappy_W(32, 380) <= 0; flappy_W(32, 381) <= 0; flappy_W(32, 382) <= 0; flappy_W(32, 383) <= 0; flappy_W(32, 384) <= 0; flappy_W(32, 385) <= 0; flappy_W(32, 386) <= 0; flappy_W(32, 387) <= 0; flappy_W(32, 388) <= 0; flappy_W(32, 389) <= 0; flappy_W(32, 390) <= 0; flappy_W(32, 391) <= 0; flappy_W(32, 392) <= 0; flappy_W(32, 393) <= 0; flappy_W(32, 394) <= 0; flappy_W(32, 395) <= 0; flappy_W(32, 396) <= 0; flappy_W(32, 397) <= 0; flappy_W(32, 398) <= 0; flappy_W(32, 399) <= 0; flappy_W(32, 400) <= 0; flappy_W(32, 401) <= 0; flappy_W(32, 402) <= 1; flappy_W(32, 403) <= 1; flappy_W(32, 404) <= 1; flappy_W(32, 405) <= 1; flappy_W(32, 406) <= 1; flappy_W(32, 407) <= 1; flappy_W(32, 408) <= 1; flappy_W(32, 409) <= 1; flappy_W(32, 410) <= 1; flappy_W(32, 411) <= 1; flappy_W(32, 412) <= 1; flappy_W(32, 413) <= 1; flappy_W(32, 414) <= 0; flappy_W(32, 415) <= 0; flappy_W(32, 416) <= 0; flappy_W(32, 417) <= 0; flappy_W(32, 418) <= 0; flappy_W(32, 419) <= 0; flappy_W(32, 420) <= 0; flappy_W(32, 421) <= 0; flappy_W(32, 422) <= 0; flappy_W(32, 423) <= 0; flappy_W(32, 424) <= 0; flappy_W(32, 425) <= 0; flappy_W(32, 426) <= 1; flappy_W(32, 427) <= 1; flappy_W(32, 428) <= 1; flappy_W(32, 429) <= 1; flappy_W(32, 430) <= 1; flappy_W(32, 431) <= 1; flappy_W(32, 432) <= 1; flappy_W(32, 433) <= 1; flappy_W(32, 434) <= 1; flappy_W(32, 435) <= 1; flappy_W(32, 436) <= 1; flappy_W(32, 437) <= 1; flappy_W(32, 438) <= 0; flappy_W(32, 439) <= 0; flappy_W(32, 440) <= 0; flappy_W(32, 441) <= 0; flappy_W(32, 442) <= 0; flappy_W(32, 443) <= 0; flappy_W(32, 444) <= 0; flappy_W(32, 445) <= 0; flappy_W(32, 446) <= 0; flappy_W(32, 447) <= 0; flappy_W(32, 448) <= 0; flappy_W(32, 449) <= 0; flappy_W(32, 450) <= 0; flappy_W(32, 451) <= 0; flappy_W(32, 452) <= 0; flappy_W(32, 453) <= 0; flappy_W(32, 454) <= 0; flappy_W(32, 455) <= 0; flappy_W(32, 456) <= 0; flappy_W(32, 457) <= 0; flappy_W(32, 458) <= 0; flappy_W(32, 459) <= 0; flappy_W(32, 460) <= 0; flappy_W(32, 461) <= 0; flappy_W(32, 462) <= 0; flappy_W(32, 463) <= 0; flappy_W(32, 464) <= 0; flappy_W(32, 465) <= 0; flappy_W(32, 466) <= 0; flappy_W(32, 467) <= 0; flappy_W(32, 468) <= 1; flappy_W(32, 469) <= 1; flappy_W(32, 470) <= 1; flappy_W(32, 471) <= 1; flappy_W(32, 472) <= 1; flappy_W(32, 473) <= 1; flappy_W(32, 474) <= 1; flappy_W(32, 475) <= 1; flappy_W(32, 476) <= 1; flappy_W(32, 477) <= 1; flappy_W(32, 478) <= 1; flappy_W(32, 479) <= 1; flappy_W(32, 480) <= 0; flappy_W(32, 481) <= 0; flappy_W(32, 482) <= 0; flappy_W(32, 483) <= 0; flappy_W(32, 484) <= 0; flappy_W(32, 485) <= 0; flappy_W(32, 486) <= 0; flappy_W(32, 487) <= 0; flappy_W(32, 488) <= 0; flappy_W(32, 489) <= 0; flappy_W(32, 490) <= 0; flappy_W(32, 491) <= 0; flappy_W(32, 492) <= 0; flappy_W(32, 493) <= 0; flappy_W(32, 494) <= 0; flappy_W(32, 495) <= 0; flappy_W(32, 496) <= 0; flappy_W(32, 497) <= 0; flappy_W(32, 498) <= 0; flappy_W(32, 499) <= 0; flappy_W(32, 500) <= 0; flappy_W(32, 501) <= 0; flappy_W(32, 502) <= 0; flappy_W(32, 503) <= 0; flappy_W(32, 504) <= 0; flappy_W(32, 505) <= 0; flappy_W(32, 506) <= 0; flappy_W(32, 507) <= 0; flappy_W(32, 508) <= 0; flappy_W(32, 509) <= 0; flappy_W(32, 510) <= 1; flappy_W(32, 511) <= 1; flappy_W(32, 512) <= 1; flappy_W(32, 513) <= 1; flappy_W(32, 514) <= 1; flappy_W(32, 515) <= 1; flappy_W(32, 516) <= 1; flappy_W(32, 517) <= 1; flappy_W(32, 518) <= 1; flappy_W(32, 519) <= 1; flappy_W(32, 520) <= 1; flappy_W(32, 521) <= 1; flappy_W(32, 522) <= 0; flappy_W(32, 523) <= 0; flappy_W(32, 524) <= 0; flappy_W(32, 525) <= 0; flappy_W(32, 526) <= 0; flappy_W(32, 527) <= 0; flappy_W(32, 528) <= 1; flappy_W(32, 529) <= 1; flappy_W(32, 530) <= 1; flappy_W(32, 531) <= 1; flappy_W(32, 532) <= 1; flappy_W(32, 533) <= 1; flappy_W(32, 534) <= 1; flappy_W(32, 535) <= 1; flappy_W(32, 536) <= 1; flappy_W(32, 537) <= 1; flappy_W(32, 538) <= 1; flappy_W(32, 539) <= 1; flappy_W(32, 540) <= 0; flappy_W(32, 541) <= 0; flappy_W(32, 542) <= 0; flappy_W(32, 543) <= 0; flappy_W(32, 544) <= 0; flappy_W(32, 545) <= 0; flappy_W(32, 546) <= 0; flappy_W(32, 547) <= 0; flappy_W(32, 548) <= 0; flappy_W(32, 549) <= 0; flappy_W(32, 550) <= 0; flappy_W(32, 551) <= 0; flappy_W(32, 552) <= 0; flappy_W(32, 553) <= 0; flappy_W(32, 554) <= 0; flappy_W(32, 555) <= 0; flappy_W(32, 556) <= 0; flappy_W(32, 557) <= 0; flappy_W(32, 558) <= 0; flappy_W(32, 559) <= 0; flappy_W(32, 560) <= 0; flappy_W(32, 561) <= 0; flappy_W(32, 562) <= 0; flappy_W(32, 563) <= 0; flappy_W(32, 564) <= 1; flappy_W(32, 565) <= 1; flappy_W(32, 566) <= 1; flappy_W(32, 567) <= 1; flappy_W(32, 568) <= 1; flappy_W(32, 569) <= 1; flappy_W(32, 570) <= 1; flappy_W(32, 571) <= 1; flappy_W(32, 572) <= 1; flappy_W(32, 573) <= 1; flappy_W(32, 574) <= 1; flappy_W(32, 575) <= 1; flappy_W(32, 576) <= 0; flappy_W(32, 577) <= 0; flappy_W(32, 578) <= 0; flappy_W(32, 579) <= 0; flappy_W(32, 580) <= 0; flappy_W(32, 581) <= 0; flappy_W(32, 582) <= 0; flappy_W(32, 583) <= 0; flappy_W(32, 584) <= 0; flappy_W(32, 585) <= 0; flappy_W(32, 586) <= 0; flappy_W(32, 587) <= 0; flappy_W(32, 588) <= 1; flappy_W(32, 589) <= 1; flappy_W(32, 590) <= 1; flappy_W(32, 591) <= 1; flappy_W(32, 592) <= 1; flappy_W(32, 593) <= 1; 
flappy_W(33, 0) <= 0; flappy_W(33, 1) <= 0; flappy_W(33, 2) <= 0; flappy_W(33, 3) <= 0; flappy_W(33, 4) <= 0; flappy_W(33, 5) <= 0; flappy_W(33, 6) <= 1; flappy_W(33, 7) <= 1; flappy_W(33, 8) <= 1; flappy_W(33, 9) <= 1; flappy_W(33, 10) <= 1; flappy_W(33, 11) <= 1; flappy_W(33, 12) <= 1; flappy_W(33, 13) <= 1; flappy_W(33, 14) <= 1; flappy_W(33, 15) <= 1; flappy_W(33, 16) <= 1; flappy_W(33, 17) <= 1; flappy_W(33, 18) <= 0; flappy_W(33, 19) <= 0; flappy_W(33, 20) <= 0; flappy_W(33, 21) <= 0; flappy_W(33, 22) <= 0; flappy_W(33, 23) <= 0; flappy_W(33, 24) <= 1; flappy_W(33, 25) <= 1; flappy_W(33, 26) <= 1; flappy_W(33, 27) <= 1; flappy_W(33, 28) <= 1; flappy_W(33, 29) <= 1; flappy_W(33, 30) <= 0; flappy_W(33, 31) <= 0; flappy_W(33, 32) <= 0; flappy_W(33, 33) <= 0; flappy_W(33, 34) <= 0; flappy_W(33, 35) <= 0; flappy_W(33, 36) <= 0; flappy_W(33, 37) <= 0; flappy_W(33, 38) <= 0; flappy_W(33, 39) <= 0; flappy_W(33, 40) <= 0; flappy_W(33, 41) <= 0; flappy_W(33, 42) <= 0; flappy_W(33, 43) <= 0; flappy_W(33, 44) <= 0; flappy_W(33, 45) <= 0; flappy_W(33, 46) <= 0; flappy_W(33, 47) <= 0; flappy_W(33, 48) <= 0; flappy_W(33, 49) <= 0; flappy_W(33, 50) <= 0; flappy_W(33, 51) <= 0; flappy_W(33, 52) <= 0; flappy_W(33, 53) <= 0; flappy_W(33, 54) <= 0; flappy_W(33, 55) <= 0; flappy_W(33, 56) <= 0; flappy_W(33, 57) <= 0; flappy_W(33, 58) <= 0; flappy_W(33, 59) <= 0; flappy_W(33, 60) <= 1; flappy_W(33, 61) <= 1; flappy_W(33, 62) <= 1; flappy_W(33, 63) <= 1; flappy_W(33, 64) <= 1; flappy_W(33, 65) <= 1; flappy_W(33, 66) <= 1; flappy_W(33, 67) <= 1; flappy_W(33, 68) <= 1; flappy_W(33, 69) <= 1; flappy_W(33, 70) <= 1; flappy_W(33, 71) <= 1; flappy_W(33, 72) <= 0; flappy_W(33, 73) <= 0; flappy_W(33, 74) <= 0; flappy_W(33, 75) <= 0; flappy_W(33, 76) <= 0; flappy_W(33, 77) <= 0; flappy_W(33, 78) <= 0; flappy_W(33, 79) <= 0; flappy_W(33, 80) <= 0; flappy_W(33, 81) <= 0; flappy_W(33, 82) <= 0; flappy_W(33, 83) <= 0; flappy_W(33, 84) <= 0; flappy_W(33, 85) <= 0; flappy_W(33, 86) <= 0; flappy_W(33, 87) <= 0; flappy_W(33, 88) <= 0; flappy_W(33, 89) <= 0; flappy_W(33, 90) <= 0; flappy_W(33, 91) <= 0; flappy_W(33, 92) <= 0; flappy_W(33, 93) <= 0; flappy_W(33, 94) <= 0; flappy_W(33, 95) <= 0; flappy_W(33, 96) <= 0; flappy_W(33, 97) <= 0; flappy_W(33, 98) <= 0; flappy_W(33, 99) <= 0; flappy_W(33, 100) <= 0; flappy_W(33, 101) <= 0; flappy_W(33, 102) <= 0; flappy_W(33, 103) <= 0; flappy_W(33, 104) <= 0; flappy_W(33, 105) <= 0; flappy_W(33, 106) <= 0; flappy_W(33, 107) <= 0; flappy_W(33, 108) <= 1; flappy_W(33, 109) <= 1; flappy_W(33, 110) <= 1; flappy_W(33, 111) <= 1; flappy_W(33, 112) <= 1; flappy_W(33, 113) <= 1; flappy_W(33, 114) <= 1; flappy_W(33, 115) <= 1; flappy_W(33, 116) <= 1; flappy_W(33, 117) <= 1; flappy_W(33, 118) <= 1; flappy_W(33, 119) <= 1; flappy_W(33, 120) <= 1; flappy_W(33, 121) <= 1; flappy_W(33, 122) <= 1; flappy_W(33, 123) <= 1; flappy_W(33, 124) <= 1; flappy_W(33, 125) <= 1; flappy_W(33, 126) <= 1; flappy_W(33, 127) <= 1; flappy_W(33, 128) <= 1; flappy_W(33, 129) <= 1; flappy_W(33, 130) <= 1; flappy_W(33, 131) <= 1; flappy_W(33, 132) <= 1; flappy_W(33, 133) <= 1; flappy_W(33, 134) <= 1; flappy_W(33, 135) <= 1; flappy_W(33, 136) <= 1; flappy_W(33, 137) <= 1; flappy_W(33, 138) <= 1; flappy_W(33, 139) <= 1; flappy_W(33, 140) <= 1; flappy_W(33, 141) <= 1; flappy_W(33, 142) <= 1; flappy_W(33, 143) <= 1; flappy_W(33, 144) <= 1; flappy_W(33, 145) <= 1; flappy_W(33, 146) <= 1; flappy_W(33, 147) <= 1; flappy_W(33, 148) <= 1; flappy_W(33, 149) <= 1; flappy_W(33, 150) <= 0; flappy_W(33, 151) <= 0; flappy_W(33, 152) <= 0; flappy_W(33, 153) <= 0; flappy_W(33, 154) <= 0; flappy_W(33, 155) <= 0; flappy_W(33, 156) <= 0; flappy_W(33, 157) <= 0; flappy_W(33, 158) <= 0; flappy_W(33, 159) <= 0; flappy_W(33, 160) <= 0; flappy_W(33, 161) <= 0; flappy_W(33, 162) <= 0; flappy_W(33, 163) <= 0; flappy_W(33, 164) <= 0; flappy_W(33, 165) <= 0; flappy_W(33, 166) <= 0; flappy_W(33, 167) <= 0; flappy_W(33, 168) <= 1; flappy_W(33, 169) <= 1; flappy_W(33, 170) <= 1; flappy_W(33, 171) <= 1; flappy_W(33, 172) <= 1; flappy_W(33, 173) <= 1; flappy_W(33, 174) <= 1; flappy_W(33, 175) <= 1; flappy_W(33, 176) <= 1; flappy_W(33, 177) <= 1; flappy_W(33, 178) <= 1; flappy_W(33, 179) <= 1; flappy_W(33, 180) <= 0; flappy_W(33, 181) <= 0; flappy_W(33, 182) <= 0; flappy_W(33, 183) <= 0; flappy_W(33, 184) <= 0; flappy_W(33, 185) <= 0; flappy_W(33, 186) <= 0; flappy_W(33, 187) <= 0; flappy_W(33, 188) <= 0; flappy_W(33, 189) <= 0; flappy_W(33, 190) <= 0; flappy_W(33, 191) <= 0; flappy_W(33, 192) <= 0; flappy_W(33, 193) <= 0; flappy_W(33, 194) <= 0; flappy_W(33, 195) <= 0; flappy_W(33, 196) <= 0; flappy_W(33, 197) <= 0; flappy_W(33, 198) <= 0; flappy_W(33, 199) <= 0; flappy_W(33, 200) <= 0; flappy_W(33, 201) <= 0; flappy_W(33, 202) <= 0; flappy_W(33, 203) <= 0; flappy_W(33, 204) <= 0; flappy_W(33, 205) <= 0; flappy_W(33, 206) <= 0; flappy_W(33, 207) <= 0; flappy_W(33, 208) <= 0; flappy_W(33, 209) <= 0; flappy_W(33, 210) <= 0; flappy_W(33, 211) <= 0; flappy_W(33, 212) <= 0; flappy_W(33, 213) <= 0; flappy_W(33, 214) <= 0; flappy_W(33, 215) <= 0; flappy_W(33, 216) <= 0; flappy_W(33, 217) <= 0; flappy_W(33, 218) <= 0; flappy_W(33, 219) <= 0; flappy_W(33, 220) <= 0; flappy_W(33, 221) <= 0; flappy_W(33, 222) <= 1; flappy_W(33, 223) <= 1; flappy_W(33, 224) <= 1; flappy_W(33, 225) <= 1; flappy_W(33, 226) <= 1; flappy_W(33, 227) <= 1; flappy_W(33, 228) <= 1; flappy_W(33, 229) <= 1; flappy_W(33, 230) <= 1; flappy_W(33, 231) <= 1; flappy_W(33, 232) <= 1; flappy_W(33, 233) <= 1; flappy_W(33, 234) <= 0; flappy_W(33, 235) <= 0; flappy_W(33, 236) <= 0; flappy_W(33, 237) <= 0; flappy_W(33, 238) <= 0; flappy_W(33, 239) <= 0; flappy_W(33, 240) <= 0; flappy_W(33, 241) <= 0; flappy_W(33, 242) <= 0; flappy_W(33, 243) <= 0; flappy_W(33, 244) <= 0; flappy_W(33, 245) <= 0; flappy_W(33, 246) <= 0; flappy_W(33, 247) <= 0; flappy_W(33, 248) <= 0; flappy_W(33, 249) <= 0; flappy_W(33, 250) <= 0; flappy_W(33, 251) <= 0; flappy_W(33, 252) <= 0; flappy_W(33, 253) <= 0; flappy_W(33, 254) <= 0; flappy_W(33, 255) <= 0; flappy_W(33, 256) <= 0; flappy_W(33, 257) <= 0; flappy_W(33, 258) <= 0; flappy_W(33, 259) <= 0; flappy_W(33, 260) <= 0; flappy_W(33, 261) <= 0; flappy_W(33, 262) <= 0; flappy_W(33, 263) <= 0; flappy_W(33, 264) <= 0; flappy_W(33, 265) <= 0; flappy_W(33, 266) <= 0; flappy_W(33, 267) <= 0; flappy_W(33, 268) <= 0; flappy_W(33, 269) <= 0; flappy_W(33, 270) <= 0; flappy_W(33, 271) <= 0; flappy_W(33, 272) <= 0; flappy_W(33, 273) <= 0; flappy_W(33, 274) <= 0; flappy_W(33, 275) <= 0; flappy_W(33, 276) <= 0; flappy_W(33, 277) <= 0; flappy_W(33, 278) <= 0; flappy_W(33, 279) <= 0; flappy_W(33, 280) <= 0; flappy_W(33, 281) <= 0; flappy_W(33, 282) <= 0; flappy_W(33, 283) <= 0; flappy_W(33, 284) <= 0; flappy_W(33, 285) <= 0; flappy_W(33, 286) <= 0; flappy_W(33, 287) <= 0; flappy_W(33, 288) <= 1; flappy_W(33, 289) <= 1; flappy_W(33, 290) <= 1; flappy_W(33, 291) <= 1; flappy_W(33, 292) <= 1; flappy_W(33, 293) <= 1; flappy_W(33, 294) <= 1; flappy_W(33, 295) <= 1; flappy_W(33, 296) <= 1; flappy_W(33, 297) <= 1; flappy_W(33, 298) <= 1; flappy_W(33, 299) <= 1; flappy_W(33, 300) <= 0; flappy_W(33, 301) <= 0; flappy_W(33, 302) <= 0; flappy_W(33, 303) <= 0; flappy_W(33, 304) <= 0; flappy_W(33, 305) <= 0; flappy_W(33, 306) <= 0; flappy_W(33, 307) <= 0; flappy_W(33, 308) <= 0; flappy_W(33, 309) <= 0; flappy_W(33, 310) <= 0; flappy_W(33, 311) <= 0; flappy_W(33, 312) <= 0; flappy_W(33, 313) <= 0; flappy_W(33, 314) <= 0; flappy_W(33, 315) <= 0; flappy_W(33, 316) <= 0; flappy_W(33, 317) <= 0; flappy_W(33, 318) <= 0; flappy_W(33, 319) <= 0; flappy_W(33, 320) <= 0; flappy_W(33, 321) <= 0; flappy_W(33, 322) <= 0; flappy_W(33, 323) <= 0; flappy_W(33, 324) <= 0; flappy_W(33, 325) <= 0; flappy_W(33, 326) <= 0; flappy_W(33, 327) <= 0; flappy_W(33, 328) <= 0; flappy_W(33, 329) <= 0; flappy_W(33, 330) <= 0; flappy_W(33, 331) <= 0; flappy_W(33, 332) <= 0; flappy_W(33, 333) <= 0; flappy_W(33, 334) <= 0; flappy_W(33, 335) <= 0; flappy_W(33, 336) <= 0; flappy_W(33, 337) <= 0; flappy_W(33, 338) <= 0; flappy_W(33, 339) <= 0; flappy_W(33, 340) <= 0; flappy_W(33, 341) <= 0; flappy_W(33, 342) <= 0; flappy_W(33, 343) <= 0; flappy_W(33, 344) <= 0; flappy_W(33, 345) <= 0; flappy_W(33, 346) <= 0; flappy_W(33, 347) <= 0; flappy_W(33, 348) <= 0; flappy_W(33, 349) <= 0; flappy_W(33, 350) <= 0; flappy_W(33, 351) <= 0; flappy_W(33, 352) <= 0; flappy_W(33, 353) <= 0; flappy_W(33, 354) <= 0; flappy_W(33, 355) <= 0; flappy_W(33, 356) <= 0; flappy_W(33, 357) <= 0; flappy_W(33, 358) <= 0; flappy_W(33, 359) <= 0; flappy_W(33, 360) <= 0; flappy_W(33, 361) <= 0; flappy_W(33, 362) <= 0; flappy_W(33, 363) <= 0; flappy_W(33, 364) <= 0; flappy_W(33, 365) <= 0; flappy_W(33, 366) <= 0; flappy_W(33, 367) <= 0; flappy_W(33, 368) <= 0; flappy_W(33, 369) <= 0; flappy_W(33, 370) <= 0; flappy_W(33, 371) <= 0; flappy_W(33, 372) <= 0; flappy_W(33, 373) <= 0; flappy_W(33, 374) <= 0; flappy_W(33, 375) <= 0; flappy_W(33, 376) <= 0; flappy_W(33, 377) <= 0; flappy_W(33, 378) <= 0; flappy_W(33, 379) <= 0; flappy_W(33, 380) <= 0; flappy_W(33, 381) <= 0; flappy_W(33, 382) <= 0; flappy_W(33, 383) <= 0; flappy_W(33, 384) <= 0; flappy_W(33, 385) <= 0; flappy_W(33, 386) <= 0; flappy_W(33, 387) <= 0; flappy_W(33, 388) <= 0; flappy_W(33, 389) <= 0; flappy_W(33, 390) <= 0; flappy_W(33, 391) <= 0; flappy_W(33, 392) <= 0; flappy_W(33, 393) <= 0; flappy_W(33, 394) <= 0; flappy_W(33, 395) <= 0; flappy_W(33, 396) <= 0; flappy_W(33, 397) <= 0; flappy_W(33, 398) <= 0; flappy_W(33, 399) <= 0; flappy_W(33, 400) <= 0; flappy_W(33, 401) <= 0; flappy_W(33, 402) <= 1; flappy_W(33, 403) <= 1; flappy_W(33, 404) <= 1; flappy_W(33, 405) <= 1; flappy_W(33, 406) <= 1; flappy_W(33, 407) <= 1; flappy_W(33, 408) <= 1; flappy_W(33, 409) <= 1; flappy_W(33, 410) <= 1; flappy_W(33, 411) <= 1; flappy_W(33, 412) <= 1; flappy_W(33, 413) <= 1; flappy_W(33, 414) <= 0; flappy_W(33, 415) <= 0; flappy_W(33, 416) <= 0; flappy_W(33, 417) <= 0; flappy_W(33, 418) <= 0; flappy_W(33, 419) <= 0; flappy_W(33, 420) <= 0; flappy_W(33, 421) <= 0; flappy_W(33, 422) <= 0; flappy_W(33, 423) <= 0; flappy_W(33, 424) <= 0; flappy_W(33, 425) <= 0; flappy_W(33, 426) <= 1; flappy_W(33, 427) <= 1; flappy_W(33, 428) <= 1; flappy_W(33, 429) <= 1; flappy_W(33, 430) <= 1; flappy_W(33, 431) <= 1; flappy_W(33, 432) <= 1; flappy_W(33, 433) <= 1; flappy_W(33, 434) <= 1; flappy_W(33, 435) <= 1; flappy_W(33, 436) <= 1; flappy_W(33, 437) <= 1; flappy_W(33, 438) <= 0; flappy_W(33, 439) <= 0; flappy_W(33, 440) <= 0; flappy_W(33, 441) <= 0; flappy_W(33, 442) <= 0; flappy_W(33, 443) <= 0; flappy_W(33, 444) <= 0; flappy_W(33, 445) <= 0; flappy_W(33, 446) <= 0; flappy_W(33, 447) <= 0; flappy_W(33, 448) <= 0; flappy_W(33, 449) <= 0; flappy_W(33, 450) <= 0; flappy_W(33, 451) <= 0; flappy_W(33, 452) <= 0; flappy_W(33, 453) <= 0; flappy_W(33, 454) <= 0; flappy_W(33, 455) <= 0; flappy_W(33, 456) <= 0; flappy_W(33, 457) <= 0; flappy_W(33, 458) <= 0; flappy_W(33, 459) <= 0; flappy_W(33, 460) <= 0; flappy_W(33, 461) <= 0; flappy_W(33, 462) <= 0; flappy_W(33, 463) <= 0; flappy_W(33, 464) <= 0; flappy_W(33, 465) <= 0; flappy_W(33, 466) <= 0; flappy_W(33, 467) <= 0; flappy_W(33, 468) <= 1; flappy_W(33, 469) <= 1; flappy_W(33, 470) <= 1; flappy_W(33, 471) <= 1; flappy_W(33, 472) <= 1; flappy_W(33, 473) <= 1; flappy_W(33, 474) <= 1; flappy_W(33, 475) <= 1; flappy_W(33, 476) <= 1; flappy_W(33, 477) <= 1; flappy_W(33, 478) <= 1; flappy_W(33, 479) <= 1; flappy_W(33, 480) <= 0; flappy_W(33, 481) <= 0; flappy_W(33, 482) <= 0; flappy_W(33, 483) <= 0; flappy_W(33, 484) <= 0; flappy_W(33, 485) <= 0; flappy_W(33, 486) <= 0; flappy_W(33, 487) <= 0; flappy_W(33, 488) <= 0; flappy_W(33, 489) <= 0; flappy_W(33, 490) <= 0; flappy_W(33, 491) <= 0; flappy_W(33, 492) <= 0; flappy_W(33, 493) <= 0; flappy_W(33, 494) <= 0; flappy_W(33, 495) <= 0; flappy_W(33, 496) <= 0; flappy_W(33, 497) <= 0; flappy_W(33, 498) <= 0; flappy_W(33, 499) <= 0; flappy_W(33, 500) <= 0; flappy_W(33, 501) <= 0; flappy_W(33, 502) <= 0; flappy_W(33, 503) <= 0; flappy_W(33, 504) <= 0; flappy_W(33, 505) <= 0; flappy_W(33, 506) <= 0; flappy_W(33, 507) <= 0; flappy_W(33, 508) <= 0; flappy_W(33, 509) <= 0; flappy_W(33, 510) <= 1; flappy_W(33, 511) <= 1; flappy_W(33, 512) <= 1; flappy_W(33, 513) <= 1; flappy_W(33, 514) <= 1; flappy_W(33, 515) <= 1; flappy_W(33, 516) <= 1; flappy_W(33, 517) <= 1; flappy_W(33, 518) <= 1; flappy_W(33, 519) <= 1; flappy_W(33, 520) <= 1; flappy_W(33, 521) <= 1; flappy_W(33, 522) <= 0; flappy_W(33, 523) <= 0; flappy_W(33, 524) <= 0; flappy_W(33, 525) <= 0; flappy_W(33, 526) <= 0; flappy_W(33, 527) <= 0; flappy_W(33, 528) <= 1; flappy_W(33, 529) <= 1; flappy_W(33, 530) <= 1; flappy_W(33, 531) <= 1; flappy_W(33, 532) <= 1; flappy_W(33, 533) <= 1; flappy_W(33, 534) <= 1; flappy_W(33, 535) <= 1; flappy_W(33, 536) <= 1; flappy_W(33, 537) <= 1; flappy_W(33, 538) <= 1; flappy_W(33, 539) <= 1; flappy_W(33, 540) <= 0; flappy_W(33, 541) <= 0; flappy_W(33, 542) <= 0; flappy_W(33, 543) <= 0; flappy_W(33, 544) <= 0; flappy_W(33, 545) <= 0; flappy_W(33, 546) <= 0; flappy_W(33, 547) <= 0; flappy_W(33, 548) <= 0; flappy_W(33, 549) <= 0; flappy_W(33, 550) <= 0; flappy_W(33, 551) <= 0; flappy_W(33, 552) <= 0; flappy_W(33, 553) <= 0; flappy_W(33, 554) <= 0; flappy_W(33, 555) <= 0; flappy_W(33, 556) <= 0; flappy_W(33, 557) <= 0; flappy_W(33, 558) <= 0; flappy_W(33, 559) <= 0; flappy_W(33, 560) <= 0; flappy_W(33, 561) <= 0; flappy_W(33, 562) <= 0; flappy_W(33, 563) <= 0; flappy_W(33, 564) <= 1; flappy_W(33, 565) <= 1; flappy_W(33, 566) <= 1; flappy_W(33, 567) <= 1; flappy_W(33, 568) <= 1; flappy_W(33, 569) <= 1; flappy_W(33, 570) <= 1; flappy_W(33, 571) <= 1; flappy_W(33, 572) <= 1; flappy_W(33, 573) <= 1; flappy_W(33, 574) <= 1; flappy_W(33, 575) <= 1; flappy_W(33, 576) <= 0; flappy_W(33, 577) <= 0; flappy_W(33, 578) <= 0; flappy_W(33, 579) <= 0; flappy_W(33, 580) <= 0; flappy_W(33, 581) <= 0; flappy_W(33, 582) <= 0; flappy_W(33, 583) <= 0; flappy_W(33, 584) <= 0; flappy_W(33, 585) <= 0; flappy_W(33, 586) <= 0; flappy_W(33, 587) <= 0; flappy_W(33, 588) <= 1; flappy_W(33, 589) <= 1; flappy_W(33, 590) <= 1; flappy_W(33, 591) <= 1; flappy_W(33, 592) <= 1; flappy_W(33, 593) <= 1; 
flappy_W(34, 0) <= 0; flappy_W(34, 1) <= 0; flappy_W(34, 2) <= 0; flappy_W(34, 3) <= 0; flappy_W(34, 4) <= 0; flappy_W(34, 5) <= 0; flappy_W(34, 6) <= 1; flappy_W(34, 7) <= 1; flappy_W(34, 8) <= 1; flappy_W(34, 9) <= 1; flappy_W(34, 10) <= 1; flappy_W(34, 11) <= 1; flappy_W(34, 12) <= 1; flappy_W(34, 13) <= 1; flappy_W(34, 14) <= 1; flappy_W(34, 15) <= 1; flappy_W(34, 16) <= 1; flappy_W(34, 17) <= 1; flappy_W(34, 18) <= 0; flappy_W(34, 19) <= 0; flappy_W(34, 20) <= 0; flappy_W(34, 21) <= 0; flappy_W(34, 22) <= 0; flappy_W(34, 23) <= 0; flappy_W(34, 24) <= 1; flappy_W(34, 25) <= 1; flappy_W(34, 26) <= 1; flappy_W(34, 27) <= 1; flappy_W(34, 28) <= 1; flappy_W(34, 29) <= 1; flappy_W(34, 30) <= 0; flappy_W(34, 31) <= 0; flappy_W(34, 32) <= 0; flappy_W(34, 33) <= 0; flappy_W(34, 34) <= 0; flappy_W(34, 35) <= 0; flappy_W(34, 36) <= 0; flappy_W(34, 37) <= 0; flappy_W(34, 38) <= 0; flappy_W(34, 39) <= 0; flappy_W(34, 40) <= 0; flappy_W(34, 41) <= 0; flappy_W(34, 42) <= 0; flappy_W(34, 43) <= 0; flappy_W(34, 44) <= 0; flappy_W(34, 45) <= 0; flappy_W(34, 46) <= 0; flappy_W(34, 47) <= 0; flappy_W(34, 48) <= 0; flappy_W(34, 49) <= 0; flappy_W(34, 50) <= 0; flappy_W(34, 51) <= 0; flappy_W(34, 52) <= 0; flappy_W(34, 53) <= 0; flappy_W(34, 54) <= 0; flappy_W(34, 55) <= 0; flappy_W(34, 56) <= 0; flappy_W(34, 57) <= 0; flappy_W(34, 58) <= 0; flappy_W(34, 59) <= 0; flappy_W(34, 60) <= 1; flappy_W(34, 61) <= 1; flappy_W(34, 62) <= 1; flappy_W(34, 63) <= 1; flappy_W(34, 64) <= 1; flappy_W(34, 65) <= 1; flappy_W(34, 66) <= 1; flappy_W(34, 67) <= 1; flappy_W(34, 68) <= 1; flappy_W(34, 69) <= 1; flappy_W(34, 70) <= 1; flappy_W(34, 71) <= 1; flappy_W(34, 72) <= 0; flappy_W(34, 73) <= 0; flappy_W(34, 74) <= 0; flappy_W(34, 75) <= 0; flappy_W(34, 76) <= 0; flappy_W(34, 77) <= 0; flappy_W(34, 78) <= 0; flappy_W(34, 79) <= 0; flappy_W(34, 80) <= 0; flappy_W(34, 81) <= 0; flappy_W(34, 82) <= 0; flappy_W(34, 83) <= 0; flappy_W(34, 84) <= 0; flappy_W(34, 85) <= 0; flappy_W(34, 86) <= 0; flappy_W(34, 87) <= 0; flappy_W(34, 88) <= 0; flappy_W(34, 89) <= 0; flappy_W(34, 90) <= 0; flappy_W(34, 91) <= 0; flappy_W(34, 92) <= 0; flappy_W(34, 93) <= 0; flappy_W(34, 94) <= 0; flappy_W(34, 95) <= 0; flappy_W(34, 96) <= 0; flappy_W(34, 97) <= 0; flappy_W(34, 98) <= 0; flappy_W(34, 99) <= 0; flappy_W(34, 100) <= 0; flappy_W(34, 101) <= 0; flappy_W(34, 102) <= 0; flappy_W(34, 103) <= 0; flappy_W(34, 104) <= 0; flappy_W(34, 105) <= 0; flappy_W(34, 106) <= 0; flappy_W(34, 107) <= 0; flappy_W(34, 108) <= 1; flappy_W(34, 109) <= 1; flappy_W(34, 110) <= 1; flappy_W(34, 111) <= 1; flappy_W(34, 112) <= 1; flappy_W(34, 113) <= 1; flappy_W(34, 114) <= 1; flappy_W(34, 115) <= 1; flappy_W(34, 116) <= 1; flappy_W(34, 117) <= 1; flappy_W(34, 118) <= 1; flappy_W(34, 119) <= 1; flappy_W(34, 120) <= 1; flappy_W(34, 121) <= 1; flappy_W(34, 122) <= 1; flappy_W(34, 123) <= 1; flappy_W(34, 124) <= 1; flappy_W(34, 125) <= 1; flappy_W(34, 126) <= 1; flappy_W(34, 127) <= 1; flappy_W(34, 128) <= 1; flappy_W(34, 129) <= 1; flappy_W(34, 130) <= 1; flappy_W(34, 131) <= 1; flappy_W(34, 132) <= 1; flappy_W(34, 133) <= 1; flappy_W(34, 134) <= 1; flappy_W(34, 135) <= 1; flappy_W(34, 136) <= 1; flappy_W(34, 137) <= 1; flappy_W(34, 138) <= 1; flappy_W(34, 139) <= 1; flappy_W(34, 140) <= 1; flappy_W(34, 141) <= 1; flappy_W(34, 142) <= 1; flappy_W(34, 143) <= 1; flappy_W(34, 144) <= 1; flappy_W(34, 145) <= 1; flappy_W(34, 146) <= 1; flappy_W(34, 147) <= 1; flappy_W(34, 148) <= 1; flappy_W(34, 149) <= 1; flappy_W(34, 150) <= 0; flappy_W(34, 151) <= 0; flappy_W(34, 152) <= 0; flappy_W(34, 153) <= 0; flappy_W(34, 154) <= 0; flappy_W(34, 155) <= 0; flappy_W(34, 156) <= 0; flappy_W(34, 157) <= 0; flappy_W(34, 158) <= 0; flappy_W(34, 159) <= 0; flappy_W(34, 160) <= 0; flappy_W(34, 161) <= 0; flappy_W(34, 162) <= 0; flappy_W(34, 163) <= 0; flappy_W(34, 164) <= 0; flappy_W(34, 165) <= 0; flappy_W(34, 166) <= 0; flappy_W(34, 167) <= 0; flappy_W(34, 168) <= 1; flappy_W(34, 169) <= 1; flappy_W(34, 170) <= 1; flappy_W(34, 171) <= 1; flappy_W(34, 172) <= 1; flappy_W(34, 173) <= 1; flappy_W(34, 174) <= 1; flappy_W(34, 175) <= 1; flappy_W(34, 176) <= 1; flappy_W(34, 177) <= 1; flappy_W(34, 178) <= 1; flappy_W(34, 179) <= 1; flappy_W(34, 180) <= 0; flappy_W(34, 181) <= 0; flappy_W(34, 182) <= 0; flappy_W(34, 183) <= 0; flappy_W(34, 184) <= 0; flappy_W(34, 185) <= 0; flappy_W(34, 186) <= 0; flappy_W(34, 187) <= 0; flappy_W(34, 188) <= 0; flappy_W(34, 189) <= 0; flappy_W(34, 190) <= 0; flappy_W(34, 191) <= 0; flappy_W(34, 192) <= 0; flappy_W(34, 193) <= 0; flappy_W(34, 194) <= 0; flappy_W(34, 195) <= 0; flappy_W(34, 196) <= 0; flappy_W(34, 197) <= 0; flappy_W(34, 198) <= 0; flappy_W(34, 199) <= 0; flappy_W(34, 200) <= 0; flappy_W(34, 201) <= 0; flappy_W(34, 202) <= 0; flappy_W(34, 203) <= 0; flappy_W(34, 204) <= 0; flappy_W(34, 205) <= 0; flappy_W(34, 206) <= 0; flappy_W(34, 207) <= 0; flappy_W(34, 208) <= 0; flappy_W(34, 209) <= 0; flappy_W(34, 210) <= 0; flappy_W(34, 211) <= 0; flappy_W(34, 212) <= 0; flappy_W(34, 213) <= 0; flappy_W(34, 214) <= 0; flappy_W(34, 215) <= 0; flappy_W(34, 216) <= 0; flappy_W(34, 217) <= 0; flappy_W(34, 218) <= 0; flappy_W(34, 219) <= 0; flappy_W(34, 220) <= 0; flappy_W(34, 221) <= 0; flappy_W(34, 222) <= 1; flappy_W(34, 223) <= 1; flappy_W(34, 224) <= 1; flappy_W(34, 225) <= 1; flappy_W(34, 226) <= 1; flappy_W(34, 227) <= 1; flappy_W(34, 228) <= 1; flappy_W(34, 229) <= 1; flappy_W(34, 230) <= 1; flappy_W(34, 231) <= 1; flappy_W(34, 232) <= 1; flappy_W(34, 233) <= 1; flappy_W(34, 234) <= 0; flappy_W(34, 235) <= 0; flappy_W(34, 236) <= 0; flappy_W(34, 237) <= 0; flappy_W(34, 238) <= 0; flappy_W(34, 239) <= 0; flappy_W(34, 240) <= 0; flappy_W(34, 241) <= 0; flappy_W(34, 242) <= 0; flappy_W(34, 243) <= 0; flappy_W(34, 244) <= 0; flappy_W(34, 245) <= 0; flappy_W(34, 246) <= 0; flappy_W(34, 247) <= 0; flappy_W(34, 248) <= 0; flappy_W(34, 249) <= 0; flappy_W(34, 250) <= 0; flappy_W(34, 251) <= 0; flappy_W(34, 252) <= 0; flappy_W(34, 253) <= 0; flappy_W(34, 254) <= 0; flappy_W(34, 255) <= 0; flappy_W(34, 256) <= 0; flappy_W(34, 257) <= 0; flappy_W(34, 258) <= 0; flappy_W(34, 259) <= 0; flappy_W(34, 260) <= 0; flappy_W(34, 261) <= 0; flappy_W(34, 262) <= 0; flappy_W(34, 263) <= 0; flappy_W(34, 264) <= 0; flappy_W(34, 265) <= 0; flappy_W(34, 266) <= 0; flappy_W(34, 267) <= 0; flappy_W(34, 268) <= 0; flappy_W(34, 269) <= 0; flappy_W(34, 270) <= 0; flappy_W(34, 271) <= 0; flappy_W(34, 272) <= 0; flappy_W(34, 273) <= 0; flappy_W(34, 274) <= 0; flappy_W(34, 275) <= 0; flappy_W(34, 276) <= 0; flappy_W(34, 277) <= 0; flappy_W(34, 278) <= 0; flappy_W(34, 279) <= 0; flappy_W(34, 280) <= 0; flappy_W(34, 281) <= 0; flappy_W(34, 282) <= 0; flappy_W(34, 283) <= 0; flappy_W(34, 284) <= 0; flappy_W(34, 285) <= 0; flappy_W(34, 286) <= 0; flappy_W(34, 287) <= 0; flappy_W(34, 288) <= 1; flappy_W(34, 289) <= 1; flappy_W(34, 290) <= 1; flappy_W(34, 291) <= 1; flappy_W(34, 292) <= 1; flappy_W(34, 293) <= 1; flappy_W(34, 294) <= 1; flappy_W(34, 295) <= 1; flappy_W(34, 296) <= 1; flappy_W(34, 297) <= 1; flappy_W(34, 298) <= 1; flappy_W(34, 299) <= 1; flappy_W(34, 300) <= 0; flappy_W(34, 301) <= 0; flappy_W(34, 302) <= 0; flappy_W(34, 303) <= 0; flappy_W(34, 304) <= 0; flappy_W(34, 305) <= 0; flappy_W(34, 306) <= 0; flappy_W(34, 307) <= 0; flappy_W(34, 308) <= 0; flappy_W(34, 309) <= 0; flappy_W(34, 310) <= 0; flappy_W(34, 311) <= 0; flappy_W(34, 312) <= 0; flappy_W(34, 313) <= 0; flappy_W(34, 314) <= 0; flappy_W(34, 315) <= 0; flappy_W(34, 316) <= 0; flappy_W(34, 317) <= 0; flappy_W(34, 318) <= 0; flappy_W(34, 319) <= 0; flappy_W(34, 320) <= 0; flappy_W(34, 321) <= 0; flappy_W(34, 322) <= 0; flappy_W(34, 323) <= 0; flappy_W(34, 324) <= 0; flappy_W(34, 325) <= 0; flappy_W(34, 326) <= 0; flappy_W(34, 327) <= 0; flappy_W(34, 328) <= 0; flappy_W(34, 329) <= 0; flappy_W(34, 330) <= 0; flappy_W(34, 331) <= 0; flappy_W(34, 332) <= 0; flappy_W(34, 333) <= 0; flappy_W(34, 334) <= 0; flappy_W(34, 335) <= 0; flappy_W(34, 336) <= 0; flappy_W(34, 337) <= 0; flappy_W(34, 338) <= 0; flappy_W(34, 339) <= 0; flappy_W(34, 340) <= 0; flappy_W(34, 341) <= 0; flappy_W(34, 342) <= 0; flappy_W(34, 343) <= 0; flappy_W(34, 344) <= 0; flappy_W(34, 345) <= 0; flappy_W(34, 346) <= 0; flappy_W(34, 347) <= 0; flappy_W(34, 348) <= 0; flappy_W(34, 349) <= 0; flappy_W(34, 350) <= 0; flappy_W(34, 351) <= 0; flappy_W(34, 352) <= 0; flappy_W(34, 353) <= 0; flappy_W(34, 354) <= 0; flappy_W(34, 355) <= 0; flappy_W(34, 356) <= 0; flappy_W(34, 357) <= 0; flappy_W(34, 358) <= 0; flappy_W(34, 359) <= 0; flappy_W(34, 360) <= 0; flappy_W(34, 361) <= 0; flappy_W(34, 362) <= 0; flappy_W(34, 363) <= 0; flappy_W(34, 364) <= 0; flappy_W(34, 365) <= 0; flappy_W(34, 366) <= 0; flappy_W(34, 367) <= 0; flappy_W(34, 368) <= 0; flappy_W(34, 369) <= 0; flappy_W(34, 370) <= 0; flappy_W(34, 371) <= 0; flappy_W(34, 372) <= 0; flappy_W(34, 373) <= 0; flappy_W(34, 374) <= 0; flappy_W(34, 375) <= 0; flappy_W(34, 376) <= 0; flappy_W(34, 377) <= 0; flappy_W(34, 378) <= 0; flappy_W(34, 379) <= 0; flappy_W(34, 380) <= 0; flappy_W(34, 381) <= 0; flappy_W(34, 382) <= 0; flappy_W(34, 383) <= 0; flappy_W(34, 384) <= 0; flappy_W(34, 385) <= 0; flappy_W(34, 386) <= 0; flappy_W(34, 387) <= 0; flappy_W(34, 388) <= 0; flappy_W(34, 389) <= 0; flappy_W(34, 390) <= 0; flappy_W(34, 391) <= 0; flappy_W(34, 392) <= 0; flappy_W(34, 393) <= 0; flappy_W(34, 394) <= 0; flappy_W(34, 395) <= 0; flappy_W(34, 396) <= 0; flappy_W(34, 397) <= 0; flappy_W(34, 398) <= 0; flappy_W(34, 399) <= 0; flappy_W(34, 400) <= 0; flappy_W(34, 401) <= 0; flappy_W(34, 402) <= 1; flappy_W(34, 403) <= 1; flappy_W(34, 404) <= 1; flappy_W(34, 405) <= 1; flappy_W(34, 406) <= 1; flappy_W(34, 407) <= 1; flappy_W(34, 408) <= 1; flappy_W(34, 409) <= 1; flappy_W(34, 410) <= 1; flappy_W(34, 411) <= 1; flappy_W(34, 412) <= 1; flappy_W(34, 413) <= 1; flappy_W(34, 414) <= 0; flappy_W(34, 415) <= 0; flappy_W(34, 416) <= 0; flappy_W(34, 417) <= 0; flappy_W(34, 418) <= 0; flappy_W(34, 419) <= 0; flappy_W(34, 420) <= 0; flappy_W(34, 421) <= 0; flappy_W(34, 422) <= 0; flappy_W(34, 423) <= 0; flappy_W(34, 424) <= 0; flappy_W(34, 425) <= 0; flappy_W(34, 426) <= 1; flappy_W(34, 427) <= 1; flappy_W(34, 428) <= 1; flappy_W(34, 429) <= 1; flappy_W(34, 430) <= 1; flappy_W(34, 431) <= 1; flappy_W(34, 432) <= 1; flappy_W(34, 433) <= 1; flappy_W(34, 434) <= 1; flappy_W(34, 435) <= 1; flappy_W(34, 436) <= 1; flappy_W(34, 437) <= 1; flappy_W(34, 438) <= 0; flappy_W(34, 439) <= 0; flappy_W(34, 440) <= 0; flappy_W(34, 441) <= 0; flappy_W(34, 442) <= 0; flappy_W(34, 443) <= 0; flappy_W(34, 444) <= 0; flappy_W(34, 445) <= 0; flappy_W(34, 446) <= 0; flappy_W(34, 447) <= 0; flappy_W(34, 448) <= 0; flappy_W(34, 449) <= 0; flappy_W(34, 450) <= 0; flappy_W(34, 451) <= 0; flappy_W(34, 452) <= 0; flappy_W(34, 453) <= 0; flappy_W(34, 454) <= 0; flappy_W(34, 455) <= 0; flappy_W(34, 456) <= 0; flappy_W(34, 457) <= 0; flappy_W(34, 458) <= 0; flappy_W(34, 459) <= 0; flappy_W(34, 460) <= 0; flappy_W(34, 461) <= 0; flappy_W(34, 462) <= 0; flappy_W(34, 463) <= 0; flappy_W(34, 464) <= 0; flappy_W(34, 465) <= 0; flappy_W(34, 466) <= 0; flappy_W(34, 467) <= 0; flappy_W(34, 468) <= 1; flappy_W(34, 469) <= 1; flappy_W(34, 470) <= 1; flappy_W(34, 471) <= 1; flappy_W(34, 472) <= 1; flappy_W(34, 473) <= 1; flappy_W(34, 474) <= 1; flappy_W(34, 475) <= 1; flappy_W(34, 476) <= 1; flappy_W(34, 477) <= 1; flappy_W(34, 478) <= 1; flappy_W(34, 479) <= 1; flappy_W(34, 480) <= 0; flappy_W(34, 481) <= 0; flappy_W(34, 482) <= 0; flappy_W(34, 483) <= 0; flappy_W(34, 484) <= 0; flappy_W(34, 485) <= 0; flappy_W(34, 486) <= 0; flappy_W(34, 487) <= 0; flappy_W(34, 488) <= 0; flappy_W(34, 489) <= 0; flappy_W(34, 490) <= 0; flappy_W(34, 491) <= 0; flappy_W(34, 492) <= 0; flappy_W(34, 493) <= 0; flappy_W(34, 494) <= 0; flappy_W(34, 495) <= 0; flappy_W(34, 496) <= 0; flappy_W(34, 497) <= 0; flappy_W(34, 498) <= 0; flappy_W(34, 499) <= 0; flappy_W(34, 500) <= 0; flappy_W(34, 501) <= 0; flappy_W(34, 502) <= 0; flappy_W(34, 503) <= 0; flappy_W(34, 504) <= 0; flappy_W(34, 505) <= 0; flappy_W(34, 506) <= 0; flappy_W(34, 507) <= 0; flappy_W(34, 508) <= 0; flappy_W(34, 509) <= 0; flappy_W(34, 510) <= 1; flappy_W(34, 511) <= 1; flappy_W(34, 512) <= 1; flappy_W(34, 513) <= 1; flappy_W(34, 514) <= 1; flappy_W(34, 515) <= 1; flappy_W(34, 516) <= 1; flappy_W(34, 517) <= 1; flappy_W(34, 518) <= 1; flappy_W(34, 519) <= 1; flappy_W(34, 520) <= 1; flappy_W(34, 521) <= 1; flappy_W(34, 522) <= 0; flappy_W(34, 523) <= 0; flappy_W(34, 524) <= 0; flappy_W(34, 525) <= 0; flappy_W(34, 526) <= 0; flappy_W(34, 527) <= 0; flappy_W(34, 528) <= 1; flappy_W(34, 529) <= 1; flappy_W(34, 530) <= 1; flappy_W(34, 531) <= 1; flappy_W(34, 532) <= 1; flappy_W(34, 533) <= 1; flappy_W(34, 534) <= 1; flappy_W(34, 535) <= 1; flappy_W(34, 536) <= 1; flappy_W(34, 537) <= 1; flappy_W(34, 538) <= 1; flappy_W(34, 539) <= 1; flappy_W(34, 540) <= 0; flappy_W(34, 541) <= 0; flappy_W(34, 542) <= 0; flappy_W(34, 543) <= 0; flappy_W(34, 544) <= 0; flappy_W(34, 545) <= 0; flappy_W(34, 546) <= 0; flappy_W(34, 547) <= 0; flappy_W(34, 548) <= 0; flappy_W(34, 549) <= 0; flappy_W(34, 550) <= 0; flappy_W(34, 551) <= 0; flappy_W(34, 552) <= 0; flappy_W(34, 553) <= 0; flappy_W(34, 554) <= 0; flappy_W(34, 555) <= 0; flappy_W(34, 556) <= 0; flappy_W(34, 557) <= 0; flappy_W(34, 558) <= 0; flappy_W(34, 559) <= 0; flappy_W(34, 560) <= 0; flappy_W(34, 561) <= 0; flappy_W(34, 562) <= 0; flappy_W(34, 563) <= 0; flappy_W(34, 564) <= 1; flappy_W(34, 565) <= 1; flappy_W(34, 566) <= 1; flappy_W(34, 567) <= 1; flappy_W(34, 568) <= 1; flappy_W(34, 569) <= 1; flappy_W(34, 570) <= 1; flappy_W(34, 571) <= 1; flappy_W(34, 572) <= 1; flappy_W(34, 573) <= 1; flappy_W(34, 574) <= 1; flappy_W(34, 575) <= 1; flappy_W(34, 576) <= 0; flappy_W(34, 577) <= 0; flappy_W(34, 578) <= 0; flappy_W(34, 579) <= 0; flappy_W(34, 580) <= 0; flappy_W(34, 581) <= 0; flappy_W(34, 582) <= 0; flappy_W(34, 583) <= 0; flappy_W(34, 584) <= 0; flappy_W(34, 585) <= 0; flappy_W(34, 586) <= 0; flappy_W(34, 587) <= 0; flappy_W(34, 588) <= 1; flappy_W(34, 589) <= 1; flappy_W(34, 590) <= 1; flappy_W(34, 591) <= 1; flappy_W(34, 592) <= 1; flappy_W(34, 593) <= 1; 
flappy_W(35, 0) <= 0; flappy_W(35, 1) <= 0; flappy_W(35, 2) <= 0; flappy_W(35, 3) <= 0; flappy_W(35, 4) <= 0; flappy_W(35, 5) <= 0; flappy_W(35, 6) <= 1; flappy_W(35, 7) <= 1; flappy_W(35, 8) <= 1; flappy_W(35, 9) <= 1; flappy_W(35, 10) <= 1; flappy_W(35, 11) <= 1; flappy_W(35, 12) <= 1; flappy_W(35, 13) <= 1; flappy_W(35, 14) <= 1; flappy_W(35, 15) <= 1; flappy_W(35, 16) <= 1; flappy_W(35, 17) <= 1; flappy_W(35, 18) <= 0; flappy_W(35, 19) <= 0; flappy_W(35, 20) <= 0; flappy_W(35, 21) <= 0; flappy_W(35, 22) <= 0; flappy_W(35, 23) <= 0; flappy_W(35, 24) <= 1; flappy_W(35, 25) <= 1; flappy_W(35, 26) <= 1; flappy_W(35, 27) <= 1; flappy_W(35, 28) <= 1; flappy_W(35, 29) <= 1; flappy_W(35, 30) <= 0; flappy_W(35, 31) <= 0; flappy_W(35, 32) <= 0; flappy_W(35, 33) <= 0; flappy_W(35, 34) <= 0; flappy_W(35, 35) <= 0; flappy_W(35, 36) <= 0; flappy_W(35, 37) <= 0; flappy_W(35, 38) <= 0; flappy_W(35, 39) <= 0; flappy_W(35, 40) <= 0; flappy_W(35, 41) <= 0; flappy_W(35, 42) <= 0; flappy_W(35, 43) <= 0; flappy_W(35, 44) <= 0; flappy_W(35, 45) <= 0; flappy_W(35, 46) <= 0; flappy_W(35, 47) <= 0; flappy_W(35, 48) <= 0; flappy_W(35, 49) <= 0; flappy_W(35, 50) <= 0; flappy_W(35, 51) <= 0; flappy_W(35, 52) <= 0; flappy_W(35, 53) <= 0; flappy_W(35, 54) <= 0; flappy_W(35, 55) <= 0; flappy_W(35, 56) <= 0; flappy_W(35, 57) <= 0; flappy_W(35, 58) <= 0; flappy_W(35, 59) <= 0; flappy_W(35, 60) <= 1; flappy_W(35, 61) <= 1; flappy_W(35, 62) <= 1; flappy_W(35, 63) <= 1; flappy_W(35, 64) <= 1; flappy_W(35, 65) <= 1; flappy_W(35, 66) <= 1; flappy_W(35, 67) <= 1; flappy_W(35, 68) <= 1; flappy_W(35, 69) <= 1; flappy_W(35, 70) <= 1; flappy_W(35, 71) <= 1; flappy_W(35, 72) <= 0; flappy_W(35, 73) <= 0; flappy_W(35, 74) <= 0; flappy_W(35, 75) <= 0; flappy_W(35, 76) <= 0; flappy_W(35, 77) <= 0; flappy_W(35, 78) <= 0; flappy_W(35, 79) <= 0; flappy_W(35, 80) <= 0; flappy_W(35, 81) <= 0; flappy_W(35, 82) <= 0; flappy_W(35, 83) <= 0; flappy_W(35, 84) <= 0; flappy_W(35, 85) <= 0; flappy_W(35, 86) <= 0; flappy_W(35, 87) <= 0; flappy_W(35, 88) <= 0; flappy_W(35, 89) <= 0; flappy_W(35, 90) <= 0; flappy_W(35, 91) <= 0; flappy_W(35, 92) <= 0; flappy_W(35, 93) <= 0; flappy_W(35, 94) <= 0; flappy_W(35, 95) <= 0; flappy_W(35, 96) <= 0; flappy_W(35, 97) <= 0; flappy_W(35, 98) <= 0; flappy_W(35, 99) <= 0; flappy_W(35, 100) <= 0; flappy_W(35, 101) <= 0; flappy_W(35, 102) <= 0; flappy_W(35, 103) <= 0; flappy_W(35, 104) <= 0; flappy_W(35, 105) <= 0; flappy_W(35, 106) <= 0; flappy_W(35, 107) <= 0; flappy_W(35, 108) <= 1; flappy_W(35, 109) <= 1; flappy_W(35, 110) <= 1; flappy_W(35, 111) <= 1; flappy_W(35, 112) <= 1; flappy_W(35, 113) <= 1; flappy_W(35, 114) <= 1; flappy_W(35, 115) <= 1; flappy_W(35, 116) <= 1; flappy_W(35, 117) <= 1; flappy_W(35, 118) <= 1; flappy_W(35, 119) <= 1; flappy_W(35, 120) <= 1; flappy_W(35, 121) <= 1; flappy_W(35, 122) <= 1; flappy_W(35, 123) <= 1; flappy_W(35, 124) <= 1; flappy_W(35, 125) <= 1; flappy_W(35, 126) <= 1; flappy_W(35, 127) <= 1; flappy_W(35, 128) <= 1; flappy_W(35, 129) <= 1; flappy_W(35, 130) <= 1; flappy_W(35, 131) <= 1; flappy_W(35, 132) <= 1; flappy_W(35, 133) <= 1; flappy_W(35, 134) <= 1; flappy_W(35, 135) <= 1; flappy_W(35, 136) <= 1; flappy_W(35, 137) <= 1; flappy_W(35, 138) <= 1; flappy_W(35, 139) <= 1; flappy_W(35, 140) <= 1; flappy_W(35, 141) <= 1; flappy_W(35, 142) <= 1; flappy_W(35, 143) <= 1; flappy_W(35, 144) <= 1; flappy_W(35, 145) <= 1; flappy_W(35, 146) <= 1; flappy_W(35, 147) <= 1; flappy_W(35, 148) <= 1; flappy_W(35, 149) <= 1; flappy_W(35, 150) <= 0; flappy_W(35, 151) <= 0; flappy_W(35, 152) <= 0; flappy_W(35, 153) <= 0; flappy_W(35, 154) <= 0; flappy_W(35, 155) <= 0; flappy_W(35, 156) <= 0; flappy_W(35, 157) <= 0; flappy_W(35, 158) <= 0; flappy_W(35, 159) <= 0; flappy_W(35, 160) <= 0; flappy_W(35, 161) <= 0; flappy_W(35, 162) <= 0; flappy_W(35, 163) <= 0; flappy_W(35, 164) <= 0; flappy_W(35, 165) <= 0; flappy_W(35, 166) <= 0; flappy_W(35, 167) <= 0; flappy_W(35, 168) <= 1; flappy_W(35, 169) <= 1; flappy_W(35, 170) <= 1; flappy_W(35, 171) <= 1; flappy_W(35, 172) <= 1; flappy_W(35, 173) <= 1; flappy_W(35, 174) <= 1; flappy_W(35, 175) <= 1; flappy_W(35, 176) <= 1; flappy_W(35, 177) <= 1; flappy_W(35, 178) <= 1; flappy_W(35, 179) <= 1; flappy_W(35, 180) <= 0; flappy_W(35, 181) <= 0; flappy_W(35, 182) <= 0; flappy_W(35, 183) <= 0; flappy_W(35, 184) <= 0; flappy_W(35, 185) <= 0; flappy_W(35, 186) <= 0; flappy_W(35, 187) <= 0; flappy_W(35, 188) <= 0; flappy_W(35, 189) <= 0; flappy_W(35, 190) <= 0; flappy_W(35, 191) <= 0; flappy_W(35, 192) <= 0; flappy_W(35, 193) <= 0; flappy_W(35, 194) <= 0; flappy_W(35, 195) <= 0; flappy_W(35, 196) <= 0; flappy_W(35, 197) <= 0; flappy_W(35, 198) <= 0; flappy_W(35, 199) <= 0; flappy_W(35, 200) <= 0; flappy_W(35, 201) <= 0; flappy_W(35, 202) <= 0; flappy_W(35, 203) <= 0; flappy_W(35, 204) <= 0; flappy_W(35, 205) <= 0; flappy_W(35, 206) <= 0; flappy_W(35, 207) <= 0; flappy_W(35, 208) <= 0; flappy_W(35, 209) <= 0; flappy_W(35, 210) <= 0; flappy_W(35, 211) <= 0; flappy_W(35, 212) <= 0; flappy_W(35, 213) <= 0; flappy_W(35, 214) <= 0; flappy_W(35, 215) <= 0; flappy_W(35, 216) <= 0; flappy_W(35, 217) <= 0; flappy_W(35, 218) <= 0; flappy_W(35, 219) <= 0; flappy_W(35, 220) <= 0; flappy_W(35, 221) <= 0; flappy_W(35, 222) <= 1; flappy_W(35, 223) <= 1; flappy_W(35, 224) <= 1; flappy_W(35, 225) <= 1; flappy_W(35, 226) <= 1; flappy_W(35, 227) <= 1; flappy_W(35, 228) <= 1; flappy_W(35, 229) <= 1; flappy_W(35, 230) <= 1; flappy_W(35, 231) <= 1; flappy_W(35, 232) <= 1; flappy_W(35, 233) <= 1; flappy_W(35, 234) <= 0; flappy_W(35, 235) <= 0; flappy_W(35, 236) <= 0; flappy_W(35, 237) <= 0; flappy_W(35, 238) <= 0; flappy_W(35, 239) <= 0; flappy_W(35, 240) <= 0; flappy_W(35, 241) <= 0; flappy_W(35, 242) <= 0; flappy_W(35, 243) <= 0; flappy_W(35, 244) <= 0; flappy_W(35, 245) <= 0; flappy_W(35, 246) <= 0; flappy_W(35, 247) <= 0; flappy_W(35, 248) <= 0; flappy_W(35, 249) <= 0; flappy_W(35, 250) <= 0; flappy_W(35, 251) <= 0; flappy_W(35, 252) <= 0; flappy_W(35, 253) <= 0; flappy_W(35, 254) <= 0; flappy_W(35, 255) <= 0; flappy_W(35, 256) <= 0; flappy_W(35, 257) <= 0; flappy_W(35, 258) <= 0; flappy_W(35, 259) <= 0; flappy_W(35, 260) <= 0; flappy_W(35, 261) <= 0; flappy_W(35, 262) <= 0; flappy_W(35, 263) <= 0; flappy_W(35, 264) <= 0; flappy_W(35, 265) <= 0; flappy_W(35, 266) <= 0; flappy_W(35, 267) <= 0; flappy_W(35, 268) <= 0; flappy_W(35, 269) <= 0; flappy_W(35, 270) <= 0; flappy_W(35, 271) <= 0; flappy_W(35, 272) <= 0; flappy_W(35, 273) <= 0; flappy_W(35, 274) <= 0; flappy_W(35, 275) <= 0; flappy_W(35, 276) <= 0; flappy_W(35, 277) <= 0; flappy_W(35, 278) <= 0; flappy_W(35, 279) <= 0; flappy_W(35, 280) <= 0; flappy_W(35, 281) <= 0; flappy_W(35, 282) <= 0; flappy_W(35, 283) <= 0; flappy_W(35, 284) <= 0; flappy_W(35, 285) <= 0; flappy_W(35, 286) <= 0; flappy_W(35, 287) <= 0; flappy_W(35, 288) <= 1; flappy_W(35, 289) <= 1; flappy_W(35, 290) <= 1; flappy_W(35, 291) <= 1; flappy_W(35, 292) <= 1; flappy_W(35, 293) <= 1; flappy_W(35, 294) <= 1; flappy_W(35, 295) <= 1; flappy_W(35, 296) <= 1; flappy_W(35, 297) <= 1; flappy_W(35, 298) <= 1; flappy_W(35, 299) <= 1; flappy_W(35, 300) <= 0; flappy_W(35, 301) <= 0; flappy_W(35, 302) <= 0; flappy_W(35, 303) <= 0; flappy_W(35, 304) <= 0; flappy_W(35, 305) <= 0; flappy_W(35, 306) <= 0; flappy_W(35, 307) <= 0; flappy_W(35, 308) <= 0; flappy_W(35, 309) <= 0; flappy_W(35, 310) <= 0; flappy_W(35, 311) <= 0; flappy_W(35, 312) <= 0; flappy_W(35, 313) <= 0; flappy_W(35, 314) <= 0; flappy_W(35, 315) <= 0; flappy_W(35, 316) <= 0; flappy_W(35, 317) <= 0; flappy_W(35, 318) <= 0; flappy_W(35, 319) <= 0; flappy_W(35, 320) <= 0; flappy_W(35, 321) <= 0; flappy_W(35, 322) <= 0; flappy_W(35, 323) <= 0; flappy_W(35, 324) <= 0; flappy_W(35, 325) <= 0; flappy_W(35, 326) <= 0; flappy_W(35, 327) <= 0; flappy_W(35, 328) <= 0; flappy_W(35, 329) <= 0; flappy_W(35, 330) <= 0; flappy_W(35, 331) <= 0; flappy_W(35, 332) <= 0; flappy_W(35, 333) <= 0; flappy_W(35, 334) <= 0; flappy_W(35, 335) <= 0; flappy_W(35, 336) <= 0; flappy_W(35, 337) <= 0; flappy_W(35, 338) <= 0; flappy_W(35, 339) <= 0; flappy_W(35, 340) <= 0; flappy_W(35, 341) <= 0; flappy_W(35, 342) <= 0; flappy_W(35, 343) <= 0; flappy_W(35, 344) <= 0; flappy_W(35, 345) <= 0; flappy_W(35, 346) <= 0; flappy_W(35, 347) <= 0; flappy_W(35, 348) <= 0; flappy_W(35, 349) <= 0; flappy_W(35, 350) <= 0; flappy_W(35, 351) <= 0; flappy_W(35, 352) <= 0; flappy_W(35, 353) <= 0; flappy_W(35, 354) <= 0; flappy_W(35, 355) <= 0; flappy_W(35, 356) <= 0; flappy_W(35, 357) <= 0; flappy_W(35, 358) <= 0; flappy_W(35, 359) <= 0; flappy_W(35, 360) <= 0; flappy_W(35, 361) <= 0; flappy_W(35, 362) <= 0; flappy_W(35, 363) <= 0; flappy_W(35, 364) <= 0; flappy_W(35, 365) <= 0; flappy_W(35, 366) <= 0; flappy_W(35, 367) <= 0; flappy_W(35, 368) <= 0; flappy_W(35, 369) <= 0; flappy_W(35, 370) <= 0; flappy_W(35, 371) <= 0; flappy_W(35, 372) <= 0; flappy_W(35, 373) <= 0; flappy_W(35, 374) <= 0; flappy_W(35, 375) <= 0; flappy_W(35, 376) <= 0; flappy_W(35, 377) <= 0; flappy_W(35, 378) <= 0; flappy_W(35, 379) <= 0; flappy_W(35, 380) <= 0; flappy_W(35, 381) <= 0; flappy_W(35, 382) <= 0; flappy_W(35, 383) <= 0; flappy_W(35, 384) <= 0; flappy_W(35, 385) <= 0; flappy_W(35, 386) <= 0; flappy_W(35, 387) <= 0; flappy_W(35, 388) <= 0; flappy_W(35, 389) <= 0; flappy_W(35, 390) <= 0; flappy_W(35, 391) <= 0; flappy_W(35, 392) <= 0; flappy_W(35, 393) <= 0; flappy_W(35, 394) <= 0; flappy_W(35, 395) <= 0; flappy_W(35, 396) <= 0; flappy_W(35, 397) <= 0; flappy_W(35, 398) <= 0; flappy_W(35, 399) <= 0; flappy_W(35, 400) <= 0; flappy_W(35, 401) <= 0; flappy_W(35, 402) <= 1; flappy_W(35, 403) <= 1; flappy_W(35, 404) <= 1; flappy_W(35, 405) <= 1; flappy_W(35, 406) <= 1; flappy_W(35, 407) <= 1; flappy_W(35, 408) <= 1; flappy_W(35, 409) <= 1; flappy_W(35, 410) <= 1; flappy_W(35, 411) <= 1; flappy_W(35, 412) <= 1; flappy_W(35, 413) <= 1; flappy_W(35, 414) <= 0; flappy_W(35, 415) <= 0; flappy_W(35, 416) <= 0; flappy_W(35, 417) <= 0; flappy_W(35, 418) <= 0; flappy_W(35, 419) <= 0; flappy_W(35, 420) <= 0; flappy_W(35, 421) <= 0; flappy_W(35, 422) <= 0; flappy_W(35, 423) <= 0; flappy_W(35, 424) <= 0; flappy_W(35, 425) <= 0; flappy_W(35, 426) <= 1; flappy_W(35, 427) <= 1; flappy_W(35, 428) <= 1; flappy_W(35, 429) <= 1; flappy_W(35, 430) <= 1; flappy_W(35, 431) <= 1; flappy_W(35, 432) <= 1; flappy_W(35, 433) <= 1; flappy_W(35, 434) <= 1; flappy_W(35, 435) <= 1; flappy_W(35, 436) <= 1; flappy_W(35, 437) <= 1; flappy_W(35, 438) <= 0; flappy_W(35, 439) <= 0; flappy_W(35, 440) <= 0; flappy_W(35, 441) <= 0; flappy_W(35, 442) <= 0; flappy_W(35, 443) <= 0; flappy_W(35, 444) <= 0; flappy_W(35, 445) <= 0; flappy_W(35, 446) <= 0; flappy_W(35, 447) <= 0; flappy_W(35, 448) <= 0; flappy_W(35, 449) <= 0; flappy_W(35, 450) <= 0; flappy_W(35, 451) <= 0; flappy_W(35, 452) <= 0; flappy_W(35, 453) <= 0; flappy_W(35, 454) <= 0; flappy_W(35, 455) <= 0; flappy_W(35, 456) <= 0; flappy_W(35, 457) <= 0; flappy_W(35, 458) <= 0; flappy_W(35, 459) <= 0; flappy_W(35, 460) <= 0; flappy_W(35, 461) <= 0; flappy_W(35, 462) <= 0; flappy_W(35, 463) <= 0; flappy_W(35, 464) <= 0; flappy_W(35, 465) <= 0; flappy_W(35, 466) <= 0; flappy_W(35, 467) <= 0; flappy_W(35, 468) <= 1; flappy_W(35, 469) <= 1; flappy_W(35, 470) <= 1; flappy_W(35, 471) <= 1; flappy_W(35, 472) <= 1; flappy_W(35, 473) <= 1; flappy_W(35, 474) <= 1; flappy_W(35, 475) <= 1; flappy_W(35, 476) <= 1; flappy_W(35, 477) <= 1; flappy_W(35, 478) <= 1; flappy_W(35, 479) <= 1; flappy_W(35, 480) <= 0; flappy_W(35, 481) <= 0; flappy_W(35, 482) <= 0; flappy_W(35, 483) <= 0; flappy_W(35, 484) <= 0; flappy_W(35, 485) <= 0; flappy_W(35, 486) <= 0; flappy_W(35, 487) <= 0; flappy_W(35, 488) <= 0; flappy_W(35, 489) <= 0; flappy_W(35, 490) <= 0; flappy_W(35, 491) <= 0; flappy_W(35, 492) <= 0; flappy_W(35, 493) <= 0; flappy_W(35, 494) <= 0; flappy_W(35, 495) <= 0; flappy_W(35, 496) <= 0; flappy_W(35, 497) <= 0; flappy_W(35, 498) <= 0; flappy_W(35, 499) <= 0; flappy_W(35, 500) <= 0; flappy_W(35, 501) <= 0; flappy_W(35, 502) <= 0; flappy_W(35, 503) <= 0; flappy_W(35, 504) <= 0; flappy_W(35, 505) <= 0; flappy_W(35, 506) <= 0; flappy_W(35, 507) <= 0; flappy_W(35, 508) <= 0; flappy_W(35, 509) <= 0; flappy_W(35, 510) <= 1; flappy_W(35, 511) <= 1; flappy_W(35, 512) <= 1; flappy_W(35, 513) <= 1; flappy_W(35, 514) <= 1; flappy_W(35, 515) <= 1; flappy_W(35, 516) <= 1; flappy_W(35, 517) <= 1; flappy_W(35, 518) <= 1; flappy_W(35, 519) <= 1; flappy_W(35, 520) <= 1; flappy_W(35, 521) <= 1; flappy_W(35, 522) <= 0; flappy_W(35, 523) <= 0; flappy_W(35, 524) <= 0; flappy_W(35, 525) <= 0; flappy_W(35, 526) <= 0; flappy_W(35, 527) <= 0; flappy_W(35, 528) <= 1; flappy_W(35, 529) <= 1; flappy_W(35, 530) <= 1; flappy_W(35, 531) <= 1; flappy_W(35, 532) <= 1; flappy_W(35, 533) <= 1; flappy_W(35, 534) <= 1; flappy_W(35, 535) <= 1; flappy_W(35, 536) <= 1; flappy_W(35, 537) <= 1; flappy_W(35, 538) <= 1; flappy_W(35, 539) <= 1; flappy_W(35, 540) <= 0; flappy_W(35, 541) <= 0; flappy_W(35, 542) <= 0; flappy_W(35, 543) <= 0; flappy_W(35, 544) <= 0; flappy_W(35, 545) <= 0; flappy_W(35, 546) <= 0; flappy_W(35, 547) <= 0; flappy_W(35, 548) <= 0; flappy_W(35, 549) <= 0; flappy_W(35, 550) <= 0; flappy_W(35, 551) <= 0; flappy_W(35, 552) <= 0; flappy_W(35, 553) <= 0; flappy_W(35, 554) <= 0; flappy_W(35, 555) <= 0; flappy_W(35, 556) <= 0; flappy_W(35, 557) <= 0; flappy_W(35, 558) <= 0; flappy_W(35, 559) <= 0; flappy_W(35, 560) <= 0; flappy_W(35, 561) <= 0; flappy_W(35, 562) <= 0; flappy_W(35, 563) <= 0; flappy_W(35, 564) <= 1; flappy_W(35, 565) <= 1; flappy_W(35, 566) <= 1; flappy_W(35, 567) <= 1; flappy_W(35, 568) <= 1; flappy_W(35, 569) <= 1; flappy_W(35, 570) <= 1; flappy_W(35, 571) <= 1; flappy_W(35, 572) <= 1; flappy_W(35, 573) <= 1; flappy_W(35, 574) <= 1; flappy_W(35, 575) <= 1; flappy_W(35, 576) <= 0; flappy_W(35, 577) <= 0; flappy_W(35, 578) <= 0; flappy_W(35, 579) <= 0; flappy_W(35, 580) <= 0; flappy_W(35, 581) <= 0; flappy_W(35, 582) <= 0; flappy_W(35, 583) <= 0; flappy_W(35, 584) <= 0; flappy_W(35, 585) <= 0; flappy_W(35, 586) <= 0; flappy_W(35, 587) <= 0; flappy_W(35, 588) <= 1; flappy_W(35, 589) <= 1; flappy_W(35, 590) <= 1; flappy_W(35, 591) <= 1; flappy_W(35, 592) <= 1; flappy_W(35, 593) <= 1; 
flappy_W(36, 0) <= 0; flappy_W(36, 1) <= 0; flappy_W(36, 2) <= 0; flappy_W(36, 3) <= 0; flappy_W(36, 4) <= 0; flappy_W(36, 5) <= 0; flappy_W(36, 6) <= 1; flappy_W(36, 7) <= 1; flappy_W(36, 8) <= 1; flappy_W(36, 9) <= 1; flappy_W(36, 10) <= 1; flappy_W(36, 11) <= 1; flappy_W(36, 12) <= 1; flappy_W(36, 13) <= 1; flappy_W(36, 14) <= 1; flappy_W(36, 15) <= 1; flappy_W(36, 16) <= 1; flappy_W(36, 17) <= 1; flappy_W(36, 18) <= 0; flappy_W(36, 19) <= 0; flappy_W(36, 20) <= 0; flappy_W(36, 21) <= 0; flappy_W(36, 22) <= 0; flappy_W(36, 23) <= 0; flappy_W(36, 24) <= 0; flappy_W(36, 25) <= 0; flappy_W(36, 26) <= 0; flappy_W(36, 27) <= 0; flappy_W(36, 28) <= 0; flappy_W(36, 29) <= 0; flappy_W(36, 30) <= 0; flappy_W(36, 31) <= 0; flappy_W(36, 32) <= 0; flappy_W(36, 33) <= 0; flappy_W(36, 34) <= 0; flappy_W(36, 35) <= 0; flappy_W(36, 36) <= 0; flappy_W(36, 37) <= 0; flappy_W(36, 38) <= 0; flappy_W(36, 39) <= 0; flappy_W(36, 40) <= 0; flappy_W(36, 41) <= 0; flappy_W(36, 42) <= 0; flappy_W(36, 43) <= 0; flappy_W(36, 44) <= 0; flappy_W(36, 45) <= 0; flappy_W(36, 46) <= 0; flappy_W(36, 47) <= 0; flappy_W(36, 48) <= 0; flappy_W(36, 49) <= 0; flappy_W(36, 50) <= 0; flappy_W(36, 51) <= 0; flappy_W(36, 52) <= 0; flappy_W(36, 53) <= 0; flappy_W(36, 54) <= 0; flappy_W(36, 55) <= 0; flappy_W(36, 56) <= 0; flappy_W(36, 57) <= 0; flappy_W(36, 58) <= 0; flappy_W(36, 59) <= 0; flappy_W(36, 60) <= 1; flappy_W(36, 61) <= 1; flappy_W(36, 62) <= 1; flappy_W(36, 63) <= 1; flappy_W(36, 64) <= 1; flappy_W(36, 65) <= 1; flappy_W(36, 66) <= 1; flappy_W(36, 67) <= 1; flappy_W(36, 68) <= 1; flappy_W(36, 69) <= 1; flappy_W(36, 70) <= 1; flappy_W(36, 71) <= 1; flappy_W(36, 72) <= 0; flappy_W(36, 73) <= 0; flappy_W(36, 74) <= 0; flappy_W(36, 75) <= 0; flappy_W(36, 76) <= 0; flappy_W(36, 77) <= 0; flappy_W(36, 78) <= 0; flappy_W(36, 79) <= 0; flappy_W(36, 80) <= 0; flappy_W(36, 81) <= 0; flappy_W(36, 82) <= 0; flappy_W(36, 83) <= 0; flappy_W(36, 84) <= 0; flappy_W(36, 85) <= 0; flappy_W(36, 86) <= 0; flappy_W(36, 87) <= 0; flappy_W(36, 88) <= 0; flappy_W(36, 89) <= 0; flappy_W(36, 90) <= 0; flappy_W(36, 91) <= 0; flappy_W(36, 92) <= 0; flappy_W(36, 93) <= 0; flappy_W(36, 94) <= 0; flappy_W(36, 95) <= 0; flappy_W(36, 96) <= 0; flappy_W(36, 97) <= 0; flappy_W(36, 98) <= 0; flappy_W(36, 99) <= 0; flappy_W(36, 100) <= 0; flappy_W(36, 101) <= 0; flappy_W(36, 102) <= 0; flappy_W(36, 103) <= 0; flappy_W(36, 104) <= 0; flappy_W(36, 105) <= 0; flappy_W(36, 106) <= 0; flappy_W(36, 107) <= 0; flappy_W(36, 108) <= 1; flappy_W(36, 109) <= 1; flappy_W(36, 110) <= 1; flappy_W(36, 111) <= 1; flappy_W(36, 112) <= 1; flappy_W(36, 113) <= 1; flappy_W(36, 114) <= 1; flappy_W(36, 115) <= 1; flappy_W(36, 116) <= 1; flappy_W(36, 117) <= 1; flappy_W(36, 118) <= 1; flappy_W(36, 119) <= 1; flappy_W(36, 120) <= 0; flappy_W(36, 121) <= 0; flappy_W(36, 122) <= 0; flappy_W(36, 123) <= 0; flappy_W(36, 124) <= 0; flappy_W(36, 125) <= 0; flappy_W(36, 126) <= 0; flappy_W(36, 127) <= 0; flappy_W(36, 128) <= 0; flappy_W(36, 129) <= 0; flappy_W(36, 130) <= 0; flappy_W(36, 131) <= 0; flappy_W(36, 132) <= 0; flappy_W(36, 133) <= 0; flappy_W(36, 134) <= 0; flappy_W(36, 135) <= 0; flappy_W(36, 136) <= 0; flappy_W(36, 137) <= 0; flappy_W(36, 138) <= 1; flappy_W(36, 139) <= 1; flappy_W(36, 140) <= 1; flappy_W(36, 141) <= 1; flappy_W(36, 142) <= 1; flappy_W(36, 143) <= 1; flappy_W(36, 144) <= 1; flappy_W(36, 145) <= 1; flappy_W(36, 146) <= 1; flappy_W(36, 147) <= 1; flappy_W(36, 148) <= 1; flappy_W(36, 149) <= 1; flappy_W(36, 150) <= 0; flappy_W(36, 151) <= 0; flappy_W(36, 152) <= 0; flappy_W(36, 153) <= 0; flappy_W(36, 154) <= 0; flappy_W(36, 155) <= 0; flappy_W(36, 156) <= 0; flappy_W(36, 157) <= 0; flappy_W(36, 158) <= 0; flappy_W(36, 159) <= 0; flappy_W(36, 160) <= 0; flappy_W(36, 161) <= 0; flappy_W(36, 162) <= 0; flappy_W(36, 163) <= 0; flappy_W(36, 164) <= 0; flappy_W(36, 165) <= 0; flappy_W(36, 166) <= 0; flappy_W(36, 167) <= 0; flappy_W(36, 168) <= 1; flappy_W(36, 169) <= 1; flappy_W(36, 170) <= 1; flappy_W(36, 171) <= 1; flappy_W(36, 172) <= 1; flappy_W(36, 173) <= 1; flappy_W(36, 174) <= 1; flappy_W(36, 175) <= 1; flappy_W(36, 176) <= 1; flappy_W(36, 177) <= 1; flappy_W(36, 178) <= 1; flappy_W(36, 179) <= 1; flappy_W(36, 180) <= 0; flappy_W(36, 181) <= 0; flappy_W(36, 182) <= 0; flappy_W(36, 183) <= 0; flappy_W(36, 184) <= 0; flappy_W(36, 185) <= 0; flappy_W(36, 186) <= 0; flappy_W(36, 187) <= 0; flappy_W(36, 188) <= 0; flappy_W(36, 189) <= 0; flappy_W(36, 190) <= 0; flappy_W(36, 191) <= 0; flappy_W(36, 192) <= 0; flappy_W(36, 193) <= 0; flappy_W(36, 194) <= 0; flappy_W(36, 195) <= 0; flappy_W(36, 196) <= 0; flappy_W(36, 197) <= 0; flappy_W(36, 198) <= 0; flappy_W(36, 199) <= 0; flappy_W(36, 200) <= 0; flappy_W(36, 201) <= 0; flappy_W(36, 202) <= 0; flappy_W(36, 203) <= 0; flappy_W(36, 204) <= 0; flappy_W(36, 205) <= 0; flappy_W(36, 206) <= 0; flappy_W(36, 207) <= 0; flappy_W(36, 208) <= 0; flappy_W(36, 209) <= 0; flappy_W(36, 210) <= 0; flappy_W(36, 211) <= 0; flappy_W(36, 212) <= 0; flappy_W(36, 213) <= 0; flappy_W(36, 214) <= 0; flappy_W(36, 215) <= 0; flappy_W(36, 216) <= 0; flappy_W(36, 217) <= 0; flappy_W(36, 218) <= 0; flappy_W(36, 219) <= 0; flappy_W(36, 220) <= 0; flappy_W(36, 221) <= 0; flappy_W(36, 222) <= 1; flappy_W(36, 223) <= 1; flappy_W(36, 224) <= 1; flappy_W(36, 225) <= 1; flappy_W(36, 226) <= 1; flappy_W(36, 227) <= 1; flappy_W(36, 228) <= 1; flappy_W(36, 229) <= 1; flappy_W(36, 230) <= 1; flappy_W(36, 231) <= 1; flappy_W(36, 232) <= 1; flappy_W(36, 233) <= 1; flappy_W(36, 234) <= 0; flappy_W(36, 235) <= 0; flappy_W(36, 236) <= 0; flappy_W(36, 237) <= 0; flappy_W(36, 238) <= 0; flappy_W(36, 239) <= 0; flappy_W(36, 240) <= 0; flappy_W(36, 241) <= 0; flappy_W(36, 242) <= 0; flappy_W(36, 243) <= 0; flappy_W(36, 244) <= 0; flappy_W(36, 245) <= 0; flappy_W(36, 246) <= 0; flappy_W(36, 247) <= 0; flappy_W(36, 248) <= 0; flappy_W(36, 249) <= 0; flappy_W(36, 250) <= 0; flappy_W(36, 251) <= 0; flappy_W(36, 252) <= 0; flappy_W(36, 253) <= 0; flappy_W(36, 254) <= 0; flappy_W(36, 255) <= 0; flappy_W(36, 256) <= 0; flappy_W(36, 257) <= 0; flappy_W(36, 258) <= 0; flappy_W(36, 259) <= 0; flappy_W(36, 260) <= 0; flappy_W(36, 261) <= 0; flappy_W(36, 262) <= 0; flappy_W(36, 263) <= 0; flappy_W(36, 264) <= 0; flappy_W(36, 265) <= 0; flappy_W(36, 266) <= 0; flappy_W(36, 267) <= 0; flappy_W(36, 268) <= 0; flappy_W(36, 269) <= 0; flappy_W(36, 270) <= 0; flappy_W(36, 271) <= 0; flappy_W(36, 272) <= 0; flappy_W(36, 273) <= 0; flappy_W(36, 274) <= 0; flappy_W(36, 275) <= 0; flappy_W(36, 276) <= 0; flappy_W(36, 277) <= 0; flappy_W(36, 278) <= 0; flappy_W(36, 279) <= 0; flappy_W(36, 280) <= 0; flappy_W(36, 281) <= 0; flappy_W(36, 282) <= 0; flappy_W(36, 283) <= 0; flappy_W(36, 284) <= 0; flappy_W(36, 285) <= 0; flappy_W(36, 286) <= 0; flappy_W(36, 287) <= 0; flappy_W(36, 288) <= 1; flappy_W(36, 289) <= 1; flappy_W(36, 290) <= 1; flappy_W(36, 291) <= 1; flappy_W(36, 292) <= 1; flappy_W(36, 293) <= 1; flappy_W(36, 294) <= 1; flappy_W(36, 295) <= 1; flappy_W(36, 296) <= 1; flappy_W(36, 297) <= 1; flappy_W(36, 298) <= 1; flappy_W(36, 299) <= 1; flappy_W(36, 300) <= 0; flappy_W(36, 301) <= 0; flappy_W(36, 302) <= 0; flappy_W(36, 303) <= 0; flappy_W(36, 304) <= 0; flappy_W(36, 305) <= 0; flappy_W(36, 306) <= 0; flappy_W(36, 307) <= 0; flappy_W(36, 308) <= 0; flappy_W(36, 309) <= 0; flappy_W(36, 310) <= 0; flappy_W(36, 311) <= 0; flappy_W(36, 312) <= 0; flappy_W(36, 313) <= 0; flappy_W(36, 314) <= 0; flappy_W(36, 315) <= 0; flappy_W(36, 316) <= 0; flappy_W(36, 317) <= 0; flappy_W(36, 318) <= 0; flappy_W(36, 319) <= 0; flappy_W(36, 320) <= 0; flappy_W(36, 321) <= 0; flappy_W(36, 322) <= 0; flappy_W(36, 323) <= 0; flappy_W(36, 324) <= 0; flappy_W(36, 325) <= 0; flappy_W(36, 326) <= 0; flappy_W(36, 327) <= 0; flappy_W(36, 328) <= 0; flappy_W(36, 329) <= 0; flappy_W(36, 330) <= 0; flappy_W(36, 331) <= 0; flappy_W(36, 332) <= 0; flappy_W(36, 333) <= 0; flappy_W(36, 334) <= 0; flappy_W(36, 335) <= 0; flappy_W(36, 336) <= 0; flappy_W(36, 337) <= 0; flappy_W(36, 338) <= 0; flappy_W(36, 339) <= 0; flappy_W(36, 340) <= 0; flappy_W(36, 341) <= 0; flappy_W(36, 342) <= 0; flappy_W(36, 343) <= 0; flappy_W(36, 344) <= 0; flappy_W(36, 345) <= 0; flappy_W(36, 346) <= 0; flappy_W(36, 347) <= 0; flappy_W(36, 348) <= 0; flappy_W(36, 349) <= 0; flappy_W(36, 350) <= 0; flappy_W(36, 351) <= 0; flappy_W(36, 352) <= 0; flappy_W(36, 353) <= 0; flappy_W(36, 354) <= 0; flappy_W(36, 355) <= 0; flappy_W(36, 356) <= 0; flappy_W(36, 357) <= 0; flappy_W(36, 358) <= 0; flappy_W(36, 359) <= 0; flappy_W(36, 360) <= 0; flappy_W(36, 361) <= 0; flappy_W(36, 362) <= 0; flappy_W(36, 363) <= 0; flappy_W(36, 364) <= 0; flappy_W(36, 365) <= 0; flappy_W(36, 366) <= 0; flappy_W(36, 367) <= 0; flappy_W(36, 368) <= 0; flappy_W(36, 369) <= 0; flappy_W(36, 370) <= 0; flappy_W(36, 371) <= 0; flappy_W(36, 372) <= 0; flappy_W(36, 373) <= 0; flappy_W(36, 374) <= 0; flappy_W(36, 375) <= 0; flappy_W(36, 376) <= 0; flappy_W(36, 377) <= 0; flappy_W(36, 378) <= 0; flappy_W(36, 379) <= 0; flappy_W(36, 380) <= 0; flappy_W(36, 381) <= 0; flappy_W(36, 382) <= 0; flappy_W(36, 383) <= 0; flappy_W(36, 384) <= 0; flappy_W(36, 385) <= 0; flappy_W(36, 386) <= 0; flappy_W(36, 387) <= 0; flappy_W(36, 388) <= 0; flappy_W(36, 389) <= 0; flappy_W(36, 390) <= 0; flappy_W(36, 391) <= 0; flappy_W(36, 392) <= 0; flappy_W(36, 393) <= 0; flappy_W(36, 394) <= 0; flappy_W(36, 395) <= 0; flappy_W(36, 396) <= 0; flappy_W(36, 397) <= 0; flappy_W(36, 398) <= 0; flappy_W(36, 399) <= 0; flappy_W(36, 400) <= 0; flappy_W(36, 401) <= 0; flappy_W(36, 402) <= 1; flappy_W(36, 403) <= 1; flappy_W(36, 404) <= 1; flappy_W(36, 405) <= 1; flappy_W(36, 406) <= 1; flappy_W(36, 407) <= 1; flappy_W(36, 408) <= 1; flappy_W(36, 409) <= 1; flappy_W(36, 410) <= 1; flappy_W(36, 411) <= 1; flappy_W(36, 412) <= 1; flappy_W(36, 413) <= 1; flappy_W(36, 414) <= 0; flappy_W(36, 415) <= 0; flappy_W(36, 416) <= 0; flappy_W(36, 417) <= 0; flappy_W(36, 418) <= 0; flappy_W(36, 419) <= 0; flappy_W(36, 420) <= 0; flappy_W(36, 421) <= 0; flappy_W(36, 422) <= 0; flappy_W(36, 423) <= 0; flappy_W(36, 424) <= 0; flappy_W(36, 425) <= 0; flappy_W(36, 426) <= 1; flappy_W(36, 427) <= 1; flappy_W(36, 428) <= 1; flappy_W(36, 429) <= 1; flappy_W(36, 430) <= 1; flappy_W(36, 431) <= 1; flappy_W(36, 432) <= 1; flappy_W(36, 433) <= 1; flappy_W(36, 434) <= 1; flappy_W(36, 435) <= 1; flappy_W(36, 436) <= 1; flappy_W(36, 437) <= 1; flappy_W(36, 438) <= 0; flappy_W(36, 439) <= 0; flappy_W(36, 440) <= 0; flappy_W(36, 441) <= 0; flappy_W(36, 442) <= 0; flappy_W(36, 443) <= 0; flappy_W(36, 444) <= 0; flappy_W(36, 445) <= 0; flappy_W(36, 446) <= 0; flappy_W(36, 447) <= 0; flappy_W(36, 448) <= 0; flappy_W(36, 449) <= 0; flappy_W(36, 450) <= 0; flappy_W(36, 451) <= 0; flappy_W(36, 452) <= 0; flappy_W(36, 453) <= 0; flappy_W(36, 454) <= 0; flappy_W(36, 455) <= 0; flappy_W(36, 456) <= 0; flappy_W(36, 457) <= 0; flappy_W(36, 458) <= 0; flappy_W(36, 459) <= 0; flappy_W(36, 460) <= 0; flappy_W(36, 461) <= 0; flappy_W(36, 462) <= 0; flappy_W(36, 463) <= 0; flappy_W(36, 464) <= 0; flappy_W(36, 465) <= 0; flappy_W(36, 466) <= 0; flappy_W(36, 467) <= 0; flappy_W(36, 468) <= 1; flappy_W(36, 469) <= 1; flappy_W(36, 470) <= 1; flappy_W(36, 471) <= 1; flappy_W(36, 472) <= 1; flappy_W(36, 473) <= 1; flappy_W(36, 474) <= 1; flappy_W(36, 475) <= 1; flappy_W(36, 476) <= 1; flappy_W(36, 477) <= 1; flappy_W(36, 478) <= 1; flappy_W(36, 479) <= 1; flappy_W(36, 480) <= 0; flappy_W(36, 481) <= 0; flappy_W(36, 482) <= 0; flappy_W(36, 483) <= 0; flappy_W(36, 484) <= 0; flappy_W(36, 485) <= 0; flappy_W(36, 486) <= 0; flappy_W(36, 487) <= 0; flappy_W(36, 488) <= 0; flappy_W(36, 489) <= 0; flappy_W(36, 490) <= 0; flappy_W(36, 491) <= 0; flappy_W(36, 492) <= 0; flappy_W(36, 493) <= 0; flappy_W(36, 494) <= 0; flappy_W(36, 495) <= 0; flappy_W(36, 496) <= 0; flappy_W(36, 497) <= 0; flappy_W(36, 498) <= 0; flappy_W(36, 499) <= 0; flappy_W(36, 500) <= 0; flappy_W(36, 501) <= 0; flappy_W(36, 502) <= 0; flappy_W(36, 503) <= 0; flappy_W(36, 504) <= 0; flappy_W(36, 505) <= 0; flappy_W(36, 506) <= 0; flappy_W(36, 507) <= 0; flappy_W(36, 508) <= 0; flappy_W(36, 509) <= 0; flappy_W(36, 510) <= 1; flappy_W(36, 511) <= 1; flappy_W(36, 512) <= 1; flappy_W(36, 513) <= 1; flappy_W(36, 514) <= 1; flappy_W(36, 515) <= 1; flappy_W(36, 516) <= 1; flappy_W(36, 517) <= 1; flappy_W(36, 518) <= 1; flappy_W(36, 519) <= 1; flappy_W(36, 520) <= 1; flappy_W(36, 521) <= 1; flappy_W(36, 522) <= 0; flappy_W(36, 523) <= 0; flappy_W(36, 524) <= 0; flappy_W(36, 525) <= 0; flappy_W(36, 526) <= 0; flappy_W(36, 527) <= 0; flappy_W(36, 528) <= 0; flappy_W(36, 529) <= 0; flappy_W(36, 530) <= 0; flappy_W(36, 531) <= 0; flappy_W(36, 532) <= 0; flappy_W(36, 533) <= 0; flappy_W(36, 534) <= 1; flappy_W(36, 535) <= 1; flappy_W(36, 536) <= 1; flappy_W(36, 537) <= 1; flappy_W(36, 538) <= 1; flappy_W(36, 539) <= 1; flappy_W(36, 540) <= 1; flappy_W(36, 541) <= 1; flappy_W(36, 542) <= 1; flappy_W(36, 543) <= 1; flappy_W(36, 544) <= 1; flappy_W(36, 545) <= 1; flappy_W(36, 546) <= 0; flappy_W(36, 547) <= 0; flappy_W(36, 548) <= 0; flappy_W(36, 549) <= 0; flappy_W(36, 550) <= 0; flappy_W(36, 551) <= 0; flappy_W(36, 552) <= 0; flappy_W(36, 553) <= 0; flappy_W(36, 554) <= 0; flappy_W(36, 555) <= 0; flappy_W(36, 556) <= 0; flappy_W(36, 557) <= 0; flappy_W(36, 558) <= 0; flappy_W(36, 559) <= 0; flappy_W(36, 560) <= 0; flappy_W(36, 561) <= 0; flappy_W(36, 562) <= 0; flappy_W(36, 563) <= 0; flappy_W(36, 564) <= 1; flappy_W(36, 565) <= 1; flappy_W(36, 566) <= 1; flappy_W(36, 567) <= 1; flappy_W(36, 568) <= 1; flappy_W(36, 569) <= 1; flappy_W(36, 570) <= 1; flappy_W(36, 571) <= 1; flappy_W(36, 572) <= 1; flappy_W(36, 573) <= 1; flappy_W(36, 574) <= 1; flappy_W(36, 575) <= 1; flappy_W(36, 576) <= 0; flappy_W(36, 577) <= 0; flappy_W(36, 578) <= 0; flappy_W(36, 579) <= 0; flappy_W(36, 580) <= 0; flappy_W(36, 581) <= 0; flappy_W(36, 582) <= 0; flappy_W(36, 583) <= 0; flappy_W(36, 584) <= 0; flappy_W(36, 585) <= 0; flappy_W(36, 586) <= 0; flappy_W(36, 587) <= 0; flappy_W(36, 588) <= 1; flappy_W(36, 589) <= 1; flappy_W(36, 590) <= 1; flappy_W(36, 591) <= 1; flappy_W(36, 592) <= 1; flappy_W(36, 593) <= 1; 
flappy_W(37, 0) <= 0; flappy_W(37, 1) <= 0; flappy_W(37, 2) <= 0; flappy_W(37, 3) <= 0; flappy_W(37, 4) <= 0; flappy_W(37, 5) <= 0; flappy_W(37, 6) <= 1; flappy_W(37, 7) <= 1; flappy_W(37, 8) <= 1; flappy_W(37, 9) <= 1; flappy_W(37, 10) <= 1; flappy_W(37, 11) <= 1; flappy_W(37, 12) <= 1; flappy_W(37, 13) <= 1; flappy_W(37, 14) <= 1; flappy_W(37, 15) <= 1; flappy_W(37, 16) <= 1; flappy_W(37, 17) <= 1; flappy_W(37, 18) <= 0; flappy_W(37, 19) <= 0; flappy_W(37, 20) <= 0; flappy_W(37, 21) <= 0; flappy_W(37, 22) <= 0; flappy_W(37, 23) <= 0; flappy_W(37, 24) <= 0; flappy_W(37, 25) <= 0; flappy_W(37, 26) <= 0; flappy_W(37, 27) <= 0; flappy_W(37, 28) <= 0; flappy_W(37, 29) <= 0; flappy_W(37, 30) <= 0; flappy_W(37, 31) <= 0; flappy_W(37, 32) <= 0; flappy_W(37, 33) <= 0; flappy_W(37, 34) <= 0; flappy_W(37, 35) <= 0; flappy_W(37, 36) <= 0; flappy_W(37, 37) <= 0; flappy_W(37, 38) <= 0; flappy_W(37, 39) <= 0; flappy_W(37, 40) <= 0; flappy_W(37, 41) <= 0; flappy_W(37, 42) <= 0; flappy_W(37, 43) <= 0; flappy_W(37, 44) <= 0; flappy_W(37, 45) <= 0; flappy_W(37, 46) <= 0; flappy_W(37, 47) <= 0; flappy_W(37, 48) <= 0; flappy_W(37, 49) <= 0; flappy_W(37, 50) <= 0; flappy_W(37, 51) <= 0; flappy_W(37, 52) <= 0; flappy_W(37, 53) <= 0; flappy_W(37, 54) <= 0; flappy_W(37, 55) <= 0; flappy_W(37, 56) <= 0; flappy_W(37, 57) <= 0; flappy_W(37, 58) <= 0; flappy_W(37, 59) <= 0; flappy_W(37, 60) <= 1; flappy_W(37, 61) <= 1; flappy_W(37, 62) <= 1; flappy_W(37, 63) <= 1; flappy_W(37, 64) <= 1; flappy_W(37, 65) <= 1; flappy_W(37, 66) <= 1; flappy_W(37, 67) <= 1; flappy_W(37, 68) <= 1; flappy_W(37, 69) <= 1; flappy_W(37, 70) <= 1; flappy_W(37, 71) <= 1; flappy_W(37, 72) <= 0; flappy_W(37, 73) <= 0; flappy_W(37, 74) <= 0; flappy_W(37, 75) <= 0; flappy_W(37, 76) <= 0; flappy_W(37, 77) <= 0; flappy_W(37, 78) <= 0; flappy_W(37, 79) <= 0; flappy_W(37, 80) <= 0; flappy_W(37, 81) <= 0; flappy_W(37, 82) <= 0; flappy_W(37, 83) <= 0; flappy_W(37, 84) <= 0; flappy_W(37, 85) <= 0; flappy_W(37, 86) <= 0; flappy_W(37, 87) <= 0; flappy_W(37, 88) <= 0; flappy_W(37, 89) <= 0; flappy_W(37, 90) <= 0; flappy_W(37, 91) <= 0; flappy_W(37, 92) <= 0; flappy_W(37, 93) <= 0; flappy_W(37, 94) <= 0; flappy_W(37, 95) <= 0; flappy_W(37, 96) <= 0; flappy_W(37, 97) <= 0; flappy_W(37, 98) <= 0; flappy_W(37, 99) <= 0; flappy_W(37, 100) <= 0; flappy_W(37, 101) <= 0; flappy_W(37, 102) <= 0; flappy_W(37, 103) <= 0; flappy_W(37, 104) <= 0; flappy_W(37, 105) <= 0; flappy_W(37, 106) <= 0; flappy_W(37, 107) <= 0; flappy_W(37, 108) <= 1; flappy_W(37, 109) <= 1; flappy_W(37, 110) <= 1; flappy_W(37, 111) <= 1; flappy_W(37, 112) <= 1; flappy_W(37, 113) <= 1; flappy_W(37, 114) <= 1; flappy_W(37, 115) <= 1; flappy_W(37, 116) <= 1; flappy_W(37, 117) <= 1; flappy_W(37, 118) <= 1; flappy_W(37, 119) <= 1; flappy_W(37, 120) <= 0; flappy_W(37, 121) <= 0; flappy_W(37, 122) <= 0; flappy_W(37, 123) <= 0; flappy_W(37, 124) <= 0; flappy_W(37, 125) <= 0; flappy_W(37, 126) <= 0; flappy_W(37, 127) <= 0; flappy_W(37, 128) <= 0; flappy_W(37, 129) <= 0; flappy_W(37, 130) <= 0; flappy_W(37, 131) <= 0; flappy_W(37, 132) <= 0; flappy_W(37, 133) <= 0; flappy_W(37, 134) <= 0; flappy_W(37, 135) <= 0; flappy_W(37, 136) <= 0; flappy_W(37, 137) <= 0; flappy_W(37, 138) <= 1; flappy_W(37, 139) <= 1; flappy_W(37, 140) <= 1; flappy_W(37, 141) <= 1; flappy_W(37, 142) <= 1; flappy_W(37, 143) <= 1; flappy_W(37, 144) <= 1; flappy_W(37, 145) <= 1; flappy_W(37, 146) <= 1; flappy_W(37, 147) <= 1; flappy_W(37, 148) <= 1; flappy_W(37, 149) <= 1; flappy_W(37, 150) <= 0; flappy_W(37, 151) <= 0; flappy_W(37, 152) <= 0; flappy_W(37, 153) <= 0; flappy_W(37, 154) <= 0; flappy_W(37, 155) <= 0; flappy_W(37, 156) <= 0; flappy_W(37, 157) <= 0; flappy_W(37, 158) <= 0; flappy_W(37, 159) <= 0; flappy_W(37, 160) <= 0; flappy_W(37, 161) <= 0; flappy_W(37, 162) <= 0; flappy_W(37, 163) <= 0; flappy_W(37, 164) <= 0; flappy_W(37, 165) <= 0; flappy_W(37, 166) <= 0; flappy_W(37, 167) <= 0; flappy_W(37, 168) <= 1; flappy_W(37, 169) <= 1; flappy_W(37, 170) <= 1; flappy_W(37, 171) <= 1; flappy_W(37, 172) <= 1; flappy_W(37, 173) <= 1; flappy_W(37, 174) <= 1; flappy_W(37, 175) <= 1; flappy_W(37, 176) <= 1; flappy_W(37, 177) <= 1; flappy_W(37, 178) <= 1; flappy_W(37, 179) <= 1; flappy_W(37, 180) <= 0; flappy_W(37, 181) <= 0; flappy_W(37, 182) <= 0; flappy_W(37, 183) <= 0; flappy_W(37, 184) <= 0; flappy_W(37, 185) <= 0; flappy_W(37, 186) <= 0; flappy_W(37, 187) <= 0; flappy_W(37, 188) <= 0; flappy_W(37, 189) <= 0; flappy_W(37, 190) <= 0; flappy_W(37, 191) <= 0; flappy_W(37, 192) <= 0; flappy_W(37, 193) <= 0; flappy_W(37, 194) <= 0; flappy_W(37, 195) <= 0; flappy_W(37, 196) <= 0; flappy_W(37, 197) <= 0; flappy_W(37, 198) <= 0; flappy_W(37, 199) <= 0; flappy_W(37, 200) <= 0; flappy_W(37, 201) <= 0; flappy_W(37, 202) <= 0; flappy_W(37, 203) <= 0; flappy_W(37, 204) <= 0; flappy_W(37, 205) <= 0; flappy_W(37, 206) <= 0; flappy_W(37, 207) <= 0; flappy_W(37, 208) <= 0; flappy_W(37, 209) <= 0; flappy_W(37, 210) <= 0; flappy_W(37, 211) <= 0; flappy_W(37, 212) <= 0; flappy_W(37, 213) <= 0; flappy_W(37, 214) <= 0; flappy_W(37, 215) <= 0; flappy_W(37, 216) <= 0; flappy_W(37, 217) <= 0; flappy_W(37, 218) <= 0; flappy_W(37, 219) <= 0; flappy_W(37, 220) <= 0; flappy_W(37, 221) <= 0; flappy_W(37, 222) <= 1; flappy_W(37, 223) <= 1; flappy_W(37, 224) <= 1; flappy_W(37, 225) <= 1; flappy_W(37, 226) <= 1; flappy_W(37, 227) <= 1; flappy_W(37, 228) <= 1; flappy_W(37, 229) <= 1; flappy_W(37, 230) <= 1; flappy_W(37, 231) <= 1; flappy_W(37, 232) <= 1; flappy_W(37, 233) <= 1; flappy_W(37, 234) <= 0; flappy_W(37, 235) <= 0; flappy_W(37, 236) <= 0; flappy_W(37, 237) <= 0; flappy_W(37, 238) <= 0; flappy_W(37, 239) <= 0; flappy_W(37, 240) <= 0; flappy_W(37, 241) <= 0; flappy_W(37, 242) <= 0; flappy_W(37, 243) <= 0; flappy_W(37, 244) <= 0; flappy_W(37, 245) <= 0; flappy_W(37, 246) <= 0; flappy_W(37, 247) <= 0; flappy_W(37, 248) <= 0; flappy_W(37, 249) <= 0; flappy_W(37, 250) <= 0; flappy_W(37, 251) <= 0; flappy_W(37, 252) <= 0; flappy_W(37, 253) <= 0; flappy_W(37, 254) <= 0; flappy_W(37, 255) <= 0; flappy_W(37, 256) <= 0; flappy_W(37, 257) <= 0; flappy_W(37, 258) <= 0; flappy_W(37, 259) <= 0; flappy_W(37, 260) <= 0; flappy_W(37, 261) <= 0; flappy_W(37, 262) <= 0; flappy_W(37, 263) <= 0; flappy_W(37, 264) <= 0; flappy_W(37, 265) <= 0; flappy_W(37, 266) <= 0; flappy_W(37, 267) <= 0; flappy_W(37, 268) <= 0; flappy_W(37, 269) <= 0; flappy_W(37, 270) <= 0; flappy_W(37, 271) <= 0; flappy_W(37, 272) <= 0; flappy_W(37, 273) <= 0; flappy_W(37, 274) <= 0; flappy_W(37, 275) <= 0; flappy_W(37, 276) <= 0; flappy_W(37, 277) <= 0; flappy_W(37, 278) <= 0; flappy_W(37, 279) <= 0; flappy_W(37, 280) <= 0; flappy_W(37, 281) <= 0; flappy_W(37, 282) <= 0; flappy_W(37, 283) <= 0; flappy_W(37, 284) <= 0; flappy_W(37, 285) <= 0; flappy_W(37, 286) <= 0; flappy_W(37, 287) <= 0; flappy_W(37, 288) <= 1; flappy_W(37, 289) <= 1; flappy_W(37, 290) <= 1; flappy_W(37, 291) <= 1; flappy_W(37, 292) <= 1; flappy_W(37, 293) <= 1; flappy_W(37, 294) <= 1; flappy_W(37, 295) <= 1; flappy_W(37, 296) <= 1; flappy_W(37, 297) <= 1; flappy_W(37, 298) <= 1; flappy_W(37, 299) <= 1; flappy_W(37, 300) <= 0; flappy_W(37, 301) <= 0; flappy_W(37, 302) <= 0; flappy_W(37, 303) <= 0; flappy_W(37, 304) <= 0; flappy_W(37, 305) <= 0; flappy_W(37, 306) <= 0; flappy_W(37, 307) <= 0; flappy_W(37, 308) <= 0; flappy_W(37, 309) <= 0; flappy_W(37, 310) <= 0; flappy_W(37, 311) <= 0; flappy_W(37, 312) <= 0; flappy_W(37, 313) <= 0; flappy_W(37, 314) <= 0; flappy_W(37, 315) <= 0; flappy_W(37, 316) <= 0; flappy_W(37, 317) <= 0; flappy_W(37, 318) <= 0; flappy_W(37, 319) <= 0; flappy_W(37, 320) <= 0; flappy_W(37, 321) <= 0; flappy_W(37, 322) <= 0; flappy_W(37, 323) <= 0; flappy_W(37, 324) <= 0; flappy_W(37, 325) <= 0; flappy_W(37, 326) <= 0; flappy_W(37, 327) <= 0; flappy_W(37, 328) <= 0; flappy_W(37, 329) <= 0; flappy_W(37, 330) <= 0; flappy_W(37, 331) <= 0; flappy_W(37, 332) <= 0; flappy_W(37, 333) <= 0; flappy_W(37, 334) <= 0; flappy_W(37, 335) <= 0; flappy_W(37, 336) <= 0; flappy_W(37, 337) <= 0; flappy_W(37, 338) <= 0; flappy_W(37, 339) <= 0; flappy_W(37, 340) <= 0; flappy_W(37, 341) <= 0; flappy_W(37, 342) <= 0; flappy_W(37, 343) <= 0; flappy_W(37, 344) <= 0; flappy_W(37, 345) <= 0; flappy_W(37, 346) <= 0; flappy_W(37, 347) <= 0; flappy_W(37, 348) <= 0; flappy_W(37, 349) <= 0; flappy_W(37, 350) <= 0; flappy_W(37, 351) <= 0; flappy_W(37, 352) <= 0; flappy_W(37, 353) <= 0; flappy_W(37, 354) <= 0; flappy_W(37, 355) <= 0; flappy_W(37, 356) <= 0; flappy_W(37, 357) <= 0; flappy_W(37, 358) <= 0; flappy_W(37, 359) <= 0; flappy_W(37, 360) <= 0; flappy_W(37, 361) <= 0; flappy_W(37, 362) <= 0; flappy_W(37, 363) <= 0; flappy_W(37, 364) <= 0; flappy_W(37, 365) <= 0; flappy_W(37, 366) <= 0; flappy_W(37, 367) <= 0; flappy_W(37, 368) <= 0; flappy_W(37, 369) <= 0; flappy_W(37, 370) <= 0; flappy_W(37, 371) <= 0; flappy_W(37, 372) <= 0; flappy_W(37, 373) <= 0; flappy_W(37, 374) <= 0; flappy_W(37, 375) <= 0; flappy_W(37, 376) <= 0; flappy_W(37, 377) <= 0; flappy_W(37, 378) <= 0; flappy_W(37, 379) <= 0; flappy_W(37, 380) <= 0; flappy_W(37, 381) <= 0; flappy_W(37, 382) <= 0; flappy_W(37, 383) <= 0; flappy_W(37, 384) <= 0; flappy_W(37, 385) <= 0; flappy_W(37, 386) <= 0; flappy_W(37, 387) <= 0; flappy_W(37, 388) <= 0; flappy_W(37, 389) <= 0; flappy_W(37, 390) <= 0; flappy_W(37, 391) <= 0; flappy_W(37, 392) <= 0; flappy_W(37, 393) <= 0; flappy_W(37, 394) <= 0; flappy_W(37, 395) <= 0; flappy_W(37, 396) <= 0; flappy_W(37, 397) <= 0; flappy_W(37, 398) <= 0; flappy_W(37, 399) <= 0; flappy_W(37, 400) <= 0; flappy_W(37, 401) <= 0; flappy_W(37, 402) <= 1; flappy_W(37, 403) <= 1; flappy_W(37, 404) <= 1; flappy_W(37, 405) <= 1; flappy_W(37, 406) <= 1; flappy_W(37, 407) <= 1; flappy_W(37, 408) <= 1; flappy_W(37, 409) <= 1; flappy_W(37, 410) <= 1; flappy_W(37, 411) <= 1; flappy_W(37, 412) <= 1; flappy_W(37, 413) <= 1; flappy_W(37, 414) <= 0; flappy_W(37, 415) <= 0; flappy_W(37, 416) <= 0; flappy_W(37, 417) <= 0; flappy_W(37, 418) <= 0; flappy_W(37, 419) <= 0; flappy_W(37, 420) <= 0; flappy_W(37, 421) <= 0; flappy_W(37, 422) <= 0; flappy_W(37, 423) <= 0; flappy_W(37, 424) <= 0; flappy_W(37, 425) <= 0; flappy_W(37, 426) <= 1; flappy_W(37, 427) <= 1; flappy_W(37, 428) <= 1; flappy_W(37, 429) <= 1; flappy_W(37, 430) <= 1; flappy_W(37, 431) <= 1; flappy_W(37, 432) <= 1; flappy_W(37, 433) <= 1; flappy_W(37, 434) <= 1; flappy_W(37, 435) <= 1; flappy_W(37, 436) <= 1; flappy_W(37, 437) <= 1; flappy_W(37, 438) <= 0; flappy_W(37, 439) <= 0; flappy_W(37, 440) <= 0; flappy_W(37, 441) <= 0; flappy_W(37, 442) <= 0; flappy_W(37, 443) <= 0; flappy_W(37, 444) <= 0; flappy_W(37, 445) <= 0; flappy_W(37, 446) <= 0; flappy_W(37, 447) <= 0; flappy_W(37, 448) <= 0; flappy_W(37, 449) <= 0; flappy_W(37, 450) <= 0; flappy_W(37, 451) <= 0; flappy_W(37, 452) <= 0; flappy_W(37, 453) <= 0; flappy_W(37, 454) <= 0; flappy_W(37, 455) <= 0; flappy_W(37, 456) <= 0; flappy_W(37, 457) <= 0; flappy_W(37, 458) <= 0; flappy_W(37, 459) <= 0; flappy_W(37, 460) <= 0; flappy_W(37, 461) <= 0; flappy_W(37, 462) <= 0; flappy_W(37, 463) <= 0; flappy_W(37, 464) <= 0; flappy_W(37, 465) <= 0; flappy_W(37, 466) <= 0; flappy_W(37, 467) <= 0; flappy_W(37, 468) <= 1; flappy_W(37, 469) <= 1; flappy_W(37, 470) <= 1; flappy_W(37, 471) <= 1; flappy_W(37, 472) <= 1; flappy_W(37, 473) <= 1; flappy_W(37, 474) <= 1; flappy_W(37, 475) <= 1; flappy_W(37, 476) <= 1; flappy_W(37, 477) <= 1; flappy_W(37, 478) <= 1; flappy_W(37, 479) <= 1; flappy_W(37, 480) <= 0; flappy_W(37, 481) <= 0; flappy_W(37, 482) <= 0; flappy_W(37, 483) <= 0; flappy_W(37, 484) <= 0; flappy_W(37, 485) <= 0; flappy_W(37, 486) <= 0; flappy_W(37, 487) <= 0; flappy_W(37, 488) <= 0; flappy_W(37, 489) <= 0; flappy_W(37, 490) <= 0; flappy_W(37, 491) <= 0; flappy_W(37, 492) <= 0; flappy_W(37, 493) <= 0; flappy_W(37, 494) <= 0; flappy_W(37, 495) <= 0; flappy_W(37, 496) <= 0; flappy_W(37, 497) <= 0; flappy_W(37, 498) <= 0; flappy_W(37, 499) <= 0; flappy_W(37, 500) <= 0; flappy_W(37, 501) <= 0; flappy_W(37, 502) <= 0; flappy_W(37, 503) <= 0; flappy_W(37, 504) <= 0; flappy_W(37, 505) <= 0; flappy_W(37, 506) <= 0; flappy_W(37, 507) <= 0; flappy_W(37, 508) <= 0; flappy_W(37, 509) <= 0; flappy_W(37, 510) <= 1; flappy_W(37, 511) <= 1; flappy_W(37, 512) <= 1; flappy_W(37, 513) <= 1; flappy_W(37, 514) <= 1; flappy_W(37, 515) <= 1; flappy_W(37, 516) <= 1; flappy_W(37, 517) <= 1; flappy_W(37, 518) <= 1; flappy_W(37, 519) <= 1; flappy_W(37, 520) <= 1; flappy_W(37, 521) <= 1; flappy_W(37, 522) <= 0; flappy_W(37, 523) <= 0; flappy_W(37, 524) <= 0; flappy_W(37, 525) <= 0; flappy_W(37, 526) <= 0; flappy_W(37, 527) <= 0; flappy_W(37, 528) <= 0; flappy_W(37, 529) <= 0; flappy_W(37, 530) <= 0; flappy_W(37, 531) <= 0; flappy_W(37, 532) <= 0; flappy_W(37, 533) <= 0; flappy_W(37, 534) <= 1; flappy_W(37, 535) <= 1; flappy_W(37, 536) <= 1; flappy_W(37, 537) <= 1; flappy_W(37, 538) <= 1; flappy_W(37, 539) <= 1; flappy_W(37, 540) <= 1; flappy_W(37, 541) <= 1; flappy_W(37, 542) <= 1; flappy_W(37, 543) <= 1; flappy_W(37, 544) <= 1; flappy_W(37, 545) <= 1; flappy_W(37, 546) <= 0; flappy_W(37, 547) <= 0; flappy_W(37, 548) <= 0; flappy_W(37, 549) <= 0; flappy_W(37, 550) <= 0; flappy_W(37, 551) <= 0; flappy_W(37, 552) <= 0; flappy_W(37, 553) <= 0; flappy_W(37, 554) <= 0; flappy_W(37, 555) <= 0; flappy_W(37, 556) <= 0; flappy_W(37, 557) <= 0; flappy_W(37, 558) <= 0; flappy_W(37, 559) <= 0; flappy_W(37, 560) <= 0; flappy_W(37, 561) <= 0; flappy_W(37, 562) <= 0; flappy_W(37, 563) <= 0; flappy_W(37, 564) <= 1; flappy_W(37, 565) <= 1; flappy_W(37, 566) <= 1; flappy_W(37, 567) <= 1; flappy_W(37, 568) <= 1; flappy_W(37, 569) <= 1; flappy_W(37, 570) <= 1; flappy_W(37, 571) <= 1; flappy_W(37, 572) <= 1; flappy_W(37, 573) <= 1; flappy_W(37, 574) <= 1; flappy_W(37, 575) <= 1; flappy_W(37, 576) <= 0; flappy_W(37, 577) <= 0; flappy_W(37, 578) <= 0; flappy_W(37, 579) <= 0; flappy_W(37, 580) <= 0; flappy_W(37, 581) <= 0; flappy_W(37, 582) <= 0; flappy_W(37, 583) <= 0; flappy_W(37, 584) <= 0; flappy_W(37, 585) <= 0; flappy_W(37, 586) <= 0; flappy_W(37, 587) <= 0; flappy_W(37, 588) <= 1; flappy_W(37, 589) <= 1; flappy_W(37, 590) <= 1; flappy_W(37, 591) <= 1; flappy_W(37, 592) <= 1; flappy_W(37, 593) <= 1; 
flappy_W(38, 0) <= 0; flappy_W(38, 1) <= 0; flappy_W(38, 2) <= 0; flappy_W(38, 3) <= 0; flappy_W(38, 4) <= 0; flappy_W(38, 5) <= 0; flappy_W(38, 6) <= 1; flappy_W(38, 7) <= 1; flappy_W(38, 8) <= 1; flappy_W(38, 9) <= 1; flappy_W(38, 10) <= 1; flappy_W(38, 11) <= 1; flappy_W(38, 12) <= 1; flappy_W(38, 13) <= 1; flappy_W(38, 14) <= 1; flappy_W(38, 15) <= 1; flappy_W(38, 16) <= 1; flappy_W(38, 17) <= 1; flappy_W(38, 18) <= 0; flappy_W(38, 19) <= 0; flappy_W(38, 20) <= 0; flappy_W(38, 21) <= 0; flappy_W(38, 22) <= 0; flappy_W(38, 23) <= 0; flappy_W(38, 24) <= 0; flappy_W(38, 25) <= 0; flappy_W(38, 26) <= 0; flappy_W(38, 27) <= 0; flappy_W(38, 28) <= 0; flappy_W(38, 29) <= 0; flappy_W(38, 30) <= 0; flappy_W(38, 31) <= 0; flappy_W(38, 32) <= 0; flappy_W(38, 33) <= 0; flappy_W(38, 34) <= 0; flappy_W(38, 35) <= 0; flappy_W(38, 36) <= 0; flappy_W(38, 37) <= 0; flappy_W(38, 38) <= 0; flappy_W(38, 39) <= 0; flappy_W(38, 40) <= 0; flappy_W(38, 41) <= 0; flappy_W(38, 42) <= 0; flappy_W(38, 43) <= 0; flappy_W(38, 44) <= 0; flappy_W(38, 45) <= 0; flappy_W(38, 46) <= 0; flappy_W(38, 47) <= 0; flappy_W(38, 48) <= 0; flappy_W(38, 49) <= 0; flappy_W(38, 50) <= 0; flappy_W(38, 51) <= 0; flappy_W(38, 52) <= 0; flappy_W(38, 53) <= 0; flappy_W(38, 54) <= 0; flappy_W(38, 55) <= 0; flappy_W(38, 56) <= 0; flappy_W(38, 57) <= 0; flappy_W(38, 58) <= 0; flappy_W(38, 59) <= 0; flappy_W(38, 60) <= 1; flappy_W(38, 61) <= 1; flappy_W(38, 62) <= 1; flappy_W(38, 63) <= 1; flappy_W(38, 64) <= 1; flappy_W(38, 65) <= 1; flappy_W(38, 66) <= 1; flappy_W(38, 67) <= 1; flappy_W(38, 68) <= 1; flappy_W(38, 69) <= 1; flappy_W(38, 70) <= 1; flappy_W(38, 71) <= 1; flappy_W(38, 72) <= 0; flappy_W(38, 73) <= 0; flappy_W(38, 74) <= 0; flappy_W(38, 75) <= 0; flappy_W(38, 76) <= 0; flappy_W(38, 77) <= 0; flappy_W(38, 78) <= 0; flappy_W(38, 79) <= 0; flappy_W(38, 80) <= 0; flappy_W(38, 81) <= 0; flappy_W(38, 82) <= 0; flappy_W(38, 83) <= 0; flappy_W(38, 84) <= 0; flappy_W(38, 85) <= 0; flappy_W(38, 86) <= 0; flappy_W(38, 87) <= 0; flappy_W(38, 88) <= 0; flappy_W(38, 89) <= 0; flappy_W(38, 90) <= 0; flappy_W(38, 91) <= 0; flappy_W(38, 92) <= 0; flappy_W(38, 93) <= 0; flappy_W(38, 94) <= 0; flappy_W(38, 95) <= 0; flappy_W(38, 96) <= 0; flappy_W(38, 97) <= 0; flappy_W(38, 98) <= 0; flappy_W(38, 99) <= 0; flappy_W(38, 100) <= 0; flappy_W(38, 101) <= 0; flappy_W(38, 102) <= 0; flappy_W(38, 103) <= 0; flappy_W(38, 104) <= 0; flappy_W(38, 105) <= 0; flappy_W(38, 106) <= 0; flappy_W(38, 107) <= 0; flappy_W(38, 108) <= 1; flappy_W(38, 109) <= 1; flappy_W(38, 110) <= 1; flappy_W(38, 111) <= 1; flappy_W(38, 112) <= 1; flappy_W(38, 113) <= 1; flappy_W(38, 114) <= 1; flappy_W(38, 115) <= 1; flappy_W(38, 116) <= 1; flappy_W(38, 117) <= 1; flappy_W(38, 118) <= 1; flappy_W(38, 119) <= 1; flappy_W(38, 120) <= 0; flappy_W(38, 121) <= 0; flappy_W(38, 122) <= 0; flappy_W(38, 123) <= 0; flappy_W(38, 124) <= 0; flappy_W(38, 125) <= 0; flappy_W(38, 126) <= 0; flappy_W(38, 127) <= 0; flappy_W(38, 128) <= 0; flappy_W(38, 129) <= 0; flappy_W(38, 130) <= 0; flappy_W(38, 131) <= 0; flappy_W(38, 132) <= 0; flappy_W(38, 133) <= 0; flappy_W(38, 134) <= 0; flappy_W(38, 135) <= 0; flappy_W(38, 136) <= 0; flappy_W(38, 137) <= 0; flappy_W(38, 138) <= 1; flappy_W(38, 139) <= 1; flappy_W(38, 140) <= 1; flappy_W(38, 141) <= 1; flappy_W(38, 142) <= 1; flappy_W(38, 143) <= 1; flappy_W(38, 144) <= 1; flappy_W(38, 145) <= 1; flappy_W(38, 146) <= 1; flappy_W(38, 147) <= 1; flappy_W(38, 148) <= 1; flappy_W(38, 149) <= 1; flappy_W(38, 150) <= 0; flappy_W(38, 151) <= 0; flappy_W(38, 152) <= 0; flappy_W(38, 153) <= 0; flappy_W(38, 154) <= 0; flappy_W(38, 155) <= 0; flappy_W(38, 156) <= 0; flappy_W(38, 157) <= 0; flappy_W(38, 158) <= 0; flappy_W(38, 159) <= 0; flappy_W(38, 160) <= 0; flappy_W(38, 161) <= 0; flappy_W(38, 162) <= 0; flappy_W(38, 163) <= 0; flappy_W(38, 164) <= 0; flappy_W(38, 165) <= 0; flappy_W(38, 166) <= 0; flappy_W(38, 167) <= 0; flappy_W(38, 168) <= 1; flappy_W(38, 169) <= 1; flappy_W(38, 170) <= 1; flappy_W(38, 171) <= 1; flappy_W(38, 172) <= 1; flappy_W(38, 173) <= 1; flappy_W(38, 174) <= 1; flappy_W(38, 175) <= 1; flappy_W(38, 176) <= 1; flappy_W(38, 177) <= 1; flappy_W(38, 178) <= 1; flappy_W(38, 179) <= 1; flappy_W(38, 180) <= 0; flappy_W(38, 181) <= 0; flappy_W(38, 182) <= 0; flappy_W(38, 183) <= 0; flappy_W(38, 184) <= 0; flappy_W(38, 185) <= 0; flappy_W(38, 186) <= 0; flappy_W(38, 187) <= 0; flappy_W(38, 188) <= 0; flappy_W(38, 189) <= 0; flappy_W(38, 190) <= 0; flappy_W(38, 191) <= 0; flappy_W(38, 192) <= 0; flappy_W(38, 193) <= 0; flappy_W(38, 194) <= 0; flappy_W(38, 195) <= 0; flappy_W(38, 196) <= 0; flappy_W(38, 197) <= 0; flappy_W(38, 198) <= 0; flappy_W(38, 199) <= 0; flappy_W(38, 200) <= 0; flappy_W(38, 201) <= 0; flappy_W(38, 202) <= 0; flappy_W(38, 203) <= 0; flappy_W(38, 204) <= 0; flappy_W(38, 205) <= 0; flappy_W(38, 206) <= 0; flappy_W(38, 207) <= 0; flappy_W(38, 208) <= 0; flappy_W(38, 209) <= 0; flappy_W(38, 210) <= 0; flappy_W(38, 211) <= 0; flappy_W(38, 212) <= 0; flappy_W(38, 213) <= 0; flappy_W(38, 214) <= 0; flappy_W(38, 215) <= 0; flappy_W(38, 216) <= 0; flappy_W(38, 217) <= 0; flappy_W(38, 218) <= 0; flappy_W(38, 219) <= 0; flappy_W(38, 220) <= 0; flappy_W(38, 221) <= 0; flappy_W(38, 222) <= 1; flappy_W(38, 223) <= 1; flappy_W(38, 224) <= 1; flappy_W(38, 225) <= 1; flappy_W(38, 226) <= 1; flappy_W(38, 227) <= 1; flappy_W(38, 228) <= 1; flappy_W(38, 229) <= 1; flappy_W(38, 230) <= 1; flappy_W(38, 231) <= 1; flappy_W(38, 232) <= 1; flappy_W(38, 233) <= 1; flappy_W(38, 234) <= 0; flappy_W(38, 235) <= 0; flappy_W(38, 236) <= 0; flappy_W(38, 237) <= 0; flappy_W(38, 238) <= 0; flappy_W(38, 239) <= 0; flappy_W(38, 240) <= 0; flappy_W(38, 241) <= 0; flappy_W(38, 242) <= 0; flappy_W(38, 243) <= 0; flappy_W(38, 244) <= 0; flappy_W(38, 245) <= 0; flappy_W(38, 246) <= 0; flappy_W(38, 247) <= 0; flappy_W(38, 248) <= 0; flappy_W(38, 249) <= 0; flappy_W(38, 250) <= 0; flappy_W(38, 251) <= 0; flappy_W(38, 252) <= 0; flappy_W(38, 253) <= 0; flappy_W(38, 254) <= 0; flappy_W(38, 255) <= 0; flappy_W(38, 256) <= 0; flappy_W(38, 257) <= 0; flappy_W(38, 258) <= 0; flappy_W(38, 259) <= 0; flappy_W(38, 260) <= 0; flappy_W(38, 261) <= 0; flappy_W(38, 262) <= 0; flappy_W(38, 263) <= 0; flappy_W(38, 264) <= 0; flappy_W(38, 265) <= 0; flappy_W(38, 266) <= 0; flappy_W(38, 267) <= 0; flappy_W(38, 268) <= 0; flappy_W(38, 269) <= 0; flappy_W(38, 270) <= 0; flappy_W(38, 271) <= 0; flappy_W(38, 272) <= 0; flappy_W(38, 273) <= 0; flappy_W(38, 274) <= 0; flappy_W(38, 275) <= 0; flappy_W(38, 276) <= 0; flappy_W(38, 277) <= 0; flappy_W(38, 278) <= 0; flappy_W(38, 279) <= 0; flappy_W(38, 280) <= 0; flappy_W(38, 281) <= 0; flappy_W(38, 282) <= 0; flappy_W(38, 283) <= 0; flappy_W(38, 284) <= 0; flappy_W(38, 285) <= 0; flappy_W(38, 286) <= 0; flappy_W(38, 287) <= 0; flappy_W(38, 288) <= 1; flappy_W(38, 289) <= 1; flappy_W(38, 290) <= 1; flappy_W(38, 291) <= 1; flappy_W(38, 292) <= 1; flappy_W(38, 293) <= 1; flappy_W(38, 294) <= 1; flappy_W(38, 295) <= 1; flappy_W(38, 296) <= 1; flappy_W(38, 297) <= 1; flappy_W(38, 298) <= 1; flappy_W(38, 299) <= 1; flappy_W(38, 300) <= 0; flappy_W(38, 301) <= 0; flappy_W(38, 302) <= 0; flappy_W(38, 303) <= 0; flappy_W(38, 304) <= 0; flappy_W(38, 305) <= 0; flappy_W(38, 306) <= 0; flappy_W(38, 307) <= 0; flappy_W(38, 308) <= 0; flappy_W(38, 309) <= 0; flappy_W(38, 310) <= 0; flappy_W(38, 311) <= 0; flappy_W(38, 312) <= 0; flappy_W(38, 313) <= 0; flappy_W(38, 314) <= 0; flappy_W(38, 315) <= 0; flappy_W(38, 316) <= 0; flappy_W(38, 317) <= 0; flappy_W(38, 318) <= 0; flappy_W(38, 319) <= 0; flappy_W(38, 320) <= 0; flappy_W(38, 321) <= 0; flappy_W(38, 322) <= 0; flappy_W(38, 323) <= 0; flappy_W(38, 324) <= 0; flappy_W(38, 325) <= 0; flappy_W(38, 326) <= 0; flappy_W(38, 327) <= 0; flappy_W(38, 328) <= 0; flappy_W(38, 329) <= 0; flappy_W(38, 330) <= 0; flappy_W(38, 331) <= 0; flappy_W(38, 332) <= 0; flappy_W(38, 333) <= 0; flappy_W(38, 334) <= 0; flappy_W(38, 335) <= 0; flappy_W(38, 336) <= 0; flappy_W(38, 337) <= 0; flappy_W(38, 338) <= 0; flappy_W(38, 339) <= 0; flappy_W(38, 340) <= 0; flappy_W(38, 341) <= 0; flappy_W(38, 342) <= 0; flappy_W(38, 343) <= 0; flappy_W(38, 344) <= 0; flappy_W(38, 345) <= 0; flappy_W(38, 346) <= 0; flappy_W(38, 347) <= 0; flappy_W(38, 348) <= 0; flappy_W(38, 349) <= 0; flappy_W(38, 350) <= 0; flappy_W(38, 351) <= 0; flappy_W(38, 352) <= 0; flappy_W(38, 353) <= 0; flappy_W(38, 354) <= 0; flappy_W(38, 355) <= 0; flappy_W(38, 356) <= 0; flappy_W(38, 357) <= 0; flappy_W(38, 358) <= 0; flappy_W(38, 359) <= 0; flappy_W(38, 360) <= 0; flappy_W(38, 361) <= 0; flappy_W(38, 362) <= 0; flappy_W(38, 363) <= 0; flappy_W(38, 364) <= 0; flappy_W(38, 365) <= 0; flappy_W(38, 366) <= 0; flappy_W(38, 367) <= 0; flappy_W(38, 368) <= 0; flappy_W(38, 369) <= 0; flappy_W(38, 370) <= 0; flappy_W(38, 371) <= 0; flappy_W(38, 372) <= 0; flappy_W(38, 373) <= 0; flappy_W(38, 374) <= 0; flappy_W(38, 375) <= 0; flappy_W(38, 376) <= 0; flappy_W(38, 377) <= 0; flappy_W(38, 378) <= 0; flappy_W(38, 379) <= 0; flappy_W(38, 380) <= 0; flappy_W(38, 381) <= 0; flappy_W(38, 382) <= 0; flappy_W(38, 383) <= 0; flappy_W(38, 384) <= 0; flappy_W(38, 385) <= 0; flappy_W(38, 386) <= 0; flappy_W(38, 387) <= 0; flappy_W(38, 388) <= 0; flappy_W(38, 389) <= 0; flappy_W(38, 390) <= 0; flappy_W(38, 391) <= 0; flappy_W(38, 392) <= 0; flappy_W(38, 393) <= 0; flappy_W(38, 394) <= 0; flappy_W(38, 395) <= 0; flappy_W(38, 396) <= 0; flappy_W(38, 397) <= 0; flappy_W(38, 398) <= 0; flappy_W(38, 399) <= 0; flappy_W(38, 400) <= 0; flappy_W(38, 401) <= 0; flappy_W(38, 402) <= 1; flappy_W(38, 403) <= 1; flappy_W(38, 404) <= 1; flappy_W(38, 405) <= 1; flappy_W(38, 406) <= 1; flappy_W(38, 407) <= 1; flappy_W(38, 408) <= 1; flappy_W(38, 409) <= 1; flappy_W(38, 410) <= 1; flappy_W(38, 411) <= 1; flappy_W(38, 412) <= 1; flappy_W(38, 413) <= 1; flappy_W(38, 414) <= 0; flappy_W(38, 415) <= 0; flappy_W(38, 416) <= 0; flappy_W(38, 417) <= 0; flappy_W(38, 418) <= 0; flappy_W(38, 419) <= 0; flappy_W(38, 420) <= 0; flappy_W(38, 421) <= 0; flappy_W(38, 422) <= 0; flappy_W(38, 423) <= 0; flappy_W(38, 424) <= 0; flappy_W(38, 425) <= 0; flappy_W(38, 426) <= 1; flappy_W(38, 427) <= 1; flappy_W(38, 428) <= 1; flappy_W(38, 429) <= 1; flappy_W(38, 430) <= 1; flappy_W(38, 431) <= 1; flappy_W(38, 432) <= 1; flappy_W(38, 433) <= 1; flappy_W(38, 434) <= 1; flappy_W(38, 435) <= 1; flappy_W(38, 436) <= 1; flappy_W(38, 437) <= 1; flappy_W(38, 438) <= 0; flappy_W(38, 439) <= 0; flappy_W(38, 440) <= 0; flappy_W(38, 441) <= 0; flappy_W(38, 442) <= 0; flappy_W(38, 443) <= 0; flappy_W(38, 444) <= 0; flappy_W(38, 445) <= 0; flappy_W(38, 446) <= 0; flappy_W(38, 447) <= 0; flappy_W(38, 448) <= 0; flappy_W(38, 449) <= 0; flappy_W(38, 450) <= 0; flappy_W(38, 451) <= 0; flappy_W(38, 452) <= 0; flappy_W(38, 453) <= 0; flappy_W(38, 454) <= 0; flappy_W(38, 455) <= 0; flappy_W(38, 456) <= 0; flappy_W(38, 457) <= 0; flappy_W(38, 458) <= 0; flappy_W(38, 459) <= 0; flappy_W(38, 460) <= 0; flappy_W(38, 461) <= 0; flappy_W(38, 462) <= 0; flappy_W(38, 463) <= 0; flappy_W(38, 464) <= 0; flappy_W(38, 465) <= 0; flappy_W(38, 466) <= 0; flappy_W(38, 467) <= 0; flappy_W(38, 468) <= 1; flappy_W(38, 469) <= 1; flappy_W(38, 470) <= 1; flappy_W(38, 471) <= 1; flappy_W(38, 472) <= 1; flappy_W(38, 473) <= 1; flappy_W(38, 474) <= 1; flappy_W(38, 475) <= 1; flappy_W(38, 476) <= 1; flappy_W(38, 477) <= 1; flappy_W(38, 478) <= 1; flappy_W(38, 479) <= 1; flappy_W(38, 480) <= 0; flappy_W(38, 481) <= 0; flappy_W(38, 482) <= 0; flappy_W(38, 483) <= 0; flappy_W(38, 484) <= 0; flappy_W(38, 485) <= 0; flappy_W(38, 486) <= 0; flappy_W(38, 487) <= 0; flappy_W(38, 488) <= 0; flappy_W(38, 489) <= 0; flappy_W(38, 490) <= 0; flappy_W(38, 491) <= 0; flappy_W(38, 492) <= 0; flappy_W(38, 493) <= 0; flappy_W(38, 494) <= 0; flappy_W(38, 495) <= 0; flappy_W(38, 496) <= 0; flappy_W(38, 497) <= 0; flappy_W(38, 498) <= 0; flappy_W(38, 499) <= 0; flappy_W(38, 500) <= 0; flappy_W(38, 501) <= 0; flappy_W(38, 502) <= 0; flappy_W(38, 503) <= 0; flappy_W(38, 504) <= 0; flappy_W(38, 505) <= 0; flappy_W(38, 506) <= 0; flappy_W(38, 507) <= 0; flappy_W(38, 508) <= 0; flappy_W(38, 509) <= 0; flappy_W(38, 510) <= 1; flappy_W(38, 511) <= 1; flappy_W(38, 512) <= 1; flappy_W(38, 513) <= 1; flappy_W(38, 514) <= 1; flappy_W(38, 515) <= 1; flappy_W(38, 516) <= 1; flappy_W(38, 517) <= 1; flappy_W(38, 518) <= 1; flappy_W(38, 519) <= 1; flappy_W(38, 520) <= 1; flappy_W(38, 521) <= 1; flappy_W(38, 522) <= 0; flappy_W(38, 523) <= 0; flappy_W(38, 524) <= 0; flappy_W(38, 525) <= 0; flappy_W(38, 526) <= 0; flappy_W(38, 527) <= 0; flappy_W(38, 528) <= 0; flappy_W(38, 529) <= 0; flappy_W(38, 530) <= 0; flappy_W(38, 531) <= 0; flappy_W(38, 532) <= 0; flappy_W(38, 533) <= 0; flappy_W(38, 534) <= 1; flappy_W(38, 535) <= 1; flappy_W(38, 536) <= 1; flappy_W(38, 537) <= 1; flappy_W(38, 538) <= 1; flappy_W(38, 539) <= 1; flappy_W(38, 540) <= 1; flappy_W(38, 541) <= 1; flappy_W(38, 542) <= 1; flappy_W(38, 543) <= 1; flappy_W(38, 544) <= 1; flappy_W(38, 545) <= 1; flappy_W(38, 546) <= 0; flappy_W(38, 547) <= 0; flappy_W(38, 548) <= 0; flappy_W(38, 549) <= 0; flappy_W(38, 550) <= 0; flappy_W(38, 551) <= 0; flappy_W(38, 552) <= 0; flappy_W(38, 553) <= 0; flappy_W(38, 554) <= 0; flappy_W(38, 555) <= 0; flappy_W(38, 556) <= 0; flappy_W(38, 557) <= 0; flappy_W(38, 558) <= 0; flappy_W(38, 559) <= 0; flappy_W(38, 560) <= 0; flappy_W(38, 561) <= 0; flappy_W(38, 562) <= 0; flappy_W(38, 563) <= 0; flappy_W(38, 564) <= 1; flappy_W(38, 565) <= 1; flappy_W(38, 566) <= 1; flappy_W(38, 567) <= 1; flappy_W(38, 568) <= 1; flappy_W(38, 569) <= 1; flappy_W(38, 570) <= 1; flappy_W(38, 571) <= 1; flappy_W(38, 572) <= 1; flappy_W(38, 573) <= 1; flappy_W(38, 574) <= 1; flappy_W(38, 575) <= 1; flappy_W(38, 576) <= 0; flappy_W(38, 577) <= 0; flappy_W(38, 578) <= 0; flappy_W(38, 579) <= 0; flappy_W(38, 580) <= 0; flappy_W(38, 581) <= 0; flappy_W(38, 582) <= 0; flappy_W(38, 583) <= 0; flappy_W(38, 584) <= 0; flappy_W(38, 585) <= 0; flappy_W(38, 586) <= 0; flappy_W(38, 587) <= 0; flappy_W(38, 588) <= 1; flappy_W(38, 589) <= 1; flappy_W(38, 590) <= 1; flappy_W(38, 591) <= 1; flappy_W(38, 592) <= 1; flappy_W(38, 593) <= 1; 
flappy_W(39, 0) <= 0; flappy_W(39, 1) <= 0; flappy_W(39, 2) <= 0; flappy_W(39, 3) <= 0; flappy_W(39, 4) <= 0; flappy_W(39, 5) <= 0; flappy_W(39, 6) <= 1; flappy_W(39, 7) <= 1; flappy_W(39, 8) <= 1; flappy_W(39, 9) <= 1; flappy_W(39, 10) <= 1; flappy_W(39, 11) <= 1; flappy_W(39, 12) <= 1; flappy_W(39, 13) <= 1; flappy_W(39, 14) <= 1; flappy_W(39, 15) <= 1; flappy_W(39, 16) <= 1; flappy_W(39, 17) <= 1; flappy_W(39, 18) <= 0; flappy_W(39, 19) <= 0; flappy_W(39, 20) <= 0; flappy_W(39, 21) <= 0; flappy_W(39, 22) <= 0; flappy_W(39, 23) <= 0; flappy_W(39, 24) <= 0; flappy_W(39, 25) <= 0; flappy_W(39, 26) <= 0; flappy_W(39, 27) <= 0; flappy_W(39, 28) <= 0; flappy_W(39, 29) <= 0; flappy_W(39, 30) <= 0; flappy_W(39, 31) <= 0; flappy_W(39, 32) <= 0; flappy_W(39, 33) <= 0; flappy_W(39, 34) <= 0; flappy_W(39, 35) <= 0; flappy_W(39, 36) <= 0; flappy_W(39, 37) <= 0; flappy_W(39, 38) <= 0; flappy_W(39, 39) <= 0; flappy_W(39, 40) <= 0; flappy_W(39, 41) <= 0; flappy_W(39, 42) <= 0; flappy_W(39, 43) <= 0; flappy_W(39, 44) <= 0; flappy_W(39, 45) <= 0; flappy_W(39, 46) <= 0; flappy_W(39, 47) <= 0; flappy_W(39, 48) <= 0; flappy_W(39, 49) <= 0; flappy_W(39, 50) <= 0; flappy_W(39, 51) <= 0; flappy_W(39, 52) <= 0; flappy_W(39, 53) <= 0; flappy_W(39, 54) <= 0; flappy_W(39, 55) <= 0; flappy_W(39, 56) <= 0; flappy_W(39, 57) <= 0; flappy_W(39, 58) <= 0; flappy_W(39, 59) <= 0; flappy_W(39, 60) <= 1; flappy_W(39, 61) <= 1; flappy_W(39, 62) <= 1; flappy_W(39, 63) <= 1; flappy_W(39, 64) <= 1; flappy_W(39, 65) <= 1; flappy_W(39, 66) <= 1; flappy_W(39, 67) <= 1; flappy_W(39, 68) <= 1; flappy_W(39, 69) <= 1; flappy_W(39, 70) <= 1; flappy_W(39, 71) <= 1; flappy_W(39, 72) <= 0; flappy_W(39, 73) <= 0; flappy_W(39, 74) <= 0; flappy_W(39, 75) <= 0; flappy_W(39, 76) <= 0; flappy_W(39, 77) <= 0; flappy_W(39, 78) <= 0; flappy_W(39, 79) <= 0; flappy_W(39, 80) <= 0; flappy_W(39, 81) <= 0; flappy_W(39, 82) <= 0; flappy_W(39, 83) <= 0; flappy_W(39, 84) <= 0; flappy_W(39, 85) <= 0; flappy_W(39, 86) <= 0; flappy_W(39, 87) <= 0; flappy_W(39, 88) <= 0; flappy_W(39, 89) <= 0; flappy_W(39, 90) <= 0; flappy_W(39, 91) <= 0; flappy_W(39, 92) <= 0; flappy_W(39, 93) <= 0; flappy_W(39, 94) <= 0; flappy_W(39, 95) <= 0; flappy_W(39, 96) <= 0; flappy_W(39, 97) <= 0; flappy_W(39, 98) <= 0; flappy_W(39, 99) <= 0; flappy_W(39, 100) <= 0; flappy_W(39, 101) <= 0; flappy_W(39, 102) <= 0; flappy_W(39, 103) <= 0; flappy_W(39, 104) <= 0; flappy_W(39, 105) <= 0; flappy_W(39, 106) <= 0; flappy_W(39, 107) <= 0; flappy_W(39, 108) <= 1; flappy_W(39, 109) <= 1; flappy_W(39, 110) <= 1; flappy_W(39, 111) <= 1; flappy_W(39, 112) <= 1; flappy_W(39, 113) <= 1; flappy_W(39, 114) <= 1; flappy_W(39, 115) <= 1; flappy_W(39, 116) <= 1; flappy_W(39, 117) <= 1; flappy_W(39, 118) <= 1; flappy_W(39, 119) <= 1; flappy_W(39, 120) <= 0; flappy_W(39, 121) <= 0; flappy_W(39, 122) <= 0; flappy_W(39, 123) <= 0; flappy_W(39, 124) <= 0; flappy_W(39, 125) <= 0; flappy_W(39, 126) <= 0; flappy_W(39, 127) <= 0; flappy_W(39, 128) <= 0; flappy_W(39, 129) <= 0; flappy_W(39, 130) <= 0; flappy_W(39, 131) <= 0; flappy_W(39, 132) <= 0; flappy_W(39, 133) <= 0; flappy_W(39, 134) <= 0; flappy_W(39, 135) <= 0; flappy_W(39, 136) <= 0; flappy_W(39, 137) <= 0; flappy_W(39, 138) <= 1; flappy_W(39, 139) <= 1; flappy_W(39, 140) <= 1; flappy_W(39, 141) <= 1; flappy_W(39, 142) <= 1; flappy_W(39, 143) <= 1; flappy_W(39, 144) <= 1; flappy_W(39, 145) <= 1; flappy_W(39, 146) <= 1; flappy_W(39, 147) <= 1; flappy_W(39, 148) <= 1; flappy_W(39, 149) <= 1; flappy_W(39, 150) <= 0; flappy_W(39, 151) <= 0; flappy_W(39, 152) <= 0; flappy_W(39, 153) <= 0; flappy_W(39, 154) <= 0; flappy_W(39, 155) <= 0; flappy_W(39, 156) <= 0; flappy_W(39, 157) <= 0; flappy_W(39, 158) <= 0; flappy_W(39, 159) <= 0; flappy_W(39, 160) <= 0; flappy_W(39, 161) <= 0; flappy_W(39, 162) <= 0; flappy_W(39, 163) <= 0; flappy_W(39, 164) <= 0; flappy_W(39, 165) <= 0; flappy_W(39, 166) <= 0; flappy_W(39, 167) <= 0; flappy_W(39, 168) <= 1; flappy_W(39, 169) <= 1; flappy_W(39, 170) <= 1; flappy_W(39, 171) <= 1; flappy_W(39, 172) <= 1; flappy_W(39, 173) <= 1; flappy_W(39, 174) <= 1; flappy_W(39, 175) <= 1; flappy_W(39, 176) <= 1; flappy_W(39, 177) <= 1; flappy_W(39, 178) <= 1; flappy_W(39, 179) <= 1; flappy_W(39, 180) <= 0; flappy_W(39, 181) <= 0; flappy_W(39, 182) <= 0; flappy_W(39, 183) <= 0; flappy_W(39, 184) <= 0; flappy_W(39, 185) <= 0; flappy_W(39, 186) <= 0; flappy_W(39, 187) <= 0; flappy_W(39, 188) <= 0; flappy_W(39, 189) <= 0; flappy_W(39, 190) <= 0; flappy_W(39, 191) <= 0; flappy_W(39, 192) <= 0; flappy_W(39, 193) <= 0; flappy_W(39, 194) <= 0; flappy_W(39, 195) <= 0; flappy_W(39, 196) <= 0; flappy_W(39, 197) <= 0; flappy_W(39, 198) <= 0; flappy_W(39, 199) <= 0; flappy_W(39, 200) <= 0; flappy_W(39, 201) <= 0; flappy_W(39, 202) <= 0; flappy_W(39, 203) <= 0; flappy_W(39, 204) <= 0; flappy_W(39, 205) <= 0; flappy_W(39, 206) <= 0; flappy_W(39, 207) <= 0; flappy_W(39, 208) <= 0; flappy_W(39, 209) <= 0; flappy_W(39, 210) <= 0; flappy_W(39, 211) <= 0; flappy_W(39, 212) <= 0; flappy_W(39, 213) <= 0; flappy_W(39, 214) <= 0; flappy_W(39, 215) <= 0; flappy_W(39, 216) <= 0; flappy_W(39, 217) <= 0; flappy_W(39, 218) <= 0; flappy_W(39, 219) <= 0; flappy_W(39, 220) <= 0; flappy_W(39, 221) <= 0; flappy_W(39, 222) <= 1; flappy_W(39, 223) <= 1; flappy_W(39, 224) <= 1; flappy_W(39, 225) <= 1; flappy_W(39, 226) <= 1; flappy_W(39, 227) <= 1; flappy_W(39, 228) <= 1; flappy_W(39, 229) <= 1; flappy_W(39, 230) <= 1; flappy_W(39, 231) <= 1; flappy_W(39, 232) <= 1; flappy_W(39, 233) <= 1; flappy_W(39, 234) <= 0; flappy_W(39, 235) <= 0; flappy_W(39, 236) <= 0; flappy_W(39, 237) <= 0; flappy_W(39, 238) <= 0; flappy_W(39, 239) <= 0; flappy_W(39, 240) <= 0; flappy_W(39, 241) <= 0; flappy_W(39, 242) <= 0; flappy_W(39, 243) <= 0; flappy_W(39, 244) <= 0; flappy_W(39, 245) <= 0; flappy_W(39, 246) <= 0; flappy_W(39, 247) <= 0; flappy_W(39, 248) <= 0; flappy_W(39, 249) <= 0; flappy_W(39, 250) <= 0; flappy_W(39, 251) <= 0; flappy_W(39, 252) <= 0; flappy_W(39, 253) <= 0; flappy_W(39, 254) <= 0; flappy_W(39, 255) <= 0; flappy_W(39, 256) <= 0; flappy_W(39, 257) <= 0; flappy_W(39, 258) <= 0; flappy_W(39, 259) <= 0; flappy_W(39, 260) <= 0; flappy_W(39, 261) <= 0; flappy_W(39, 262) <= 0; flappy_W(39, 263) <= 0; flappy_W(39, 264) <= 0; flappy_W(39, 265) <= 0; flappy_W(39, 266) <= 0; flappy_W(39, 267) <= 0; flappy_W(39, 268) <= 0; flappy_W(39, 269) <= 0; flappy_W(39, 270) <= 0; flappy_W(39, 271) <= 0; flappy_W(39, 272) <= 0; flappy_W(39, 273) <= 0; flappy_W(39, 274) <= 0; flappy_W(39, 275) <= 0; flappy_W(39, 276) <= 0; flappy_W(39, 277) <= 0; flappy_W(39, 278) <= 0; flappy_W(39, 279) <= 0; flappy_W(39, 280) <= 0; flappy_W(39, 281) <= 0; flappy_W(39, 282) <= 0; flappy_W(39, 283) <= 0; flappy_W(39, 284) <= 0; flappy_W(39, 285) <= 0; flappy_W(39, 286) <= 0; flappy_W(39, 287) <= 0; flappy_W(39, 288) <= 1; flappy_W(39, 289) <= 1; flappy_W(39, 290) <= 1; flappy_W(39, 291) <= 1; flappy_W(39, 292) <= 1; flappy_W(39, 293) <= 1; flappy_W(39, 294) <= 1; flappy_W(39, 295) <= 1; flappy_W(39, 296) <= 1; flappy_W(39, 297) <= 1; flappy_W(39, 298) <= 1; flappy_W(39, 299) <= 1; flappy_W(39, 300) <= 0; flappy_W(39, 301) <= 0; flappy_W(39, 302) <= 0; flappy_W(39, 303) <= 0; flappy_W(39, 304) <= 0; flappy_W(39, 305) <= 0; flappy_W(39, 306) <= 0; flappy_W(39, 307) <= 0; flappy_W(39, 308) <= 0; flappy_W(39, 309) <= 0; flappy_W(39, 310) <= 0; flappy_W(39, 311) <= 0; flappy_W(39, 312) <= 0; flappy_W(39, 313) <= 0; flappy_W(39, 314) <= 0; flappy_W(39, 315) <= 0; flappy_W(39, 316) <= 0; flappy_W(39, 317) <= 0; flappy_W(39, 318) <= 0; flappy_W(39, 319) <= 0; flappy_W(39, 320) <= 0; flappy_W(39, 321) <= 0; flappy_W(39, 322) <= 0; flappy_W(39, 323) <= 0; flappy_W(39, 324) <= 0; flappy_W(39, 325) <= 0; flappy_W(39, 326) <= 0; flappy_W(39, 327) <= 0; flappy_W(39, 328) <= 0; flappy_W(39, 329) <= 0; flappy_W(39, 330) <= 0; flappy_W(39, 331) <= 0; flappy_W(39, 332) <= 0; flappy_W(39, 333) <= 0; flappy_W(39, 334) <= 0; flappy_W(39, 335) <= 0; flappy_W(39, 336) <= 0; flappy_W(39, 337) <= 0; flappy_W(39, 338) <= 0; flappy_W(39, 339) <= 0; flappy_W(39, 340) <= 0; flappy_W(39, 341) <= 0; flappy_W(39, 342) <= 0; flappy_W(39, 343) <= 0; flappy_W(39, 344) <= 0; flappy_W(39, 345) <= 0; flappy_W(39, 346) <= 0; flappy_W(39, 347) <= 0; flappy_W(39, 348) <= 0; flappy_W(39, 349) <= 0; flappy_W(39, 350) <= 0; flappy_W(39, 351) <= 0; flappy_W(39, 352) <= 0; flappy_W(39, 353) <= 0; flappy_W(39, 354) <= 0; flappy_W(39, 355) <= 0; flappy_W(39, 356) <= 0; flappy_W(39, 357) <= 0; flappy_W(39, 358) <= 0; flappy_W(39, 359) <= 0; flappy_W(39, 360) <= 0; flappy_W(39, 361) <= 0; flappy_W(39, 362) <= 0; flappy_W(39, 363) <= 0; flappy_W(39, 364) <= 0; flappy_W(39, 365) <= 0; flappy_W(39, 366) <= 0; flappy_W(39, 367) <= 0; flappy_W(39, 368) <= 0; flappy_W(39, 369) <= 0; flappy_W(39, 370) <= 0; flappy_W(39, 371) <= 0; flappy_W(39, 372) <= 0; flappy_W(39, 373) <= 0; flappy_W(39, 374) <= 0; flappy_W(39, 375) <= 0; flappy_W(39, 376) <= 0; flappy_W(39, 377) <= 0; flappy_W(39, 378) <= 0; flappy_W(39, 379) <= 0; flappy_W(39, 380) <= 0; flappy_W(39, 381) <= 0; flappy_W(39, 382) <= 0; flappy_W(39, 383) <= 0; flappy_W(39, 384) <= 0; flappy_W(39, 385) <= 0; flappy_W(39, 386) <= 0; flappy_W(39, 387) <= 0; flappy_W(39, 388) <= 0; flappy_W(39, 389) <= 0; flappy_W(39, 390) <= 0; flappy_W(39, 391) <= 0; flappy_W(39, 392) <= 0; flappy_W(39, 393) <= 0; flappy_W(39, 394) <= 0; flappy_W(39, 395) <= 0; flappy_W(39, 396) <= 0; flappy_W(39, 397) <= 0; flappy_W(39, 398) <= 0; flappy_W(39, 399) <= 0; flappy_W(39, 400) <= 0; flappy_W(39, 401) <= 0; flappy_W(39, 402) <= 1; flappy_W(39, 403) <= 1; flappy_W(39, 404) <= 1; flappy_W(39, 405) <= 1; flappy_W(39, 406) <= 1; flappy_W(39, 407) <= 1; flappy_W(39, 408) <= 1; flappy_W(39, 409) <= 1; flappy_W(39, 410) <= 1; flappy_W(39, 411) <= 1; flappy_W(39, 412) <= 1; flappy_W(39, 413) <= 1; flappy_W(39, 414) <= 0; flappy_W(39, 415) <= 0; flappy_W(39, 416) <= 0; flappy_W(39, 417) <= 0; flappy_W(39, 418) <= 0; flappy_W(39, 419) <= 0; flappy_W(39, 420) <= 0; flappy_W(39, 421) <= 0; flappy_W(39, 422) <= 0; flappy_W(39, 423) <= 0; flappy_W(39, 424) <= 0; flappy_W(39, 425) <= 0; flappy_W(39, 426) <= 1; flappy_W(39, 427) <= 1; flappy_W(39, 428) <= 1; flappy_W(39, 429) <= 1; flappy_W(39, 430) <= 1; flappy_W(39, 431) <= 1; flappy_W(39, 432) <= 1; flappy_W(39, 433) <= 1; flappy_W(39, 434) <= 1; flappy_W(39, 435) <= 1; flappy_W(39, 436) <= 1; flappy_W(39, 437) <= 1; flappy_W(39, 438) <= 0; flappy_W(39, 439) <= 0; flappy_W(39, 440) <= 0; flappy_W(39, 441) <= 0; flappy_W(39, 442) <= 0; flappy_W(39, 443) <= 0; flappy_W(39, 444) <= 0; flappy_W(39, 445) <= 0; flappy_W(39, 446) <= 0; flappy_W(39, 447) <= 0; flappy_W(39, 448) <= 0; flappy_W(39, 449) <= 0; flappy_W(39, 450) <= 0; flappy_W(39, 451) <= 0; flappy_W(39, 452) <= 0; flappy_W(39, 453) <= 0; flappy_W(39, 454) <= 0; flappy_W(39, 455) <= 0; flappy_W(39, 456) <= 0; flappy_W(39, 457) <= 0; flappy_W(39, 458) <= 0; flappy_W(39, 459) <= 0; flappy_W(39, 460) <= 0; flappy_W(39, 461) <= 0; flappy_W(39, 462) <= 0; flappy_W(39, 463) <= 0; flappy_W(39, 464) <= 0; flappy_W(39, 465) <= 0; flappy_W(39, 466) <= 0; flappy_W(39, 467) <= 0; flappy_W(39, 468) <= 1; flappy_W(39, 469) <= 1; flappy_W(39, 470) <= 1; flappy_W(39, 471) <= 1; flappy_W(39, 472) <= 1; flappy_W(39, 473) <= 1; flappy_W(39, 474) <= 1; flappy_W(39, 475) <= 1; flappy_W(39, 476) <= 1; flappy_W(39, 477) <= 1; flappy_W(39, 478) <= 1; flappy_W(39, 479) <= 1; flappy_W(39, 480) <= 0; flappy_W(39, 481) <= 0; flappy_W(39, 482) <= 0; flappy_W(39, 483) <= 0; flappy_W(39, 484) <= 0; flappy_W(39, 485) <= 0; flappy_W(39, 486) <= 0; flappy_W(39, 487) <= 0; flappy_W(39, 488) <= 0; flappy_W(39, 489) <= 0; flappy_W(39, 490) <= 0; flappy_W(39, 491) <= 0; flappy_W(39, 492) <= 0; flappy_W(39, 493) <= 0; flappy_W(39, 494) <= 0; flappy_W(39, 495) <= 0; flappy_W(39, 496) <= 0; flappy_W(39, 497) <= 0; flappy_W(39, 498) <= 0; flappy_W(39, 499) <= 0; flappy_W(39, 500) <= 0; flappy_W(39, 501) <= 0; flappy_W(39, 502) <= 0; flappy_W(39, 503) <= 0; flappy_W(39, 504) <= 0; flappy_W(39, 505) <= 0; flappy_W(39, 506) <= 0; flappy_W(39, 507) <= 0; flappy_W(39, 508) <= 0; flappy_W(39, 509) <= 0; flappy_W(39, 510) <= 1; flappy_W(39, 511) <= 1; flappy_W(39, 512) <= 1; flappy_W(39, 513) <= 1; flappy_W(39, 514) <= 1; flappy_W(39, 515) <= 1; flappy_W(39, 516) <= 1; flappy_W(39, 517) <= 1; flappy_W(39, 518) <= 1; flappy_W(39, 519) <= 1; flappy_W(39, 520) <= 1; flappy_W(39, 521) <= 1; flappy_W(39, 522) <= 0; flappy_W(39, 523) <= 0; flappy_W(39, 524) <= 0; flappy_W(39, 525) <= 0; flappy_W(39, 526) <= 0; flappy_W(39, 527) <= 0; flappy_W(39, 528) <= 0; flappy_W(39, 529) <= 0; flappy_W(39, 530) <= 0; flappy_W(39, 531) <= 0; flappy_W(39, 532) <= 0; flappy_W(39, 533) <= 0; flappy_W(39, 534) <= 1; flappy_W(39, 535) <= 1; flappy_W(39, 536) <= 1; flappy_W(39, 537) <= 1; flappy_W(39, 538) <= 1; flappy_W(39, 539) <= 1; flappy_W(39, 540) <= 1; flappy_W(39, 541) <= 1; flappy_W(39, 542) <= 1; flappy_W(39, 543) <= 1; flappy_W(39, 544) <= 1; flappy_W(39, 545) <= 1; flappy_W(39, 546) <= 0; flappy_W(39, 547) <= 0; flappy_W(39, 548) <= 0; flappy_W(39, 549) <= 0; flappy_W(39, 550) <= 0; flappy_W(39, 551) <= 0; flappy_W(39, 552) <= 0; flappy_W(39, 553) <= 0; flappy_W(39, 554) <= 0; flappy_W(39, 555) <= 0; flappy_W(39, 556) <= 0; flappy_W(39, 557) <= 0; flappy_W(39, 558) <= 0; flappy_W(39, 559) <= 0; flappy_W(39, 560) <= 0; flappy_W(39, 561) <= 0; flappy_W(39, 562) <= 0; flappy_W(39, 563) <= 0; flappy_W(39, 564) <= 1; flappy_W(39, 565) <= 1; flappy_W(39, 566) <= 1; flappy_W(39, 567) <= 1; flappy_W(39, 568) <= 1; flappy_W(39, 569) <= 1; flappy_W(39, 570) <= 1; flappy_W(39, 571) <= 1; flappy_W(39, 572) <= 1; flappy_W(39, 573) <= 1; flappy_W(39, 574) <= 1; flappy_W(39, 575) <= 1; flappy_W(39, 576) <= 0; flappy_W(39, 577) <= 0; flappy_W(39, 578) <= 0; flappy_W(39, 579) <= 0; flappy_W(39, 580) <= 0; flappy_W(39, 581) <= 0; flappy_W(39, 582) <= 0; flappy_W(39, 583) <= 0; flappy_W(39, 584) <= 0; flappy_W(39, 585) <= 0; flappy_W(39, 586) <= 0; flappy_W(39, 587) <= 0; flappy_W(39, 588) <= 1; flappy_W(39, 589) <= 1; flappy_W(39, 590) <= 1; flappy_W(39, 591) <= 1; flappy_W(39, 592) <= 1; flappy_W(39, 593) <= 1; 
flappy_W(40, 0) <= 0; flappy_W(40, 1) <= 0; flappy_W(40, 2) <= 0; flappy_W(40, 3) <= 0; flappy_W(40, 4) <= 0; flappy_W(40, 5) <= 0; flappy_W(40, 6) <= 1; flappy_W(40, 7) <= 1; flappy_W(40, 8) <= 1; flappy_W(40, 9) <= 1; flappy_W(40, 10) <= 1; flappy_W(40, 11) <= 1; flappy_W(40, 12) <= 1; flappy_W(40, 13) <= 1; flappy_W(40, 14) <= 1; flappy_W(40, 15) <= 1; flappy_W(40, 16) <= 1; flappy_W(40, 17) <= 1; flappy_W(40, 18) <= 0; flappy_W(40, 19) <= 0; flappy_W(40, 20) <= 0; flappy_W(40, 21) <= 0; flappy_W(40, 22) <= 0; flappy_W(40, 23) <= 0; flappy_W(40, 24) <= 0; flappy_W(40, 25) <= 0; flappy_W(40, 26) <= 0; flappy_W(40, 27) <= 0; flappy_W(40, 28) <= 0; flappy_W(40, 29) <= 0; flappy_W(40, 30) <= 0; flappy_W(40, 31) <= 0; flappy_W(40, 32) <= 0; flappy_W(40, 33) <= 0; flappy_W(40, 34) <= 0; flappy_W(40, 35) <= 0; flappy_W(40, 36) <= 0; flappy_W(40, 37) <= 0; flappy_W(40, 38) <= 0; flappy_W(40, 39) <= 0; flappy_W(40, 40) <= 0; flappy_W(40, 41) <= 0; flappy_W(40, 42) <= 0; flappy_W(40, 43) <= 0; flappy_W(40, 44) <= 0; flappy_W(40, 45) <= 0; flappy_W(40, 46) <= 0; flappy_W(40, 47) <= 0; flappy_W(40, 48) <= 0; flappy_W(40, 49) <= 0; flappy_W(40, 50) <= 0; flappy_W(40, 51) <= 0; flappy_W(40, 52) <= 0; flappy_W(40, 53) <= 0; flappy_W(40, 54) <= 0; flappy_W(40, 55) <= 0; flappy_W(40, 56) <= 0; flappy_W(40, 57) <= 0; flappy_W(40, 58) <= 0; flappy_W(40, 59) <= 0; flappy_W(40, 60) <= 1; flappy_W(40, 61) <= 1; flappy_W(40, 62) <= 1; flappy_W(40, 63) <= 1; flappy_W(40, 64) <= 1; flappy_W(40, 65) <= 1; flappy_W(40, 66) <= 1; flappy_W(40, 67) <= 1; flappy_W(40, 68) <= 1; flappy_W(40, 69) <= 1; flappy_W(40, 70) <= 1; flappy_W(40, 71) <= 1; flappy_W(40, 72) <= 0; flappy_W(40, 73) <= 0; flappy_W(40, 74) <= 0; flappy_W(40, 75) <= 0; flappy_W(40, 76) <= 0; flappy_W(40, 77) <= 0; flappy_W(40, 78) <= 0; flappy_W(40, 79) <= 0; flappy_W(40, 80) <= 0; flappy_W(40, 81) <= 0; flappy_W(40, 82) <= 0; flappy_W(40, 83) <= 0; flappy_W(40, 84) <= 0; flappy_W(40, 85) <= 0; flappy_W(40, 86) <= 0; flappy_W(40, 87) <= 0; flappy_W(40, 88) <= 0; flappy_W(40, 89) <= 0; flappy_W(40, 90) <= 0; flappy_W(40, 91) <= 0; flappy_W(40, 92) <= 0; flappy_W(40, 93) <= 0; flappy_W(40, 94) <= 0; flappy_W(40, 95) <= 0; flappy_W(40, 96) <= 0; flappy_W(40, 97) <= 0; flappy_W(40, 98) <= 0; flappy_W(40, 99) <= 0; flappy_W(40, 100) <= 0; flappy_W(40, 101) <= 0; flappy_W(40, 102) <= 0; flappy_W(40, 103) <= 0; flappy_W(40, 104) <= 0; flappy_W(40, 105) <= 0; flappy_W(40, 106) <= 0; flappy_W(40, 107) <= 0; flappy_W(40, 108) <= 1; flappy_W(40, 109) <= 1; flappy_W(40, 110) <= 1; flappy_W(40, 111) <= 1; flappy_W(40, 112) <= 1; flappy_W(40, 113) <= 1; flappy_W(40, 114) <= 1; flappy_W(40, 115) <= 1; flappy_W(40, 116) <= 1; flappy_W(40, 117) <= 1; flappy_W(40, 118) <= 1; flappy_W(40, 119) <= 1; flappy_W(40, 120) <= 0; flappy_W(40, 121) <= 0; flappy_W(40, 122) <= 0; flappy_W(40, 123) <= 0; flappy_W(40, 124) <= 0; flappy_W(40, 125) <= 0; flappy_W(40, 126) <= 0; flappy_W(40, 127) <= 0; flappy_W(40, 128) <= 0; flappy_W(40, 129) <= 0; flappy_W(40, 130) <= 0; flappy_W(40, 131) <= 0; flappy_W(40, 132) <= 0; flappy_W(40, 133) <= 0; flappy_W(40, 134) <= 0; flappy_W(40, 135) <= 0; flappy_W(40, 136) <= 0; flappy_W(40, 137) <= 0; flappy_W(40, 138) <= 1; flappy_W(40, 139) <= 1; flappy_W(40, 140) <= 1; flappy_W(40, 141) <= 1; flappy_W(40, 142) <= 1; flappy_W(40, 143) <= 1; flappy_W(40, 144) <= 1; flappy_W(40, 145) <= 1; flappy_W(40, 146) <= 1; flappy_W(40, 147) <= 1; flappy_W(40, 148) <= 1; flappy_W(40, 149) <= 1; flappy_W(40, 150) <= 0; flappy_W(40, 151) <= 0; flappy_W(40, 152) <= 0; flappy_W(40, 153) <= 0; flappy_W(40, 154) <= 0; flappy_W(40, 155) <= 0; flappy_W(40, 156) <= 0; flappy_W(40, 157) <= 0; flappy_W(40, 158) <= 0; flappy_W(40, 159) <= 0; flappy_W(40, 160) <= 0; flappy_W(40, 161) <= 0; flappy_W(40, 162) <= 0; flappy_W(40, 163) <= 0; flappy_W(40, 164) <= 0; flappy_W(40, 165) <= 0; flappy_W(40, 166) <= 0; flappy_W(40, 167) <= 0; flappy_W(40, 168) <= 1; flappy_W(40, 169) <= 1; flappy_W(40, 170) <= 1; flappy_W(40, 171) <= 1; flappy_W(40, 172) <= 1; flappy_W(40, 173) <= 1; flappy_W(40, 174) <= 1; flappy_W(40, 175) <= 1; flappy_W(40, 176) <= 1; flappy_W(40, 177) <= 1; flappy_W(40, 178) <= 1; flappy_W(40, 179) <= 1; flappy_W(40, 180) <= 0; flappy_W(40, 181) <= 0; flappy_W(40, 182) <= 0; flappy_W(40, 183) <= 0; flappy_W(40, 184) <= 0; flappy_W(40, 185) <= 0; flappy_W(40, 186) <= 0; flappy_W(40, 187) <= 0; flappy_W(40, 188) <= 0; flappy_W(40, 189) <= 0; flappy_W(40, 190) <= 0; flappy_W(40, 191) <= 0; flappy_W(40, 192) <= 0; flappy_W(40, 193) <= 0; flappy_W(40, 194) <= 0; flappy_W(40, 195) <= 0; flappy_W(40, 196) <= 0; flappy_W(40, 197) <= 0; flappy_W(40, 198) <= 0; flappy_W(40, 199) <= 0; flappy_W(40, 200) <= 0; flappy_W(40, 201) <= 0; flappy_W(40, 202) <= 0; flappy_W(40, 203) <= 0; flappy_W(40, 204) <= 0; flappy_W(40, 205) <= 0; flappy_W(40, 206) <= 0; flappy_W(40, 207) <= 0; flappy_W(40, 208) <= 0; flappy_W(40, 209) <= 0; flappy_W(40, 210) <= 0; flappy_W(40, 211) <= 0; flappy_W(40, 212) <= 0; flappy_W(40, 213) <= 0; flappy_W(40, 214) <= 0; flappy_W(40, 215) <= 0; flappy_W(40, 216) <= 0; flappy_W(40, 217) <= 0; flappy_W(40, 218) <= 0; flappy_W(40, 219) <= 0; flappy_W(40, 220) <= 0; flappy_W(40, 221) <= 0; flappy_W(40, 222) <= 1; flappy_W(40, 223) <= 1; flappy_W(40, 224) <= 1; flappy_W(40, 225) <= 1; flappy_W(40, 226) <= 1; flappy_W(40, 227) <= 1; flappy_W(40, 228) <= 1; flappy_W(40, 229) <= 1; flappy_W(40, 230) <= 1; flappy_W(40, 231) <= 1; flappy_W(40, 232) <= 1; flappy_W(40, 233) <= 1; flappy_W(40, 234) <= 0; flappy_W(40, 235) <= 0; flappy_W(40, 236) <= 0; flappy_W(40, 237) <= 0; flappy_W(40, 238) <= 0; flappy_W(40, 239) <= 0; flappy_W(40, 240) <= 0; flappy_W(40, 241) <= 0; flappy_W(40, 242) <= 0; flappy_W(40, 243) <= 0; flappy_W(40, 244) <= 0; flappy_W(40, 245) <= 0; flappy_W(40, 246) <= 0; flappy_W(40, 247) <= 0; flappy_W(40, 248) <= 0; flappy_W(40, 249) <= 0; flappy_W(40, 250) <= 0; flappy_W(40, 251) <= 0; flappy_W(40, 252) <= 0; flappy_W(40, 253) <= 0; flappy_W(40, 254) <= 0; flappy_W(40, 255) <= 0; flappy_W(40, 256) <= 0; flappy_W(40, 257) <= 0; flappy_W(40, 258) <= 0; flappy_W(40, 259) <= 0; flappy_W(40, 260) <= 0; flappy_W(40, 261) <= 0; flappy_W(40, 262) <= 0; flappy_W(40, 263) <= 0; flappy_W(40, 264) <= 0; flappy_W(40, 265) <= 0; flappy_W(40, 266) <= 0; flappy_W(40, 267) <= 0; flappy_W(40, 268) <= 0; flappy_W(40, 269) <= 0; flappy_W(40, 270) <= 0; flappy_W(40, 271) <= 0; flappy_W(40, 272) <= 0; flappy_W(40, 273) <= 0; flappy_W(40, 274) <= 0; flappy_W(40, 275) <= 0; flappy_W(40, 276) <= 0; flappy_W(40, 277) <= 0; flappy_W(40, 278) <= 0; flappy_W(40, 279) <= 0; flappy_W(40, 280) <= 0; flappy_W(40, 281) <= 0; flappy_W(40, 282) <= 0; flappy_W(40, 283) <= 0; flappy_W(40, 284) <= 0; flappy_W(40, 285) <= 0; flappy_W(40, 286) <= 0; flappy_W(40, 287) <= 0; flappy_W(40, 288) <= 1; flappy_W(40, 289) <= 1; flappy_W(40, 290) <= 1; flappy_W(40, 291) <= 1; flappy_W(40, 292) <= 1; flappy_W(40, 293) <= 1; flappy_W(40, 294) <= 1; flappy_W(40, 295) <= 1; flappy_W(40, 296) <= 1; flappy_W(40, 297) <= 1; flappy_W(40, 298) <= 1; flappy_W(40, 299) <= 1; flappy_W(40, 300) <= 0; flappy_W(40, 301) <= 0; flappy_W(40, 302) <= 0; flappy_W(40, 303) <= 0; flappy_W(40, 304) <= 0; flappy_W(40, 305) <= 0; flappy_W(40, 306) <= 0; flappy_W(40, 307) <= 0; flappy_W(40, 308) <= 0; flappy_W(40, 309) <= 0; flappy_W(40, 310) <= 0; flappy_W(40, 311) <= 0; flappy_W(40, 312) <= 0; flappy_W(40, 313) <= 0; flappy_W(40, 314) <= 0; flappy_W(40, 315) <= 0; flappy_W(40, 316) <= 0; flappy_W(40, 317) <= 0; flappy_W(40, 318) <= 0; flappy_W(40, 319) <= 0; flappy_W(40, 320) <= 0; flappy_W(40, 321) <= 0; flappy_W(40, 322) <= 0; flappy_W(40, 323) <= 0; flappy_W(40, 324) <= 0; flappy_W(40, 325) <= 0; flappy_W(40, 326) <= 0; flappy_W(40, 327) <= 0; flappy_W(40, 328) <= 0; flappy_W(40, 329) <= 0; flappy_W(40, 330) <= 0; flappy_W(40, 331) <= 0; flappy_W(40, 332) <= 0; flappy_W(40, 333) <= 0; flappy_W(40, 334) <= 0; flappy_W(40, 335) <= 0; flappy_W(40, 336) <= 0; flappy_W(40, 337) <= 0; flappy_W(40, 338) <= 0; flappy_W(40, 339) <= 0; flappy_W(40, 340) <= 0; flappy_W(40, 341) <= 0; flappy_W(40, 342) <= 0; flappy_W(40, 343) <= 0; flappy_W(40, 344) <= 0; flappy_W(40, 345) <= 0; flappy_W(40, 346) <= 0; flappy_W(40, 347) <= 0; flappy_W(40, 348) <= 0; flappy_W(40, 349) <= 0; flappy_W(40, 350) <= 0; flappy_W(40, 351) <= 0; flappy_W(40, 352) <= 0; flappy_W(40, 353) <= 0; flappy_W(40, 354) <= 0; flappy_W(40, 355) <= 0; flappy_W(40, 356) <= 0; flappy_W(40, 357) <= 0; flappy_W(40, 358) <= 0; flappy_W(40, 359) <= 0; flappy_W(40, 360) <= 0; flappy_W(40, 361) <= 0; flappy_W(40, 362) <= 0; flappy_W(40, 363) <= 0; flappy_W(40, 364) <= 0; flappy_W(40, 365) <= 0; flappy_W(40, 366) <= 0; flappy_W(40, 367) <= 0; flappy_W(40, 368) <= 0; flappy_W(40, 369) <= 0; flappy_W(40, 370) <= 0; flappy_W(40, 371) <= 0; flappy_W(40, 372) <= 0; flappy_W(40, 373) <= 0; flappy_W(40, 374) <= 0; flappy_W(40, 375) <= 0; flappy_W(40, 376) <= 0; flappy_W(40, 377) <= 0; flappy_W(40, 378) <= 0; flappy_W(40, 379) <= 0; flappy_W(40, 380) <= 0; flappy_W(40, 381) <= 0; flappy_W(40, 382) <= 0; flappy_W(40, 383) <= 0; flappy_W(40, 384) <= 0; flappy_W(40, 385) <= 0; flappy_W(40, 386) <= 0; flappy_W(40, 387) <= 0; flappy_W(40, 388) <= 0; flappy_W(40, 389) <= 0; flappy_W(40, 390) <= 0; flappy_W(40, 391) <= 0; flappy_W(40, 392) <= 0; flappy_W(40, 393) <= 0; flappy_W(40, 394) <= 0; flappy_W(40, 395) <= 0; flappy_W(40, 396) <= 0; flappy_W(40, 397) <= 0; flappy_W(40, 398) <= 0; flappy_W(40, 399) <= 0; flappy_W(40, 400) <= 0; flappy_W(40, 401) <= 0; flappy_W(40, 402) <= 1; flappy_W(40, 403) <= 1; flappy_W(40, 404) <= 1; flappy_W(40, 405) <= 1; flappy_W(40, 406) <= 1; flappy_W(40, 407) <= 1; flappy_W(40, 408) <= 1; flappy_W(40, 409) <= 1; flappy_W(40, 410) <= 1; flappy_W(40, 411) <= 1; flappy_W(40, 412) <= 1; flappy_W(40, 413) <= 1; flappy_W(40, 414) <= 0; flappy_W(40, 415) <= 0; flappy_W(40, 416) <= 0; flappy_W(40, 417) <= 0; flappy_W(40, 418) <= 0; flappy_W(40, 419) <= 0; flappy_W(40, 420) <= 0; flappy_W(40, 421) <= 0; flappy_W(40, 422) <= 0; flappy_W(40, 423) <= 0; flappy_W(40, 424) <= 0; flappy_W(40, 425) <= 0; flappy_W(40, 426) <= 1; flappy_W(40, 427) <= 1; flappy_W(40, 428) <= 1; flappy_W(40, 429) <= 1; flappy_W(40, 430) <= 1; flappy_W(40, 431) <= 1; flappy_W(40, 432) <= 1; flappy_W(40, 433) <= 1; flappy_W(40, 434) <= 1; flappy_W(40, 435) <= 1; flappy_W(40, 436) <= 1; flappy_W(40, 437) <= 1; flappy_W(40, 438) <= 0; flappy_W(40, 439) <= 0; flappy_W(40, 440) <= 0; flappy_W(40, 441) <= 0; flappy_W(40, 442) <= 0; flappy_W(40, 443) <= 0; flappy_W(40, 444) <= 0; flappy_W(40, 445) <= 0; flappy_W(40, 446) <= 0; flappy_W(40, 447) <= 0; flappy_W(40, 448) <= 0; flappy_W(40, 449) <= 0; flappy_W(40, 450) <= 0; flappy_W(40, 451) <= 0; flappy_W(40, 452) <= 0; flappy_W(40, 453) <= 0; flappy_W(40, 454) <= 0; flappy_W(40, 455) <= 0; flappy_W(40, 456) <= 0; flappy_W(40, 457) <= 0; flappy_W(40, 458) <= 0; flappy_W(40, 459) <= 0; flappy_W(40, 460) <= 0; flappy_W(40, 461) <= 0; flappy_W(40, 462) <= 0; flappy_W(40, 463) <= 0; flappy_W(40, 464) <= 0; flappy_W(40, 465) <= 0; flappy_W(40, 466) <= 0; flappy_W(40, 467) <= 0; flappy_W(40, 468) <= 1; flappy_W(40, 469) <= 1; flappy_W(40, 470) <= 1; flappy_W(40, 471) <= 1; flappy_W(40, 472) <= 1; flappy_W(40, 473) <= 1; flappy_W(40, 474) <= 1; flappy_W(40, 475) <= 1; flappy_W(40, 476) <= 1; flappy_W(40, 477) <= 1; flappy_W(40, 478) <= 1; flappy_W(40, 479) <= 1; flappy_W(40, 480) <= 0; flappy_W(40, 481) <= 0; flappy_W(40, 482) <= 0; flappy_W(40, 483) <= 0; flappy_W(40, 484) <= 0; flappy_W(40, 485) <= 0; flappy_W(40, 486) <= 0; flappy_W(40, 487) <= 0; flappy_W(40, 488) <= 0; flappy_W(40, 489) <= 0; flappy_W(40, 490) <= 0; flappy_W(40, 491) <= 0; flappy_W(40, 492) <= 0; flappy_W(40, 493) <= 0; flappy_W(40, 494) <= 0; flappy_W(40, 495) <= 0; flappy_W(40, 496) <= 0; flappy_W(40, 497) <= 0; flappy_W(40, 498) <= 0; flappy_W(40, 499) <= 0; flappy_W(40, 500) <= 0; flappy_W(40, 501) <= 0; flappy_W(40, 502) <= 0; flappy_W(40, 503) <= 0; flappy_W(40, 504) <= 0; flappy_W(40, 505) <= 0; flappy_W(40, 506) <= 0; flappy_W(40, 507) <= 0; flappy_W(40, 508) <= 0; flappy_W(40, 509) <= 0; flappy_W(40, 510) <= 1; flappy_W(40, 511) <= 1; flappy_W(40, 512) <= 1; flappy_W(40, 513) <= 1; flappy_W(40, 514) <= 1; flappy_W(40, 515) <= 1; flappy_W(40, 516) <= 1; flappy_W(40, 517) <= 1; flappy_W(40, 518) <= 1; flappy_W(40, 519) <= 1; flappy_W(40, 520) <= 1; flappy_W(40, 521) <= 1; flappy_W(40, 522) <= 0; flappy_W(40, 523) <= 0; flappy_W(40, 524) <= 0; flappy_W(40, 525) <= 0; flappy_W(40, 526) <= 0; flappy_W(40, 527) <= 0; flappy_W(40, 528) <= 0; flappy_W(40, 529) <= 0; flappy_W(40, 530) <= 0; flappy_W(40, 531) <= 0; flappy_W(40, 532) <= 0; flappy_W(40, 533) <= 0; flappy_W(40, 534) <= 1; flappy_W(40, 535) <= 1; flappy_W(40, 536) <= 1; flappy_W(40, 537) <= 1; flappy_W(40, 538) <= 1; flappy_W(40, 539) <= 1; flappy_W(40, 540) <= 1; flappy_W(40, 541) <= 1; flappy_W(40, 542) <= 1; flappy_W(40, 543) <= 1; flappy_W(40, 544) <= 1; flappy_W(40, 545) <= 1; flappy_W(40, 546) <= 0; flappy_W(40, 547) <= 0; flappy_W(40, 548) <= 0; flappy_W(40, 549) <= 0; flappy_W(40, 550) <= 0; flappy_W(40, 551) <= 0; flappy_W(40, 552) <= 0; flappy_W(40, 553) <= 0; flappy_W(40, 554) <= 0; flappy_W(40, 555) <= 0; flappy_W(40, 556) <= 0; flappy_W(40, 557) <= 0; flappy_W(40, 558) <= 0; flappy_W(40, 559) <= 0; flappy_W(40, 560) <= 0; flappy_W(40, 561) <= 0; flappy_W(40, 562) <= 0; flappy_W(40, 563) <= 0; flappy_W(40, 564) <= 1; flappy_W(40, 565) <= 1; flappy_W(40, 566) <= 1; flappy_W(40, 567) <= 1; flappy_W(40, 568) <= 1; flappy_W(40, 569) <= 1; flappy_W(40, 570) <= 1; flappy_W(40, 571) <= 1; flappy_W(40, 572) <= 1; flappy_W(40, 573) <= 1; flappy_W(40, 574) <= 1; flappy_W(40, 575) <= 1; flappy_W(40, 576) <= 0; flappy_W(40, 577) <= 0; flappy_W(40, 578) <= 0; flappy_W(40, 579) <= 0; flappy_W(40, 580) <= 0; flappy_W(40, 581) <= 0; flappy_W(40, 582) <= 0; flappy_W(40, 583) <= 0; flappy_W(40, 584) <= 0; flappy_W(40, 585) <= 0; flappy_W(40, 586) <= 0; flappy_W(40, 587) <= 0; flappy_W(40, 588) <= 1; flappy_W(40, 589) <= 1; flappy_W(40, 590) <= 1; flappy_W(40, 591) <= 1; flappy_W(40, 592) <= 1; flappy_W(40, 593) <= 1; 
flappy_W(41, 0) <= 0; flappy_W(41, 1) <= 0; flappy_W(41, 2) <= 0; flappy_W(41, 3) <= 0; flappy_W(41, 4) <= 0; flappy_W(41, 5) <= 0; flappy_W(41, 6) <= 1; flappy_W(41, 7) <= 1; flappy_W(41, 8) <= 1; flappy_W(41, 9) <= 1; flappy_W(41, 10) <= 1; flappy_W(41, 11) <= 1; flappy_W(41, 12) <= 1; flappy_W(41, 13) <= 1; flappy_W(41, 14) <= 1; flappy_W(41, 15) <= 1; flappy_W(41, 16) <= 1; flappy_W(41, 17) <= 1; flappy_W(41, 18) <= 0; flappy_W(41, 19) <= 0; flappy_W(41, 20) <= 0; flappy_W(41, 21) <= 0; flappy_W(41, 22) <= 0; flappy_W(41, 23) <= 0; flappy_W(41, 24) <= 0; flappy_W(41, 25) <= 0; flappy_W(41, 26) <= 0; flappy_W(41, 27) <= 0; flappy_W(41, 28) <= 0; flappy_W(41, 29) <= 0; flappy_W(41, 30) <= 0; flappy_W(41, 31) <= 0; flappy_W(41, 32) <= 0; flappy_W(41, 33) <= 0; flappy_W(41, 34) <= 0; flappy_W(41, 35) <= 0; flappy_W(41, 36) <= 0; flappy_W(41, 37) <= 0; flappy_W(41, 38) <= 0; flappy_W(41, 39) <= 0; flappy_W(41, 40) <= 0; flappy_W(41, 41) <= 0; flappy_W(41, 42) <= 0; flappy_W(41, 43) <= 0; flappy_W(41, 44) <= 0; flappy_W(41, 45) <= 0; flappy_W(41, 46) <= 0; flappy_W(41, 47) <= 0; flappy_W(41, 48) <= 0; flappy_W(41, 49) <= 0; flappy_W(41, 50) <= 0; flappy_W(41, 51) <= 0; flappy_W(41, 52) <= 0; flappy_W(41, 53) <= 0; flappy_W(41, 54) <= 0; flappy_W(41, 55) <= 0; flappy_W(41, 56) <= 0; flappy_W(41, 57) <= 0; flappy_W(41, 58) <= 0; flappy_W(41, 59) <= 0; flappy_W(41, 60) <= 1; flappy_W(41, 61) <= 1; flappy_W(41, 62) <= 1; flappy_W(41, 63) <= 1; flappy_W(41, 64) <= 1; flappy_W(41, 65) <= 1; flappy_W(41, 66) <= 1; flappy_W(41, 67) <= 1; flappy_W(41, 68) <= 1; flappy_W(41, 69) <= 1; flappy_W(41, 70) <= 1; flappy_W(41, 71) <= 1; flappy_W(41, 72) <= 0; flappy_W(41, 73) <= 0; flappy_W(41, 74) <= 0; flappy_W(41, 75) <= 0; flappy_W(41, 76) <= 0; flappy_W(41, 77) <= 0; flappy_W(41, 78) <= 0; flappy_W(41, 79) <= 0; flappy_W(41, 80) <= 0; flappy_W(41, 81) <= 0; flappy_W(41, 82) <= 0; flappy_W(41, 83) <= 0; flappy_W(41, 84) <= 0; flappy_W(41, 85) <= 0; flappy_W(41, 86) <= 0; flappy_W(41, 87) <= 0; flappy_W(41, 88) <= 0; flappy_W(41, 89) <= 0; flappy_W(41, 90) <= 0; flappy_W(41, 91) <= 0; flappy_W(41, 92) <= 0; flappy_W(41, 93) <= 0; flappy_W(41, 94) <= 0; flappy_W(41, 95) <= 0; flappy_W(41, 96) <= 0; flappy_W(41, 97) <= 0; flappy_W(41, 98) <= 0; flappy_W(41, 99) <= 0; flappy_W(41, 100) <= 0; flappy_W(41, 101) <= 0; flappy_W(41, 102) <= 0; flappy_W(41, 103) <= 0; flappy_W(41, 104) <= 0; flappy_W(41, 105) <= 0; flappy_W(41, 106) <= 0; flappy_W(41, 107) <= 0; flappy_W(41, 108) <= 1; flappy_W(41, 109) <= 1; flappy_W(41, 110) <= 1; flappy_W(41, 111) <= 1; flappy_W(41, 112) <= 1; flappy_W(41, 113) <= 1; flappy_W(41, 114) <= 1; flappy_W(41, 115) <= 1; flappy_W(41, 116) <= 1; flappy_W(41, 117) <= 1; flappy_W(41, 118) <= 1; flappy_W(41, 119) <= 1; flappy_W(41, 120) <= 0; flappy_W(41, 121) <= 0; flappy_W(41, 122) <= 0; flappy_W(41, 123) <= 0; flappy_W(41, 124) <= 0; flappy_W(41, 125) <= 0; flappy_W(41, 126) <= 0; flappy_W(41, 127) <= 0; flappy_W(41, 128) <= 0; flappy_W(41, 129) <= 0; flappy_W(41, 130) <= 0; flappy_W(41, 131) <= 0; flappy_W(41, 132) <= 0; flappy_W(41, 133) <= 0; flappy_W(41, 134) <= 0; flappy_W(41, 135) <= 0; flappy_W(41, 136) <= 0; flappy_W(41, 137) <= 0; flappy_W(41, 138) <= 1; flappy_W(41, 139) <= 1; flappy_W(41, 140) <= 1; flappy_W(41, 141) <= 1; flappy_W(41, 142) <= 1; flappy_W(41, 143) <= 1; flappy_W(41, 144) <= 1; flappy_W(41, 145) <= 1; flappy_W(41, 146) <= 1; flappy_W(41, 147) <= 1; flappy_W(41, 148) <= 1; flappy_W(41, 149) <= 1; flappy_W(41, 150) <= 0; flappy_W(41, 151) <= 0; flappy_W(41, 152) <= 0; flappy_W(41, 153) <= 0; flappy_W(41, 154) <= 0; flappy_W(41, 155) <= 0; flappy_W(41, 156) <= 0; flappy_W(41, 157) <= 0; flappy_W(41, 158) <= 0; flappy_W(41, 159) <= 0; flappy_W(41, 160) <= 0; flappy_W(41, 161) <= 0; flappy_W(41, 162) <= 0; flappy_W(41, 163) <= 0; flappy_W(41, 164) <= 0; flappy_W(41, 165) <= 0; flappy_W(41, 166) <= 0; flappy_W(41, 167) <= 0; flappy_W(41, 168) <= 1; flappy_W(41, 169) <= 1; flappy_W(41, 170) <= 1; flappy_W(41, 171) <= 1; flappy_W(41, 172) <= 1; flappy_W(41, 173) <= 1; flappy_W(41, 174) <= 1; flappy_W(41, 175) <= 1; flappy_W(41, 176) <= 1; flappy_W(41, 177) <= 1; flappy_W(41, 178) <= 1; flappy_W(41, 179) <= 1; flappy_W(41, 180) <= 0; flappy_W(41, 181) <= 0; flappy_W(41, 182) <= 0; flappy_W(41, 183) <= 0; flappy_W(41, 184) <= 0; flappy_W(41, 185) <= 0; flappy_W(41, 186) <= 0; flappy_W(41, 187) <= 0; flappy_W(41, 188) <= 0; flappy_W(41, 189) <= 0; flappy_W(41, 190) <= 0; flappy_W(41, 191) <= 0; flappy_W(41, 192) <= 0; flappy_W(41, 193) <= 0; flappy_W(41, 194) <= 0; flappy_W(41, 195) <= 0; flappy_W(41, 196) <= 0; flappy_W(41, 197) <= 0; flappy_W(41, 198) <= 0; flappy_W(41, 199) <= 0; flappy_W(41, 200) <= 0; flappy_W(41, 201) <= 0; flappy_W(41, 202) <= 0; flappy_W(41, 203) <= 0; flappy_W(41, 204) <= 0; flappy_W(41, 205) <= 0; flappy_W(41, 206) <= 0; flappy_W(41, 207) <= 0; flappy_W(41, 208) <= 0; flappy_W(41, 209) <= 0; flappy_W(41, 210) <= 0; flappy_W(41, 211) <= 0; flappy_W(41, 212) <= 0; flappy_W(41, 213) <= 0; flappy_W(41, 214) <= 0; flappy_W(41, 215) <= 0; flappy_W(41, 216) <= 0; flappy_W(41, 217) <= 0; flappy_W(41, 218) <= 0; flappy_W(41, 219) <= 0; flappy_W(41, 220) <= 0; flappy_W(41, 221) <= 0; flappy_W(41, 222) <= 1; flappy_W(41, 223) <= 1; flappy_W(41, 224) <= 1; flappy_W(41, 225) <= 1; flappy_W(41, 226) <= 1; flappy_W(41, 227) <= 1; flappy_W(41, 228) <= 1; flappy_W(41, 229) <= 1; flappy_W(41, 230) <= 1; flappy_W(41, 231) <= 1; flappy_W(41, 232) <= 1; flappy_W(41, 233) <= 1; flappy_W(41, 234) <= 0; flappy_W(41, 235) <= 0; flappy_W(41, 236) <= 0; flappy_W(41, 237) <= 0; flappy_W(41, 238) <= 0; flappy_W(41, 239) <= 0; flappy_W(41, 240) <= 0; flappy_W(41, 241) <= 0; flappy_W(41, 242) <= 0; flappy_W(41, 243) <= 0; flappy_W(41, 244) <= 0; flappy_W(41, 245) <= 0; flappy_W(41, 246) <= 0; flappy_W(41, 247) <= 0; flappy_W(41, 248) <= 0; flappy_W(41, 249) <= 0; flappy_W(41, 250) <= 0; flappy_W(41, 251) <= 0; flappy_W(41, 252) <= 0; flappy_W(41, 253) <= 0; flappy_W(41, 254) <= 0; flappy_W(41, 255) <= 0; flappy_W(41, 256) <= 0; flappy_W(41, 257) <= 0; flappy_W(41, 258) <= 0; flappy_W(41, 259) <= 0; flappy_W(41, 260) <= 0; flappy_W(41, 261) <= 0; flappy_W(41, 262) <= 0; flappy_W(41, 263) <= 0; flappy_W(41, 264) <= 0; flappy_W(41, 265) <= 0; flappy_W(41, 266) <= 0; flappy_W(41, 267) <= 0; flappy_W(41, 268) <= 0; flappy_W(41, 269) <= 0; flappy_W(41, 270) <= 0; flappy_W(41, 271) <= 0; flappy_W(41, 272) <= 0; flappy_W(41, 273) <= 0; flappy_W(41, 274) <= 0; flappy_W(41, 275) <= 0; flappy_W(41, 276) <= 0; flappy_W(41, 277) <= 0; flappy_W(41, 278) <= 0; flappy_W(41, 279) <= 0; flappy_W(41, 280) <= 0; flappy_W(41, 281) <= 0; flappy_W(41, 282) <= 0; flappy_W(41, 283) <= 0; flappy_W(41, 284) <= 0; flappy_W(41, 285) <= 0; flappy_W(41, 286) <= 0; flappy_W(41, 287) <= 0; flappy_W(41, 288) <= 1; flappy_W(41, 289) <= 1; flappy_W(41, 290) <= 1; flappy_W(41, 291) <= 1; flappy_W(41, 292) <= 1; flappy_W(41, 293) <= 1; flappy_W(41, 294) <= 1; flappy_W(41, 295) <= 1; flappy_W(41, 296) <= 1; flappy_W(41, 297) <= 1; flappy_W(41, 298) <= 1; flappy_W(41, 299) <= 1; flappy_W(41, 300) <= 0; flappy_W(41, 301) <= 0; flappy_W(41, 302) <= 0; flappy_W(41, 303) <= 0; flappy_W(41, 304) <= 0; flappy_W(41, 305) <= 0; flappy_W(41, 306) <= 0; flappy_W(41, 307) <= 0; flappy_W(41, 308) <= 0; flappy_W(41, 309) <= 0; flappy_W(41, 310) <= 0; flappy_W(41, 311) <= 0; flappy_W(41, 312) <= 0; flappy_W(41, 313) <= 0; flappy_W(41, 314) <= 0; flappy_W(41, 315) <= 0; flappy_W(41, 316) <= 0; flappy_W(41, 317) <= 0; flappy_W(41, 318) <= 0; flappy_W(41, 319) <= 0; flappy_W(41, 320) <= 0; flappy_W(41, 321) <= 0; flappy_W(41, 322) <= 0; flappy_W(41, 323) <= 0; flappy_W(41, 324) <= 0; flappy_W(41, 325) <= 0; flappy_W(41, 326) <= 0; flappy_W(41, 327) <= 0; flappy_W(41, 328) <= 0; flappy_W(41, 329) <= 0; flappy_W(41, 330) <= 0; flappy_W(41, 331) <= 0; flappy_W(41, 332) <= 0; flappy_W(41, 333) <= 0; flappy_W(41, 334) <= 0; flappy_W(41, 335) <= 0; flappy_W(41, 336) <= 0; flappy_W(41, 337) <= 0; flappy_W(41, 338) <= 0; flappy_W(41, 339) <= 0; flappy_W(41, 340) <= 0; flappy_W(41, 341) <= 0; flappy_W(41, 342) <= 0; flappy_W(41, 343) <= 0; flappy_W(41, 344) <= 0; flappy_W(41, 345) <= 0; flappy_W(41, 346) <= 0; flappy_W(41, 347) <= 0; flappy_W(41, 348) <= 0; flappy_W(41, 349) <= 0; flappy_W(41, 350) <= 0; flappy_W(41, 351) <= 0; flappy_W(41, 352) <= 0; flappy_W(41, 353) <= 0; flappy_W(41, 354) <= 0; flappy_W(41, 355) <= 0; flappy_W(41, 356) <= 0; flappy_W(41, 357) <= 0; flappy_W(41, 358) <= 0; flappy_W(41, 359) <= 0; flappy_W(41, 360) <= 0; flappy_W(41, 361) <= 0; flappy_W(41, 362) <= 0; flappy_W(41, 363) <= 0; flappy_W(41, 364) <= 0; flappy_W(41, 365) <= 0; flappy_W(41, 366) <= 0; flappy_W(41, 367) <= 0; flappy_W(41, 368) <= 0; flappy_W(41, 369) <= 0; flappy_W(41, 370) <= 0; flappy_W(41, 371) <= 0; flappy_W(41, 372) <= 0; flappy_W(41, 373) <= 0; flappy_W(41, 374) <= 0; flappy_W(41, 375) <= 0; flappy_W(41, 376) <= 0; flappy_W(41, 377) <= 0; flappy_W(41, 378) <= 0; flappy_W(41, 379) <= 0; flappy_W(41, 380) <= 0; flappy_W(41, 381) <= 0; flappy_W(41, 382) <= 0; flappy_W(41, 383) <= 0; flappy_W(41, 384) <= 0; flappy_W(41, 385) <= 0; flappy_W(41, 386) <= 0; flappy_W(41, 387) <= 0; flappy_W(41, 388) <= 0; flappy_W(41, 389) <= 0; flappy_W(41, 390) <= 0; flappy_W(41, 391) <= 0; flappy_W(41, 392) <= 0; flappy_W(41, 393) <= 0; flappy_W(41, 394) <= 0; flappy_W(41, 395) <= 0; flappy_W(41, 396) <= 0; flappy_W(41, 397) <= 0; flappy_W(41, 398) <= 0; flappy_W(41, 399) <= 0; flappy_W(41, 400) <= 0; flappy_W(41, 401) <= 0; flappy_W(41, 402) <= 1; flappy_W(41, 403) <= 1; flappy_W(41, 404) <= 1; flappy_W(41, 405) <= 1; flappy_W(41, 406) <= 1; flappy_W(41, 407) <= 1; flappy_W(41, 408) <= 1; flappy_W(41, 409) <= 1; flappy_W(41, 410) <= 1; flappy_W(41, 411) <= 1; flappy_W(41, 412) <= 1; flappy_W(41, 413) <= 1; flappy_W(41, 414) <= 0; flappy_W(41, 415) <= 0; flappy_W(41, 416) <= 0; flappy_W(41, 417) <= 0; flappy_W(41, 418) <= 0; flappy_W(41, 419) <= 0; flappy_W(41, 420) <= 0; flappy_W(41, 421) <= 0; flappy_W(41, 422) <= 0; flappy_W(41, 423) <= 0; flappy_W(41, 424) <= 0; flappy_W(41, 425) <= 0; flappy_W(41, 426) <= 1; flappy_W(41, 427) <= 1; flappy_W(41, 428) <= 1; flappy_W(41, 429) <= 1; flappy_W(41, 430) <= 1; flappy_W(41, 431) <= 1; flappy_W(41, 432) <= 1; flappy_W(41, 433) <= 1; flappy_W(41, 434) <= 1; flappy_W(41, 435) <= 1; flappy_W(41, 436) <= 1; flappy_W(41, 437) <= 1; flappy_W(41, 438) <= 0; flappy_W(41, 439) <= 0; flappy_W(41, 440) <= 0; flappy_W(41, 441) <= 0; flappy_W(41, 442) <= 0; flappy_W(41, 443) <= 0; flappy_W(41, 444) <= 0; flappy_W(41, 445) <= 0; flappy_W(41, 446) <= 0; flappy_W(41, 447) <= 0; flappy_W(41, 448) <= 0; flappy_W(41, 449) <= 0; flappy_W(41, 450) <= 0; flappy_W(41, 451) <= 0; flappy_W(41, 452) <= 0; flappy_W(41, 453) <= 0; flappy_W(41, 454) <= 0; flappy_W(41, 455) <= 0; flappy_W(41, 456) <= 0; flappy_W(41, 457) <= 0; flappy_W(41, 458) <= 0; flappy_W(41, 459) <= 0; flappy_W(41, 460) <= 0; flappy_W(41, 461) <= 0; flappy_W(41, 462) <= 0; flappy_W(41, 463) <= 0; flappy_W(41, 464) <= 0; flappy_W(41, 465) <= 0; flappy_W(41, 466) <= 0; flappy_W(41, 467) <= 0; flappy_W(41, 468) <= 1; flappy_W(41, 469) <= 1; flappy_W(41, 470) <= 1; flappy_W(41, 471) <= 1; flappy_W(41, 472) <= 1; flappy_W(41, 473) <= 1; flappy_W(41, 474) <= 1; flappy_W(41, 475) <= 1; flappy_W(41, 476) <= 1; flappy_W(41, 477) <= 1; flappy_W(41, 478) <= 1; flappy_W(41, 479) <= 1; flappy_W(41, 480) <= 0; flappy_W(41, 481) <= 0; flappy_W(41, 482) <= 0; flappy_W(41, 483) <= 0; flappy_W(41, 484) <= 0; flappy_W(41, 485) <= 0; flappy_W(41, 486) <= 0; flappy_W(41, 487) <= 0; flappy_W(41, 488) <= 0; flappy_W(41, 489) <= 0; flappy_W(41, 490) <= 0; flappy_W(41, 491) <= 0; flappy_W(41, 492) <= 0; flappy_W(41, 493) <= 0; flappy_W(41, 494) <= 0; flappy_W(41, 495) <= 0; flappy_W(41, 496) <= 0; flappy_W(41, 497) <= 0; flappy_W(41, 498) <= 0; flappy_W(41, 499) <= 0; flappy_W(41, 500) <= 0; flappy_W(41, 501) <= 0; flappy_W(41, 502) <= 0; flappy_W(41, 503) <= 0; flappy_W(41, 504) <= 0; flappy_W(41, 505) <= 0; flappy_W(41, 506) <= 0; flappy_W(41, 507) <= 0; flappy_W(41, 508) <= 0; flappy_W(41, 509) <= 0; flappy_W(41, 510) <= 1; flappy_W(41, 511) <= 1; flappy_W(41, 512) <= 1; flappy_W(41, 513) <= 1; flappy_W(41, 514) <= 1; flappy_W(41, 515) <= 1; flappy_W(41, 516) <= 1; flappy_W(41, 517) <= 1; flappy_W(41, 518) <= 1; flappy_W(41, 519) <= 1; flappy_W(41, 520) <= 1; flappy_W(41, 521) <= 1; flappy_W(41, 522) <= 0; flappy_W(41, 523) <= 0; flappy_W(41, 524) <= 0; flappy_W(41, 525) <= 0; flappy_W(41, 526) <= 0; flappy_W(41, 527) <= 0; flappy_W(41, 528) <= 0; flappy_W(41, 529) <= 0; flappy_W(41, 530) <= 0; flappy_W(41, 531) <= 0; flappy_W(41, 532) <= 0; flappy_W(41, 533) <= 0; flappy_W(41, 534) <= 1; flappy_W(41, 535) <= 1; flappy_W(41, 536) <= 1; flappy_W(41, 537) <= 1; flappy_W(41, 538) <= 1; flappy_W(41, 539) <= 1; flappy_W(41, 540) <= 1; flappy_W(41, 541) <= 1; flappy_W(41, 542) <= 1; flappy_W(41, 543) <= 1; flappy_W(41, 544) <= 1; flappy_W(41, 545) <= 1; flappy_W(41, 546) <= 0; flappy_W(41, 547) <= 0; flappy_W(41, 548) <= 0; flappy_W(41, 549) <= 0; flappy_W(41, 550) <= 0; flappy_W(41, 551) <= 0; flappy_W(41, 552) <= 0; flappy_W(41, 553) <= 0; flappy_W(41, 554) <= 0; flappy_W(41, 555) <= 0; flappy_W(41, 556) <= 0; flappy_W(41, 557) <= 0; flappy_W(41, 558) <= 0; flappy_W(41, 559) <= 0; flappy_W(41, 560) <= 0; flappy_W(41, 561) <= 0; flappy_W(41, 562) <= 0; flappy_W(41, 563) <= 0; flappy_W(41, 564) <= 1; flappy_W(41, 565) <= 1; flappy_W(41, 566) <= 1; flappy_W(41, 567) <= 1; flappy_W(41, 568) <= 1; flappy_W(41, 569) <= 1; flappy_W(41, 570) <= 1; flappy_W(41, 571) <= 1; flappy_W(41, 572) <= 1; flappy_W(41, 573) <= 1; flappy_W(41, 574) <= 1; flappy_W(41, 575) <= 1; flappy_W(41, 576) <= 0; flappy_W(41, 577) <= 0; flappy_W(41, 578) <= 0; flappy_W(41, 579) <= 0; flappy_W(41, 580) <= 0; flappy_W(41, 581) <= 0; flappy_W(41, 582) <= 0; flappy_W(41, 583) <= 0; flappy_W(41, 584) <= 0; flappy_W(41, 585) <= 0; flappy_W(41, 586) <= 0; flappy_W(41, 587) <= 0; flappy_W(41, 588) <= 1; flappy_W(41, 589) <= 1; flappy_W(41, 590) <= 1; flappy_W(41, 591) <= 1; flappy_W(41, 592) <= 1; flappy_W(41, 593) <= 1; 
flappy_W(42, 0) <= 0; flappy_W(42, 1) <= 0; flappy_W(42, 2) <= 0; flappy_W(42, 3) <= 0; flappy_W(42, 4) <= 0; flappy_W(42, 5) <= 0; flappy_W(42, 6) <= 1; flappy_W(42, 7) <= 1; flappy_W(42, 8) <= 1; flappy_W(42, 9) <= 1; flappy_W(42, 10) <= 1; flappy_W(42, 11) <= 1; flappy_W(42, 12) <= 1; flappy_W(42, 13) <= 1; flappy_W(42, 14) <= 1; flappy_W(42, 15) <= 1; flappy_W(42, 16) <= 1; flappy_W(42, 17) <= 1; flappy_W(42, 18) <= 0; flappy_W(42, 19) <= 0; flappy_W(42, 20) <= 0; flappy_W(42, 21) <= 0; flappy_W(42, 22) <= 0; flappy_W(42, 23) <= 0; flappy_W(42, 24) <= 0; flappy_W(42, 25) <= 0; flappy_W(42, 26) <= 0; flappy_W(42, 27) <= 0; flappy_W(42, 28) <= 0; flappy_W(42, 29) <= 0; flappy_W(42, 30) <= 0; flappy_W(42, 31) <= 0; flappy_W(42, 32) <= 0; flappy_W(42, 33) <= 0; flappy_W(42, 34) <= 0; flappy_W(42, 35) <= 0; flappy_W(42, 36) <= 0; flappy_W(42, 37) <= 0; flappy_W(42, 38) <= 0; flappy_W(42, 39) <= 0; flappy_W(42, 40) <= 0; flappy_W(42, 41) <= 0; flappy_W(42, 42) <= 0; flappy_W(42, 43) <= 0; flappy_W(42, 44) <= 0; flappy_W(42, 45) <= 0; flappy_W(42, 46) <= 0; flappy_W(42, 47) <= 0; flappy_W(42, 48) <= 0; flappy_W(42, 49) <= 0; flappy_W(42, 50) <= 0; flappy_W(42, 51) <= 0; flappy_W(42, 52) <= 0; flappy_W(42, 53) <= 0; flappy_W(42, 54) <= 0; flappy_W(42, 55) <= 0; flappy_W(42, 56) <= 0; flappy_W(42, 57) <= 0; flappy_W(42, 58) <= 0; flappy_W(42, 59) <= 0; flappy_W(42, 60) <= 1; flappy_W(42, 61) <= 1; flappy_W(42, 62) <= 1; flappy_W(42, 63) <= 1; flappy_W(42, 64) <= 1; flappy_W(42, 65) <= 1; flappy_W(42, 66) <= 1; flappy_W(42, 67) <= 1; flappy_W(42, 68) <= 1; flappy_W(42, 69) <= 1; flappy_W(42, 70) <= 1; flappy_W(42, 71) <= 1; flappy_W(42, 72) <= 0; flappy_W(42, 73) <= 0; flappy_W(42, 74) <= 0; flappy_W(42, 75) <= 0; flappy_W(42, 76) <= 0; flappy_W(42, 77) <= 0; flappy_W(42, 78) <= 0; flappy_W(42, 79) <= 0; flappy_W(42, 80) <= 0; flappy_W(42, 81) <= 0; flappy_W(42, 82) <= 0; flappy_W(42, 83) <= 0; flappy_W(42, 84) <= 0; flappy_W(42, 85) <= 0; flappy_W(42, 86) <= 0; flappy_W(42, 87) <= 0; flappy_W(42, 88) <= 0; flappy_W(42, 89) <= 0; flappy_W(42, 90) <= 1; flappy_W(42, 91) <= 1; flappy_W(42, 92) <= 1; flappy_W(42, 93) <= 1; flappy_W(42, 94) <= 1; flappy_W(42, 95) <= 1; flappy_W(42, 96) <= 0; flappy_W(42, 97) <= 0; flappy_W(42, 98) <= 0; flappy_W(42, 99) <= 0; flappy_W(42, 100) <= 0; flappy_W(42, 101) <= 0; flappy_W(42, 102) <= 0; flappy_W(42, 103) <= 0; flappy_W(42, 104) <= 0; flappy_W(42, 105) <= 0; flappy_W(42, 106) <= 0; flappy_W(42, 107) <= 0; flappy_W(42, 108) <= 1; flappy_W(42, 109) <= 1; flappy_W(42, 110) <= 1; flappy_W(42, 111) <= 1; flappy_W(42, 112) <= 1; flappy_W(42, 113) <= 1; flappy_W(42, 114) <= 1; flappy_W(42, 115) <= 1; flappy_W(42, 116) <= 1; flappy_W(42, 117) <= 1; flappy_W(42, 118) <= 1; flappy_W(42, 119) <= 1; flappy_W(42, 120) <= 0; flappy_W(42, 121) <= 0; flappy_W(42, 122) <= 0; flappy_W(42, 123) <= 0; flappy_W(42, 124) <= 0; flappy_W(42, 125) <= 0; flappy_W(42, 126) <= 0; flappy_W(42, 127) <= 0; flappy_W(42, 128) <= 0; flappy_W(42, 129) <= 0; flappy_W(42, 130) <= 0; flappy_W(42, 131) <= 0; flappy_W(42, 132) <= 0; flappy_W(42, 133) <= 0; flappy_W(42, 134) <= 0; flappy_W(42, 135) <= 0; flappy_W(42, 136) <= 0; flappy_W(42, 137) <= 0; flappy_W(42, 138) <= 1; flappy_W(42, 139) <= 1; flappy_W(42, 140) <= 1; flappy_W(42, 141) <= 1; flappy_W(42, 142) <= 1; flappy_W(42, 143) <= 1; flappy_W(42, 144) <= 1; flappy_W(42, 145) <= 1; flappy_W(42, 146) <= 1; flappy_W(42, 147) <= 1; flappy_W(42, 148) <= 1; flappy_W(42, 149) <= 1; flappy_W(42, 150) <= 0; flappy_W(42, 151) <= 0; flappy_W(42, 152) <= 0; flappy_W(42, 153) <= 0; flappy_W(42, 154) <= 0; flappy_W(42, 155) <= 0; flappy_W(42, 156) <= 0; flappy_W(42, 157) <= 0; flappy_W(42, 158) <= 0; flappy_W(42, 159) <= 0; flappy_W(42, 160) <= 0; flappy_W(42, 161) <= 0; flappy_W(42, 162) <= 0; flappy_W(42, 163) <= 0; flappy_W(42, 164) <= 0; flappy_W(42, 165) <= 0; flappy_W(42, 166) <= 0; flappy_W(42, 167) <= 0; flappy_W(42, 168) <= 1; flappy_W(42, 169) <= 1; flappy_W(42, 170) <= 1; flappy_W(42, 171) <= 1; flappy_W(42, 172) <= 1; flappy_W(42, 173) <= 1; flappy_W(42, 174) <= 1; flappy_W(42, 175) <= 1; flappy_W(42, 176) <= 1; flappy_W(42, 177) <= 1; flappy_W(42, 178) <= 1; flappy_W(42, 179) <= 1; flappy_W(42, 180) <= 0; flappy_W(42, 181) <= 0; flappy_W(42, 182) <= 0; flappy_W(42, 183) <= 0; flappy_W(42, 184) <= 0; flappy_W(42, 185) <= 0; flappy_W(42, 186) <= 0; flappy_W(42, 187) <= 0; flappy_W(42, 188) <= 0; flappy_W(42, 189) <= 0; flappy_W(42, 190) <= 0; flappy_W(42, 191) <= 0; flappy_W(42, 192) <= 0; flappy_W(42, 193) <= 0; flappy_W(42, 194) <= 0; flappy_W(42, 195) <= 0; flappy_W(42, 196) <= 0; flappy_W(42, 197) <= 0; flappy_W(42, 198) <= 0; flappy_W(42, 199) <= 0; flappy_W(42, 200) <= 0; flappy_W(42, 201) <= 0; flappy_W(42, 202) <= 0; flappy_W(42, 203) <= 0; flappy_W(42, 204) <= 0; flappy_W(42, 205) <= 0; flappy_W(42, 206) <= 0; flappy_W(42, 207) <= 0; flappy_W(42, 208) <= 0; flappy_W(42, 209) <= 0; flappy_W(42, 210) <= 0; flappy_W(42, 211) <= 0; flappy_W(42, 212) <= 0; flappy_W(42, 213) <= 0; flappy_W(42, 214) <= 0; flappy_W(42, 215) <= 0; flappy_W(42, 216) <= 0; flappy_W(42, 217) <= 0; flappy_W(42, 218) <= 0; flappy_W(42, 219) <= 0; flappy_W(42, 220) <= 0; flappy_W(42, 221) <= 0; flappy_W(42, 222) <= 1; flappy_W(42, 223) <= 1; flappy_W(42, 224) <= 1; flappy_W(42, 225) <= 1; flappy_W(42, 226) <= 1; flappy_W(42, 227) <= 1; flappy_W(42, 228) <= 1; flappy_W(42, 229) <= 1; flappy_W(42, 230) <= 1; flappy_W(42, 231) <= 1; flappy_W(42, 232) <= 1; flappy_W(42, 233) <= 1; flappy_W(42, 234) <= 0; flappy_W(42, 235) <= 0; flappy_W(42, 236) <= 0; flappy_W(42, 237) <= 0; flappy_W(42, 238) <= 0; flappy_W(42, 239) <= 0; flappy_W(42, 240) <= 0; flappy_W(42, 241) <= 0; flappy_W(42, 242) <= 0; flappy_W(42, 243) <= 0; flappy_W(42, 244) <= 0; flappy_W(42, 245) <= 0; flappy_W(42, 246) <= 0; flappy_W(42, 247) <= 0; flappy_W(42, 248) <= 0; flappy_W(42, 249) <= 0; flappy_W(42, 250) <= 0; flappy_W(42, 251) <= 0; flappy_W(42, 252) <= 0; flappy_W(42, 253) <= 0; flappy_W(42, 254) <= 0; flappy_W(42, 255) <= 0; flappy_W(42, 256) <= 0; flappy_W(42, 257) <= 0; flappy_W(42, 258) <= 0; flappy_W(42, 259) <= 0; flappy_W(42, 260) <= 0; flappy_W(42, 261) <= 0; flappy_W(42, 262) <= 0; flappy_W(42, 263) <= 0; flappy_W(42, 264) <= 0; flappy_W(42, 265) <= 0; flappy_W(42, 266) <= 0; flappy_W(42, 267) <= 0; flappy_W(42, 268) <= 0; flappy_W(42, 269) <= 0; flappy_W(42, 270) <= 0; flappy_W(42, 271) <= 0; flappy_W(42, 272) <= 0; flappy_W(42, 273) <= 0; flappy_W(42, 274) <= 0; flappy_W(42, 275) <= 0; flappy_W(42, 276) <= 0; flappy_W(42, 277) <= 0; flappy_W(42, 278) <= 0; flappy_W(42, 279) <= 0; flappy_W(42, 280) <= 0; flappy_W(42, 281) <= 0; flappy_W(42, 282) <= 0; flappy_W(42, 283) <= 0; flappy_W(42, 284) <= 0; flappy_W(42, 285) <= 0; flappy_W(42, 286) <= 0; flappy_W(42, 287) <= 0; flappy_W(42, 288) <= 1; flappy_W(42, 289) <= 1; flappy_W(42, 290) <= 1; flappy_W(42, 291) <= 1; flappy_W(42, 292) <= 1; flappy_W(42, 293) <= 1; flappy_W(42, 294) <= 1; flappy_W(42, 295) <= 1; flappy_W(42, 296) <= 1; flappy_W(42, 297) <= 1; flappy_W(42, 298) <= 1; flappy_W(42, 299) <= 1; flappy_W(42, 300) <= 0; flappy_W(42, 301) <= 0; flappy_W(42, 302) <= 0; flappy_W(42, 303) <= 0; flappy_W(42, 304) <= 0; flappy_W(42, 305) <= 0; flappy_W(42, 306) <= 0; flappy_W(42, 307) <= 0; flappy_W(42, 308) <= 0; flappy_W(42, 309) <= 0; flappy_W(42, 310) <= 0; flappy_W(42, 311) <= 0; flappy_W(42, 312) <= 0; flappy_W(42, 313) <= 0; flappy_W(42, 314) <= 0; flappy_W(42, 315) <= 0; flappy_W(42, 316) <= 0; flappy_W(42, 317) <= 0; flappy_W(42, 318) <= 0; flappy_W(42, 319) <= 0; flappy_W(42, 320) <= 0; flappy_W(42, 321) <= 0; flappy_W(42, 322) <= 0; flappy_W(42, 323) <= 0; flappy_W(42, 324) <= 0; flappy_W(42, 325) <= 0; flappy_W(42, 326) <= 0; flappy_W(42, 327) <= 0; flappy_W(42, 328) <= 0; flappy_W(42, 329) <= 0; flappy_W(42, 330) <= 0; flappy_W(42, 331) <= 0; flappy_W(42, 332) <= 0; flappy_W(42, 333) <= 0; flappy_W(42, 334) <= 0; flappy_W(42, 335) <= 0; flappy_W(42, 336) <= 0; flappy_W(42, 337) <= 0; flappy_W(42, 338) <= 0; flappy_W(42, 339) <= 0; flappy_W(42, 340) <= 0; flappy_W(42, 341) <= 0; flappy_W(42, 342) <= 0; flappy_W(42, 343) <= 0; flappy_W(42, 344) <= 0; flappy_W(42, 345) <= 0; flappy_W(42, 346) <= 0; flappy_W(42, 347) <= 0; flappy_W(42, 348) <= 0; flappy_W(42, 349) <= 0; flappy_W(42, 350) <= 0; flappy_W(42, 351) <= 0; flappy_W(42, 352) <= 0; flappy_W(42, 353) <= 0; flappy_W(42, 354) <= 0; flappy_W(42, 355) <= 0; flappy_W(42, 356) <= 0; flappy_W(42, 357) <= 0; flappy_W(42, 358) <= 0; flappy_W(42, 359) <= 0; flappy_W(42, 360) <= 0; flappy_W(42, 361) <= 0; flappy_W(42, 362) <= 0; flappy_W(42, 363) <= 0; flappy_W(42, 364) <= 0; flappy_W(42, 365) <= 0; flappy_W(42, 366) <= 0; flappy_W(42, 367) <= 0; flappy_W(42, 368) <= 0; flappy_W(42, 369) <= 0; flappy_W(42, 370) <= 0; flappy_W(42, 371) <= 0; flappy_W(42, 372) <= 0; flappy_W(42, 373) <= 0; flappy_W(42, 374) <= 0; flappy_W(42, 375) <= 0; flappy_W(42, 376) <= 0; flappy_W(42, 377) <= 0; flappy_W(42, 378) <= 0; flappy_W(42, 379) <= 0; flappy_W(42, 380) <= 0; flappy_W(42, 381) <= 0; flappy_W(42, 382) <= 0; flappy_W(42, 383) <= 0; flappy_W(42, 384) <= 0; flappy_W(42, 385) <= 0; flappy_W(42, 386) <= 0; flappy_W(42, 387) <= 0; flappy_W(42, 388) <= 0; flappy_W(42, 389) <= 0; flappy_W(42, 390) <= 0; flappy_W(42, 391) <= 0; flappy_W(42, 392) <= 0; flappy_W(42, 393) <= 0; flappy_W(42, 394) <= 0; flappy_W(42, 395) <= 0; flappy_W(42, 396) <= 0; flappy_W(42, 397) <= 0; flappy_W(42, 398) <= 0; flappy_W(42, 399) <= 0; flappy_W(42, 400) <= 0; flappy_W(42, 401) <= 0; flappy_W(42, 402) <= 1; flappy_W(42, 403) <= 1; flappy_W(42, 404) <= 1; flappy_W(42, 405) <= 1; flappy_W(42, 406) <= 1; flappy_W(42, 407) <= 1; flappy_W(42, 408) <= 1; flappy_W(42, 409) <= 1; flappy_W(42, 410) <= 1; flappy_W(42, 411) <= 1; flappy_W(42, 412) <= 1; flappy_W(42, 413) <= 1; flappy_W(42, 414) <= 0; flappy_W(42, 415) <= 0; flappy_W(42, 416) <= 0; flappy_W(42, 417) <= 0; flappy_W(42, 418) <= 0; flappy_W(42, 419) <= 0; flappy_W(42, 420) <= 0; flappy_W(42, 421) <= 0; flappy_W(42, 422) <= 0; flappy_W(42, 423) <= 0; flappy_W(42, 424) <= 0; flappy_W(42, 425) <= 0; flappy_W(42, 426) <= 1; flappy_W(42, 427) <= 1; flappy_W(42, 428) <= 1; flappy_W(42, 429) <= 1; flappy_W(42, 430) <= 1; flappy_W(42, 431) <= 1; flappy_W(42, 432) <= 1; flappy_W(42, 433) <= 1; flappy_W(42, 434) <= 1; flappy_W(42, 435) <= 1; flappy_W(42, 436) <= 1; flappy_W(42, 437) <= 1; flappy_W(42, 438) <= 0; flappy_W(42, 439) <= 0; flappy_W(42, 440) <= 0; flappy_W(42, 441) <= 0; flappy_W(42, 442) <= 0; flappy_W(42, 443) <= 0; flappy_W(42, 444) <= 0; flappy_W(42, 445) <= 0; flappy_W(42, 446) <= 0; flappy_W(42, 447) <= 0; flappy_W(42, 448) <= 0; flappy_W(42, 449) <= 0; flappy_W(42, 450) <= 0; flappy_W(42, 451) <= 0; flappy_W(42, 452) <= 0; flappy_W(42, 453) <= 0; flappy_W(42, 454) <= 0; flappy_W(42, 455) <= 0; flappy_W(42, 456) <= 0; flappy_W(42, 457) <= 0; flappy_W(42, 458) <= 0; flappy_W(42, 459) <= 0; flappy_W(42, 460) <= 0; flappy_W(42, 461) <= 0; flappy_W(42, 462) <= 0; flappy_W(42, 463) <= 0; flappy_W(42, 464) <= 0; flappy_W(42, 465) <= 0; flappy_W(42, 466) <= 0; flappy_W(42, 467) <= 0; flappy_W(42, 468) <= 1; flappy_W(42, 469) <= 1; flappy_W(42, 470) <= 1; flappy_W(42, 471) <= 1; flappy_W(42, 472) <= 1; flappy_W(42, 473) <= 1; flappy_W(42, 474) <= 1; flappy_W(42, 475) <= 1; flappy_W(42, 476) <= 1; flappy_W(42, 477) <= 1; flappy_W(42, 478) <= 1; flappy_W(42, 479) <= 1; flappy_W(42, 480) <= 0; flappy_W(42, 481) <= 0; flappy_W(42, 482) <= 0; flappy_W(42, 483) <= 0; flappy_W(42, 484) <= 0; flappy_W(42, 485) <= 0; flappy_W(42, 486) <= 0; flappy_W(42, 487) <= 0; flappy_W(42, 488) <= 0; flappy_W(42, 489) <= 0; flappy_W(42, 490) <= 0; flappy_W(42, 491) <= 0; flappy_W(42, 492) <= 0; flappy_W(42, 493) <= 0; flappy_W(42, 494) <= 0; flappy_W(42, 495) <= 0; flappy_W(42, 496) <= 0; flappy_W(42, 497) <= 0; flappy_W(42, 498) <= 0; flappy_W(42, 499) <= 0; flappy_W(42, 500) <= 0; flappy_W(42, 501) <= 0; flappy_W(42, 502) <= 0; flappy_W(42, 503) <= 0; flappy_W(42, 504) <= 0; flappy_W(42, 505) <= 0; flappy_W(42, 506) <= 0; flappy_W(42, 507) <= 0; flappy_W(42, 508) <= 0; flappy_W(42, 509) <= 0; flappy_W(42, 510) <= 1; flappy_W(42, 511) <= 1; flappy_W(42, 512) <= 1; flappy_W(42, 513) <= 1; flappy_W(42, 514) <= 1; flappy_W(42, 515) <= 1; flappy_W(42, 516) <= 1; flappy_W(42, 517) <= 1; flappy_W(42, 518) <= 1; flappy_W(42, 519) <= 1; flappy_W(42, 520) <= 1; flappy_W(42, 521) <= 1; flappy_W(42, 522) <= 0; flappy_W(42, 523) <= 0; flappy_W(42, 524) <= 0; flappy_W(42, 525) <= 0; flappy_W(42, 526) <= 0; flappy_W(42, 527) <= 0; flappy_W(42, 528) <= 0; flappy_W(42, 529) <= 0; flappy_W(42, 530) <= 0; flappy_W(42, 531) <= 0; flappy_W(42, 532) <= 0; flappy_W(42, 533) <= 0; flappy_W(42, 534) <= 1; flappy_W(42, 535) <= 1; flappy_W(42, 536) <= 1; flappy_W(42, 537) <= 1; flappy_W(42, 538) <= 1; flappy_W(42, 539) <= 1; flappy_W(42, 540) <= 1; flappy_W(42, 541) <= 1; flappy_W(42, 542) <= 1; flappy_W(42, 543) <= 1; flappy_W(42, 544) <= 1; flappy_W(42, 545) <= 1; flappy_W(42, 546) <= 0; flappy_W(42, 547) <= 0; flappy_W(42, 548) <= 0; flappy_W(42, 549) <= 0; flappy_W(42, 550) <= 0; flappy_W(42, 551) <= 0; flappy_W(42, 552) <= 0; flappy_W(42, 553) <= 0; flappy_W(42, 554) <= 0; flappy_W(42, 555) <= 0; flappy_W(42, 556) <= 0; flappy_W(42, 557) <= 0; flappy_W(42, 558) <= 0; flappy_W(42, 559) <= 0; flappy_W(42, 560) <= 0; flappy_W(42, 561) <= 0; flappy_W(42, 562) <= 0; flappy_W(42, 563) <= 0; flappy_W(42, 564) <= 1; flappy_W(42, 565) <= 1; flappy_W(42, 566) <= 1; flappy_W(42, 567) <= 1; flappy_W(42, 568) <= 1; flappy_W(42, 569) <= 1; flappy_W(42, 570) <= 1; flappy_W(42, 571) <= 1; flappy_W(42, 572) <= 1; flappy_W(42, 573) <= 1; flappy_W(42, 574) <= 1; flappy_W(42, 575) <= 1; flappy_W(42, 576) <= 0; flappy_W(42, 577) <= 0; flappy_W(42, 578) <= 0; flappy_W(42, 579) <= 0; flappy_W(42, 580) <= 0; flappy_W(42, 581) <= 0; flappy_W(42, 582) <= 0; flappy_W(42, 583) <= 0; flappy_W(42, 584) <= 0; flappy_W(42, 585) <= 0; flappy_W(42, 586) <= 0; flappy_W(42, 587) <= 0; flappy_W(42, 588) <= 1; flappy_W(42, 589) <= 1; flappy_W(42, 590) <= 1; flappy_W(42, 591) <= 1; flappy_W(42, 592) <= 1; flappy_W(42, 593) <= 1; 
flappy_W(43, 0) <= 0; flappy_W(43, 1) <= 0; flappy_W(43, 2) <= 0; flappy_W(43, 3) <= 0; flappy_W(43, 4) <= 0; flappy_W(43, 5) <= 0; flappy_W(43, 6) <= 1; flappy_W(43, 7) <= 1; flappy_W(43, 8) <= 1; flappy_W(43, 9) <= 1; flappy_W(43, 10) <= 1; flappy_W(43, 11) <= 1; flappy_W(43, 12) <= 1; flappy_W(43, 13) <= 1; flappy_W(43, 14) <= 1; flappy_W(43, 15) <= 1; flappy_W(43, 16) <= 1; flappy_W(43, 17) <= 1; flappy_W(43, 18) <= 0; flappy_W(43, 19) <= 0; flappy_W(43, 20) <= 0; flappy_W(43, 21) <= 0; flappy_W(43, 22) <= 0; flappy_W(43, 23) <= 0; flappy_W(43, 24) <= 0; flappy_W(43, 25) <= 0; flappy_W(43, 26) <= 0; flappy_W(43, 27) <= 0; flappy_W(43, 28) <= 0; flappy_W(43, 29) <= 0; flappy_W(43, 30) <= 0; flappy_W(43, 31) <= 0; flappy_W(43, 32) <= 0; flappy_W(43, 33) <= 0; flappy_W(43, 34) <= 0; flappy_W(43, 35) <= 0; flappy_W(43, 36) <= 0; flappy_W(43, 37) <= 0; flappy_W(43, 38) <= 0; flappy_W(43, 39) <= 0; flappy_W(43, 40) <= 0; flappy_W(43, 41) <= 0; flappy_W(43, 42) <= 0; flappy_W(43, 43) <= 0; flappy_W(43, 44) <= 0; flappy_W(43, 45) <= 0; flappy_W(43, 46) <= 0; flappy_W(43, 47) <= 0; flappy_W(43, 48) <= 0; flappy_W(43, 49) <= 0; flappy_W(43, 50) <= 0; flappy_W(43, 51) <= 0; flappy_W(43, 52) <= 0; flappy_W(43, 53) <= 0; flappy_W(43, 54) <= 0; flappy_W(43, 55) <= 0; flappy_W(43, 56) <= 0; flappy_W(43, 57) <= 0; flappy_W(43, 58) <= 0; flappy_W(43, 59) <= 0; flappy_W(43, 60) <= 1; flappy_W(43, 61) <= 1; flappy_W(43, 62) <= 1; flappy_W(43, 63) <= 1; flappy_W(43, 64) <= 1; flappy_W(43, 65) <= 1; flappy_W(43, 66) <= 1; flappy_W(43, 67) <= 1; flappy_W(43, 68) <= 1; flappy_W(43, 69) <= 1; flappy_W(43, 70) <= 1; flappy_W(43, 71) <= 1; flappy_W(43, 72) <= 0; flappy_W(43, 73) <= 0; flappy_W(43, 74) <= 0; flappy_W(43, 75) <= 0; flappy_W(43, 76) <= 0; flappy_W(43, 77) <= 0; flappy_W(43, 78) <= 0; flappy_W(43, 79) <= 0; flappy_W(43, 80) <= 0; flappy_W(43, 81) <= 0; flappy_W(43, 82) <= 0; flappy_W(43, 83) <= 0; flappy_W(43, 84) <= 0; flappy_W(43, 85) <= 0; flappy_W(43, 86) <= 0; flappy_W(43, 87) <= 0; flappy_W(43, 88) <= 0; flappy_W(43, 89) <= 0; flappy_W(43, 90) <= 1; flappy_W(43, 91) <= 1; flappy_W(43, 92) <= 1; flappy_W(43, 93) <= 1; flappy_W(43, 94) <= 1; flappy_W(43, 95) <= 1; flappy_W(43, 96) <= 0; flappy_W(43, 97) <= 0; flappy_W(43, 98) <= 0; flappy_W(43, 99) <= 0; flappy_W(43, 100) <= 0; flappy_W(43, 101) <= 0; flappy_W(43, 102) <= 0; flappy_W(43, 103) <= 0; flappy_W(43, 104) <= 0; flappy_W(43, 105) <= 0; flappy_W(43, 106) <= 0; flappy_W(43, 107) <= 0; flappy_W(43, 108) <= 1; flappy_W(43, 109) <= 1; flappy_W(43, 110) <= 1; flappy_W(43, 111) <= 1; flappy_W(43, 112) <= 1; flappy_W(43, 113) <= 1; flappy_W(43, 114) <= 1; flappy_W(43, 115) <= 1; flappy_W(43, 116) <= 1; flappy_W(43, 117) <= 1; flappy_W(43, 118) <= 1; flappy_W(43, 119) <= 1; flappy_W(43, 120) <= 0; flappy_W(43, 121) <= 0; flappy_W(43, 122) <= 0; flappy_W(43, 123) <= 0; flappy_W(43, 124) <= 0; flappy_W(43, 125) <= 0; flappy_W(43, 126) <= 0; flappy_W(43, 127) <= 0; flappy_W(43, 128) <= 0; flappy_W(43, 129) <= 0; flappy_W(43, 130) <= 0; flappy_W(43, 131) <= 0; flappy_W(43, 132) <= 0; flappy_W(43, 133) <= 0; flappy_W(43, 134) <= 0; flappy_W(43, 135) <= 0; flappy_W(43, 136) <= 0; flappy_W(43, 137) <= 0; flappy_W(43, 138) <= 1; flappy_W(43, 139) <= 1; flappy_W(43, 140) <= 1; flappy_W(43, 141) <= 1; flappy_W(43, 142) <= 1; flappy_W(43, 143) <= 1; flappy_W(43, 144) <= 1; flappy_W(43, 145) <= 1; flappy_W(43, 146) <= 1; flappy_W(43, 147) <= 1; flappy_W(43, 148) <= 1; flappy_W(43, 149) <= 1; flappy_W(43, 150) <= 0; flappy_W(43, 151) <= 0; flappy_W(43, 152) <= 0; flappy_W(43, 153) <= 0; flappy_W(43, 154) <= 0; flappy_W(43, 155) <= 0; flappy_W(43, 156) <= 0; flappy_W(43, 157) <= 0; flappy_W(43, 158) <= 0; flappy_W(43, 159) <= 0; flappy_W(43, 160) <= 0; flappy_W(43, 161) <= 0; flappy_W(43, 162) <= 0; flappy_W(43, 163) <= 0; flappy_W(43, 164) <= 0; flappy_W(43, 165) <= 0; flappy_W(43, 166) <= 0; flappy_W(43, 167) <= 0; flappy_W(43, 168) <= 1; flappy_W(43, 169) <= 1; flappy_W(43, 170) <= 1; flappy_W(43, 171) <= 1; flappy_W(43, 172) <= 1; flappy_W(43, 173) <= 1; flappy_W(43, 174) <= 1; flappy_W(43, 175) <= 1; flappy_W(43, 176) <= 1; flappy_W(43, 177) <= 1; flappy_W(43, 178) <= 1; flappy_W(43, 179) <= 1; flappy_W(43, 180) <= 0; flappy_W(43, 181) <= 0; flappy_W(43, 182) <= 0; flappy_W(43, 183) <= 0; flappy_W(43, 184) <= 0; flappy_W(43, 185) <= 0; flappy_W(43, 186) <= 0; flappy_W(43, 187) <= 0; flappy_W(43, 188) <= 0; flappy_W(43, 189) <= 0; flappy_W(43, 190) <= 0; flappy_W(43, 191) <= 0; flappy_W(43, 192) <= 0; flappy_W(43, 193) <= 0; flappy_W(43, 194) <= 0; flappy_W(43, 195) <= 0; flappy_W(43, 196) <= 0; flappy_W(43, 197) <= 0; flappy_W(43, 198) <= 0; flappy_W(43, 199) <= 0; flappy_W(43, 200) <= 0; flappy_W(43, 201) <= 0; flappy_W(43, 202) <= 0; flappy_W(43, 203) <= 0; flappy_W(43, 204) <= 0; flappy_W(43, 205) <= 0; flappy_W(43, 206) <= 0; flappy_W(43, 207) <= 0; flappy_W(43, 208) <= 0; flappy_W(43, 209) <= 0; flappy_W(43, 210) <= 0; flappy_W(43, 211) <= 0; flappy_W(43, 212) <= 0; flappy_W(43, 213) <= 0; flappy_W(43, 214) <= 0; flappy_W(43, 215) <= 0; flappy_W(43, 216) <= 0; flappy_W(43, 217) <= 0; flappy_W(43, 218) <= 0; flappy_W(43, 219) <= 0; flappy_W(43, 220) <= 0; flappy_W(43, 221) <= 0; flappy_W(43, 222) <= 1; flappy_W(43, 223) <= 1; flappy_W(43, 224) <= 1; flappy_W(43, 225) <= 1; flappy_W(43, 226) <= 1; flappy_W(43, 227) <= 1; flappy_W(43, 228) <= 1; flappy_W(43, 229) <= 1; flappy_W(43, 230) <= 1; flappy_W(43, 231) <= 1; flappy_W(43, 232) <= 1; flappy_W(43, 233) <= 1; flappy_W(43, 234) <= 0; flappy_W(43, 235) <= 0; flappy_W(43, 236) <= 0; flappy_W(43, 237) <= 0; flappy_W(43, 238) <= 0; flappy_W(43, 239) <= 0; flappy_W(43, 240) <= 0; flappy_W(43, 241) <= 0; flappy_W(43, 242) <= 0; flappy_W(43, 243) <= 0; flappy_W(43, 244) <= 0; flappy_W(43, 245) <= 0; flappy_W(43, 246) <= 0; flappy_W(43, 247) <= 0; flappy_W(43, 248) <= 0; flappy_W(43, 249) <= 0; flappy_W(43, 250) <= 0; flappy_W(43, 251) <= 0; flappy_W(43, 252) <= 0; flappy_W(43, 253) <= 0; flappy_W(43, 254) <= 0; flappy_W(43, 255) <= 0; flappy_W(43, 256) <= 0; flappy_W(43, 257) <= 0; flappy_W(43, 258) <= 0; flappy_W(43, 259) <= 0; flappy_W(43, 260) <= 0; flappy_W(43, 261) <= 0; flappy_W(43, 262) <= 0; flappy_W(43, 263) <= 0; flappy_W(43, 264) <= 0; flappy_W(43, 265) <= 0; flappy_W(43, 266) <= 0; flappy_W(43, 267) <= 0; flappy_W(43, 268) <= 0; flappy_W(43, 269) <= 0; flappy_W(43, 270) <= 0; flappy_W(43, 271) <= 0; flappy_W(43, 272) <= 0; flappy_W(43, 273) <= 0; flappy_W(43, 274) <= 0; flappy_W(43, 275) <= 0; flappy_W(43, 276) <= 0; flappy_W(43, 277) <= 0; flappy_W(43, 278) <= 0; flappy_W(43, 279) <= 0; flappy_W(43, 280) <= 0; flappy_W(43, 281) <= 0; flappy_W(43, 282) <= 0; flappy_W(43, 283) <= 0; flappy_W(43, 284) <= 0; flappy_W(43, 285) <= 0; flappy_W(43, 286) <= 0; flappy_W(43, 287) <= 0; flappy_W(43, 288) <= 1; flappy_W(43, 289) <= 1; flappy_W(43, 290) <= 1; flappy_W(43, 291) <= 1; flappy_W(43, 292) <= 1; flappy_W(43, 293) <= 1; flappy_W(43, 294) <= 1; flappy_W(43, 295) <= 1; flappy_W(43, 296) <= 1; flappy_W(43, 297) <= 1; flappy_W(43, 298) <= 1; flappy_W(43, 299) <= 1; flappy_W(43, 300) <= 0; flappy_W(43, 301) <= 0; flappy_W(43, 302) <= 0; flappy_W(43, 303) <= 0; flappy_W(43, 304) <= 0; flappy_W(43, 305) <= 0; flappy_W(43, 306) <= 0; flappy_W(43, 307) <= 0; flappy_W(43, 308) <= 0; flappy_W(43, 309) <= 0; flappy_W(43, 310) <= 0; flappy_W(43, 311) <= 0; flappy_W(43, 312) <= 0; flappy_W(43, 313) <= 0; flappy_W(43, 314) <= 0; flappy_W(43, 315) <= 0; flappy_W(43, 316) <= 0; flappy_W(43, 317) <= 0; flappy_W(43, 318) <= 0; flappy_W(43, 319) <= 0; flappy_W(43, 320) <= 0; flappy_W(43, 321) <= 0; flappy_W(43, 322) <= 0; flappy_W(43, 323) <= 0; flappy_W(43, 324) <= 0; flappy_W(43, 325) <= 0; flappy_W(43, 326) <= 0; flappy_W(43, 327) <= 0; flappy_W(43, 328) <= 0; flappy_W(43, 329) <= 0; flappy_W(43, 330) <= 0; flappy_W(43, 331) <= 0; flappy_W(43, 332) <= 0; flappy_W(43, 333) <= 0; flappy_W(43, 334) <= 0; flappy_W(43, 335) <= 0; flappy_W(43, 336) <= 0; flappy_W(43, 337) <= 0; flappy_W(43, 338) <= 0; flappy_W(43, 339) <= 0; flappy_W(43, 340) <= 0; flappy_W(43, 341) <= 0; flappy_W(43, 342) <= 0; flappy_W(43, 343) <= 0; flappy_W(43, 344) <= 0; flappy_W(43, 345) <= 0; flappy_W(43, 346) <= 0; flappy_W(43, 347) <= 0; flappy_W(43, 348) <= 0; flappy_W(43, 349) <= 0; flappy_W(43, 350) <= 0; flappy_W(43, 351) <= 0; flappy_W(43, 352) <= 0; flappy_W(43, 353) <= 0; flappy_W(43, 354) <= 0; flappy_W(43, 355) <= 0; flappy_W(43, 356) <= 0; flappy_W(43, 357) <= 0; flappy_W(43, 358) <= 0; flappy_W(43, 359) <= 0; flappy_W(43, 360) <= 0; flappy_W(43, 361) <= 0; flappy_W(43, 362) <= 0; flappy_W(43, 363) <= 0; flappy_W(43, 364) <= 0; flappy_W(43, 365) <= 0; flappy_W(43, 366) <= 0; flappy_W(43, 367) <= 0; flappy_W(43, 368) <= 0; flappy_W(43, 369) <= 0; flappy_W(43, 370) <= 0; flappy_W(43, 371) <= 0; flappy_W(43, 372) <= 0; flappy_W(43, 373) <= 0; flappy_W(43, 374) <= 0; flappy_W(43, 375) <= 0; flappy_W(43, 376) <= 0; flappy_W(43, 377) <= 0; flappy_W(43, 378) <= 0; flappy_W(43, 379) <= 0; flappy_W(43, 380) <= 0; flappy_W(43, 381) <= 0; flappy_W(43, 382) <= 0; flappy_W(43, 383) <= 0; flappy_W(43, 384) <= 0; flappy_W(43, 385) <= 0; flappy_W(43, 386) <= 0; flappy_W(43, 387) <= 0; flappy_W(43, 388) <= 0; flappy_W(43, 389) <= 0; flappy_W(43, 390) <= 0; flappy_W(43, 391) <= 0; flappy_W(43, 392) <= 0; flappy_W(43, 393) <= 0; flappy_W(43, 394) <= 0; flappy_W(43, 395) <= 0; flappy_W(43, 396) <= 0; flappy_W(43, 397) <= 0; flappy_W(43, 398) <= 0; flappy_W(43, 399) <= 0; flappy_W(43, 400) <= 0; flappy_W(43, 401) <= 0; flappy_W(43, 402) <= 1; flappy_W(43, 403) <= 1; flappy_W(43, 404) <= 1; flappy_W(43, 405) <= 1; flappy_W(43, 406) <= 1; flappy_W(43, 407) <= 1; flappy_W(43, 408) <= 1; flappy_W(43, 409) <= 1; flappy_W(43, 410) <= 1; flappy_W(43, 411) <= 1; flappy_W(43, 412) <= 1; flappy_W(43, 413) <= 1; flappy_W(43, 414) <= 0; flappy_W(43, 415) <= 0; flappy_W(43, 416) <= 0; flappy_W(43, 417) <= 0; flappy_W(43, 418) <= 0; flappy_W(43, 419) <= 0; flappy_W(43, 420) <= 0; flappy_W(43, 421) <= 0; flappy_W(43, 422) <= 0; flappy_W(43, 423) <= 0; flappy_W(43, 424) <= 0; flappy_W(43, 425) <= 0; flappy_W(43, 426) <= 1; flappy_W(43, 427) <= 1; flappy_W(43, 428) <= 1; flappy_W(43, 429) <= 1; flappy_W(43, 430) <= 1; flappy_W(43, 431) <= 1; flappy_W(43, 432) <= 1; flappy_W(43, 433) <= 1; flappy_W(43, 434) <= 1; flappy_W(43, 435) <= 1; flappy_W(43, 436) <= 1; flappy_W(43, 437) <= 1; flappy_W(43, 438) <= 0; flappy_W(43, 439) <= 0; flappy_W(43, 440) <= 0; flappy_W(43, 441) <= 0; flappy_W(43, 442) <= 0; flappy_W(43, 443) <= 0; flappy_W(43, 444) <= 0; flappy_W(43, 445) <= 0; flappy_W(43, 446) <= 0; flappy_W(43, 447) <= 0; flappy_W(43, 448) <= 0; flappy_W(43, 449) <= 0; flappy_W(43, 450) <= 0; flappy_W(43, 451) <= 0; flappy_W(43, 452) <= 0; flappy_W(43, 453) <= 0; flappy_W(43, 454) <= 0; flappy_W(43, 455) <= 0; flappy_W(43, 456) <= 0; flappy_W(43, 457) <= 0; flappy_W(43, 458) <= 0; flappy_W(43, 459) <= 0; flappy_W(43, 460) <= 0; flappy_W(43, 461) <= 0; flappy_W(43, 462) <= 0; flappy_W(43, 463) <= 0; flappy_W(43, 464) <= 0; flappy_W(43, 465) <= 0; flappy_W(43, 466) <= 0; flappy_W(43, 467) <= 0; flappy_W(43, 468) <= 1; flappy_W(43, 469) <= 1; flappy_W(43, 470) <= 1; flappy_W(43, 471) <= 1; flappy_W(43, 472) <= 1; flappy_W(43, 473) <= 1; flappy_W(43, 474) <= 1; flappy_W(43, 475) <= 1; flappy_W(43, 476) <= 1; flappy_W(43, 477) <= 1; flappy_W(43, 478) <= 1; flappy_W(43, 479) <= 1; flappy_W(43, 480) <= 0; flappy_W(43, 481) <= 0; flappy_W(43, 482) <= 0; flappy_W(43, 483) <= 0; flappy_W(43, 484) <= 0; flappy_W(43, 485) <= 0; flappy_W(43, 486) <= 0; flappy_W(43, 487) <= 0; flappy_W(43, 488) <= 0; flappy_W(43, 489) <= 0; flappy_W(43, 490) <= 0; flappy_W(43, 491) <= 0; flappy_W(43, 492) <= 0; flappy_W(43, 493) <= 0; flappy_W(43, 494) <= 0; flappy_W(43, 495) <= 0; flappy_W(43, 496) <= 0; flappy_W(43, 497) <= 0; flappy_W(43, 498) <= 0; flappy_W(43, 499) <= 0; flappy_W(43, 500) <= 0; flappy_W(43, 501) <= 0; flappy_W(43, 502) <= 0; flappy_W(43, 503) <= 0; flappy_W(43, 504) <= 0; flappy_W(43, 505) <= 0; flappy_W(43, 506) <= 0; flappy_W(43, 507) <= 0; flappy_W(43, 508) <= 0; flappy_W(43, 509) <= 0; flappy_W(43, 510) <= 1; flappy_W(43, 511) <= 1; flappy_W(43, 512) <= 1; flappy_W(43, 513) <= 1; flappy_W(43, 514) <= 1; flappy_W(43, 515) <= 1; flappy_W(43, 516) <= 1; flappy_W(43, 517) <= 1; flappy_W(43, 518) <= 1; flappy_W(43, 519) <= 1; flappy_W(43, 520) <= 1; flappy_W(43, 521) <= 1; flappy_W(43, 522) <= 0; flappy_W(43, 523) <= 0; flappy_W(43, 524) <= 0; flappy_W(43, 525) <= 0; flappy_W(43, 526) <= 0; flappy_W(43, 527) <= 0; flappy_W(43, 528) <= 0; flappy_W(43, 529) <= 0; flappy_W(43, 530) <= 0; flappy_W(43, 531) <= 0; flappy_W(43, 532) <= 0; flappy_W(43, 533) <= 0; flappy_W(43, 534) <= 1; flappy_W(43, 535) <= 1; flappy_W(43, 536) <= 1; flappy_W(43, 537) <= 1; flappy_W(43, 538) <= 1; flappy_W(43, 539) <= 1; flappy_W(43, 540) <= 1; flappy_W(43, 541) <= 1; flappy_W(43, 542) <= 1; flappy_W(43, 543) <= 1; flappy_W(43, 544) <= 1; flappy_W(43, 545) <= 1; flappy_W(43, 546) <= 0; flappy_W(43, 547) <= 0; flappy_W(43, 548) <= 0; flappy_W(43, 549) <= 0; flappy_W(43, 550) <= 0; flappy_W(43, 551) <= 0; flappy_W(43, 552) <= 0; flappy_W(43, 553) <= 0; flappy_W(43, 554) <= 0; flappy_W(43, 555) <= 0; flappy_W(43, 556) <= 0; flappy_W(43, 557) <= 0; flappy_W(43, 558) <= 0; flappy_W(43, 559) <= 0; flappy_W(43, 560) <= 0; flappy_W(43, 561) <= 0; flappy_W(43, 562) <= 0; flappy_W(43, 563) <= 0; flappy_W(43, 564) <= 1; flappy_W(43, 565) <= 1; flappy_W(43, 566) <= 1; flappy_W(43, 567) <= 1; flappy_W(43, 568) <= 1; flappy_W(43, 569) <= 1; flappy_W(43, 570) <= 1; flappy_W(43, 571) <= 1; flappy_W(43, 572) <= 1; flappy_W(43, 573) <= 1; flappy_W(43, 574) <= 1; flappy_W(43, 575) <= 1; flappy_W(43, 576) <= 0; flappy_W(43, 577) <= 0; flappy_W(43, 578) <= 0; flappy_W(43, 579) <= 0; flappy_W(43, 580) <= 0; flappy_W(43, 581) <= 0; flappy_W(43, 582) <= 0; flappy_W(43, 583) <= 0; flappy_W(43, 584) <= 0; flappy_W(43, 585) <= 0; flappy_W(43, 586) <= 0; flappy_W(43, 587) <= 0; flappy_W(43, 588) <= 1; flappy_W(43, 589) <= 1; flappy_W(43, 590) <= 1; flappy_W(43, 591) <= 1; flappy_W(43, 592) <= 1; flappy_W(43, 593) <= 1; 
flappy_W(44, 0) <= 0; flappy_W(44, 1) <= 0; flappy_W(44, 2) <= 0; flappy_W(44, 3) <= 0; flappy_W(44, 4) <= 0; flappy_W(44, 5) <= 0; flappy_W(44, 6) <= 1; flappy_W(44, 7) <= 1; flappy_W(44, 8) <= 1; flappy_W(44, 9) <= 1; flappy_W(44, 10) <= 1; flappy_W(44, 11) <= 1; flappy_W(44, 12) <= 1; flappy_W(44, 13) <= 1; flappy_W(44, 14) <= 1; flappy_W(44, 15) <= 1; flappy_W(44, 16) <= 1; flappy_W(44, 17) <= 1; flappy_W(44, 18) <= 0; flappy_W(44, 19) <= 0; flappy_W(44, 20) <= 0; flappy_W(44, 21) <= 0; flappy_W(44, 22) <= 0; flappy_W(44, 23) <= 0; flappy_W(44, 24) <= 0; flappy_W(44, 25) <= 0; flappy_W(44, 26) <= 0; flappy_W(44, 27) <= 0; flappy_W(44, 28) <= 0; flappy_W(44, 29) <= 0; flappy_W(44, 30) <= 0; flappy_W(44, 31) <= 0; flappy_W(44, 32) <= 0; flappy_W(44, 33) <= 0; flappy_W(44, 34) <= 0; flappy_W(44, 35) <= 0; flappy_W(44, 36) <= 0; flappy_W(44, 37) <= 0; flappy_W(44, 38) <= 0; flappy_W(44, 39) <= 0; flappy_W(44, 40) <= 0; flappy_W(44, 41) <= 0; flappy_W(44, 42) <= 0; flappy_W(44, 43) <= 0; flappy_W(44, 44) <= 0; flappy_W(44, 45) <= 0; flappy_W(44, 46) <= 0; flappy_W(44, 47) <= 0; flappy_W(44, 48) <= 0; flappy_W(44, 49) <= 0; flappy_W(44, 50) <= 0; flappy_W(44, 51) <= 0; flappy_W(44, 52) <= 0; flappy_W(44, 53) <= 0; flappy_W(44, 54) <= 0; flappy_W(44, 55) <= 0; flappy_W(44, 56) <= 0; flappy_W(44, 57) <= 0; flappy_W(44, 58) <= 0; flappy_W(44, 59) <= 0; flappy_W(44, 60) <= 1; flappy_W(44, 61) <= 1; flappy_W(44, 62) <= 1; flappy_W(44, 63) <= 1; flappy_W(44, 64) <= 1; flappy_W(44, 65) <= 1; flappy_W(44, 66) <= 1; flappy_W(44, 67) <= 1; flappy_W(44, 68) <= 1; flappy_W(44, 69) <= 1; flappy_W(44, 70) <= 1; flappy_W(44, 71) <= 1; flappy_W(44, 72) <= 0; flappy_W(44, 73) <= 0; flappy_W(44, 74) <= 0; flappy_W(44, 75) <= 0; flappy_W(44, 76) <= 0; flappy_W(44, 77) <= 0; flappy_W(44, 78) <= 0; flappy_W(44, 79) <= 0; flappy_W(44, 80) <= 0; flappy_W(44, 81) <= 0; flappy_W(44, 82) <= 0; flappy_W(44, 83) <= 0; flappy_W(44, 84) <= 0; flappy_W(44, 85) <= 0; flappy_W(44, 86) <= 0; flappy_W(44, 87) <= 0; flappy_W(44, 88) <= 0; flappy_W(44, 89) <= 0; flappy_W(44, 90) <= 1; flappy_W(44, 91) <= 1; flappy_W(44, 92) <= 1; flappy_W(44, 93) <= 1; flappy_W(44, 94) <= 1; flappy_W(44, 95) <= 1; flappy_W(44, 96) <= 0; flappy_W(44, 97) <= 0; flappy_W(44, 98) <= 0; flappy_W(44, 99) <= 0; flappy_W(44, 100) <= 0; flappy_W(44, 101) <= 0; flappy_W(44, 102) <= 0; flappy_W(44, 103) <= 0; flappy_W(44, 104) <= 0; flappy_W(44, 105) <= 0; flappy_W(44, 106) <= 0; flappy_W(44, 107) <= 0; flappy_W(44, 108) <= 1; flappy_W(44, 109) <= 1; flappy_W(44, 110) <= 1; flappy_W(44, 111) <= 1; flappy_W(44, 112) <= 1; flappy_W(44, 113) <= 1; flappy_W(44, 114) <= 1; flappy_W(44, 115) <= 1; flappy_W(44, 116) <= 1; flappy_W(44, 117) <= 1; flappy_W(44, 118) <= 1; flappy_W(44, 119) <= 1; flappy_W(44, 120) <= 0; flappy_W(44, 121) <= 0; flappy_W(44, 122) <= 0; flappy_W(44, 123) <= 0; flappy_W(44, 124) <= 0; flappy_W(44, 125) <= 0; flappy_W(44, 126) <= 0; flappy_W(44, 127) <= 0; flappy_W(44, 128) <= 0; flappy_W(44, 129) <= 0; flappy_W(44, 130) <= 0; flappy_W(44, 131) <= 0; flappy_W(44, 132) <= 0; flappy_W(44, 133) <= 0; flappy_W(44, 134) <= 0; flappy_W(44, 135) <= 0; flappy_W(44, 136) <= 0; flappy_W(44, 137) <= 0; flappy_W(44, 138) <= 1; flappy_W(44, 139) <= 1; flappy_W(44, 140) <= 1; flappy_W(44, 141) <= 1; flappy_W(44, 142) <= 1; flappy_W(44, 143) <= 1; flappy_W(44, 144) <= 1; flappy_W(44, 145) <= 1; flappy_W(44, 146) <= 1; flappy_W(44, 147) <= 1; flappy_W(44, 148) <= 1; flappy_W(44, 149) <= 1; flappy_W(44, 150) <= 0; flappy_W(44, 151) <= 0; flappy_W(44, 152) <= 0; flappy_W(44, 153) <= 0; flappy_W(44, 154) <= 0; flappy_W(44, 155) <= 0; flappy_W(44, 156) <= 0; flappy_W(44, 157) <= 0; flappy_W(44, 158) <= 0; flappy_W(44, 159) <= 0; flappy_W(44, 160) <= 0; flappy_W(44, 161) <= 0; flappy_W(44, 162) <= 0; flappy_W(44, 163) <= 0; flappy_W(44, 164) <= 0; flappy_W(44, 165) <= 0; flappy_W(44, 166) <= 0; flappy_W(44, 167) <= 0; flappy_W(44, 168) <= 1; flappy_W(44, 169) <= 1; flappy_W(44, 170) <= 1; flappy_W(44, 171) <= 1; flappy_W(44, 172) <= 1; flappy_W(44, 173) <= 1; flappy_W(44, 174) <= 1; flappy_W(44, 175) <= 1; flappy_W(44, 176) <= 1; flappy_W(44, 177) <= 1; flappy_W(44, 178) <= 1; flappy_W(44, 179) <= 1; flappy_W(44, 180) <= 0; flappy_W(44, 181) <= 0; flappy_W(44, 182) <= 0; flappy_W(44, 183) <= 0; flappy_W(44, 184) <= 0; flappy_W(44, 185) <= 0; flappy_W(44, 186) <= 0; flappy_W(44, 187) <= 0; flappy_W(44, 188) <= 0; flappy_W(44, 189) <= 0; flappy_W(44, 190) <= 0; flappy_W(44, 191) <= 0; flappy_W(44, 192) <= 0; flappy_W(44, 193) <= 0; flappy_W(44, 194) <= 0; flappy_W(44, 195) <= 0; flappy_W(44, 196) <= 0; flappy_W(44, 197) <= 0; flappy_W(44, 198) <= 0; flappy_W(44, 199) <= 0; flappy_W(44, 200) <= 0; flappy_W(44, 201) <= 0; flappy_W(44, 202) <= 0; flappy_W(44, 203) <= 0; flappy_W(44, 204) <= 0; flappy_W(44, 205) <= 0; flappy_W(44, 206) <= 0; flappy_W(44, 207) <= 0; flappy_W(44, 208) <= 0; flappy_W(44, 209) <= 0; flappy_W(44, 210) <= 0; flappy_W(44, 211) <= 0; flappy_W(44, 212) <= 0; flappy_W(44, 213) <= 0; flappy_W(44, 214) <= 0; flappy_W(44, 215) <= 0; flappy_W(44, 216) <= 0; flappy_W(44, 217) <= 0; flappy_W(44, 218) <= 0; flappy_W(44, 219) <= 0; flappy_W(44, 220) <= 0; flappy_W(44, 221) <= 0; flappy_W(44, 222) <= 1; flappy_W(44, 223) <= 1; flappy_W(44, 224) <= 1; flappy_W(44, 225) <= 1; flappy_W(44, 226) <= 1; flappy_W(44, 227) <= 1; flappy_W(44, 228) <= 1; flappy_W(44, 229) <= 1; flappy_W(44, 230) <= 1; flappy_W(44, 231) <= 1; flappy_W(44, 232) <= 1; flappy_W(44, 233) <= 1; flappy_W(44, 234) <= 0; flappy_W(44, 235) <= 0; flappy_W(44, 236) <= 0; flappy_W(44, 237) <= 0; flappy_W(44, 238) <= 0; flappy_W(44, 239) <= 0; flappy_W(44, 240) <= 0; flappy_W(44, 241) <= 0; flappy_W(44, 242) <= 0; flappy_W(44, 243) <= 0; flappy_W(44, 244) <= 0; flappy_W(44, 245) <= 0; flappy_W(44, 246) <= 0; flappy_W(44, 247) <= 0; flappy_W(44, 248) <= 0; flappy_W(44, 249) <= 0; flappy_W(44, 250) <= 0; flappy_W(44, 251) <= 0; flappy_W(44, 252) <= 0; flappy_W(44, 253) <= 0; flappy_W(44, 254) <= 0; flappy_W(44, 255) <= 0; flappy_W(44, 256) <= 0; flappy_W(44, 257) <= 0; flappy_W(44, 258) <= 0; flappy_W(44, 259) <= 0; flappy_W(44, 260) <= 0; flappy_W(44, 261) <= 0; flappy_W(44, 262) <= 0; flappy_W(44, 263) <= 0; flappy_W(44, 264) <= 0; flappy_W(44, 265) <= 0; flappy_W(44, 266) <= 0; flappy_W(44, 267) <= 0; flappy_W(44, 268) <= 0; flappy_W(44, 269) <= 0; flappy_W(44, 270) <= 0; flappy_W(44, 271) <= 0; flappy_W(44, 272) <= 0; flappy_W(44, 273) <= 0; flappy_W(44, 274) <= 0; flappy_W(44, 275) <= 0; flappy_W(44, 276) <= 0; flappy_W(44, 277) <= 0; flappy_W(44, 278) <= 0; flappy_W(44, 279) <= 0; flappy_W(44, 280) <= 0; flappy_W(44, 281) <= 0; flappy_W(44, 282) <= 0; flappy_W(44, 283) <= 0; flappy_W(44, 284) <= 0; flappy_W(44, 285) <= 0; flappy_W(44, 286) <= 0; flappy_W(44, 287) <= 0; flappy_W(44, 288) <= 1; flappy_W(44, 289) <= 1; flappy_W(44, 290) <= 1; flappy_W(44, 291) <= 1; flappy_W(44, 292) <= 1; flappy_W(44, 293) <= 1; flappy_W(44, 294) <= 1; flappy_W(44, 295) <= 1; flappy_W(44, 296) <= 1; flappy_W(44, 297) <= 1; flappy_W(44, 298) <= 1; flappy_W(44, 299) <= 1; flappy_W(44, 300) <= 0; flappy_W(44, 301) <= 0; flappy_W(44, 302) <= 0; flappy_W(44, 303) <= 0; flappy_W(44, 304) <= 0; flappy_W(44, 305) <= 0; flappy_W(44, 306) <= 0; flappy_W(44, 307) <= 0; flappy_W(44, 308) <= 0; flappy_W(44, 309) <= 0; flappy_W(44, 310) <= 0; flappy_W(44, 311) <= 0; flappy_W(44, 312) <= 0; flappy_W(44, 313) <= 0; flappy_W(44, 314) <= 0; flappy_W(44, 315) <= 0; flappy_W(44, 316) <= 0; flappy_W(44, 317) <= 0; flappy_W(44, 318) <= 0; flappy_W(44, 319) <= 0; flappy_W(44, 320) <= 0; flappy_W(44, 321) <= 0; flappy_W(44, 322) <= 0; flappy_W(44, 323) <= 0; flappy_W(44, 324) <= 0; flappy_W(44, 325) <= 0; flappy_W(44, 326) <= 0; flappy_W(44, 327) <= 0; flappy_W(44, 328) <= 0; flappy_W(44, 329) <= 0; flappy_W(44, 330) <= 0; flappy_W(44, 331) <= 0; flappy_W(44, 332) <= 0; flappy_W(44, 333) <= 0; flappy_W(44, 334) <= 0; flappy_W(44, 335) <= 0; flappy_W(44, 336) <= 0; flappy_W(44, 337) <= 0; flappy_W(44, 338) <= 0; flappy_W(44, 339) <= 0; flappy_W(44, 340) <= 0; flappy_W(44, 341) <= 0; flappy_W(44, 342) <= 0; flappy_W(44, 343) <= 0; flappy_W(44, 344) <= 0; flappy_W(44, 345) <= 0; flappy_W(44, 346) <= 0; flappy_W(44, 347) <= 0; flappy_W(44, 348) <= 0; flappy_W(44, 349) <= 0; flappy_W(44, 350) <= 0; flappy_W(44, 351) <= 0; flappy_W(44, 352) <= 0; flappy_W(44, 353) <= 0; flappy_W(44, 354) <= 0; flappy_W(44, 355) <= 0; flappy_W(44, 356) <= 0; flappy_W(44, 357) <= 0; flappy_W(44, 358) <= 0; flappy_W(44, 359) <= 0; flappy_W(44, 360) <= 0; flappy_W(44, 361) <= 0; flappy_W(44, 362) <= 0; flappy_W(44, 363) <= 0; flappy_W(44, 364) <= 0; flappy_W(44, 365) <= 0; flappy_W(44, 366) <= 0; flappy_W(44, 367) <= 0; flappy_W(44, 368) <= 0; flappy_W(44, 369) <= 0; flappy_W(44, 370) <= 0; flappy_W(44, 371) <= 0; flappy_W(44, 372) <= 0; flappy_W(44, 373) <= 0; flappy_W(44, 374) <= 0; flappy_W(44, 375) <= 0; flappy_W(44, 376) <= 0; flappy_W(44, 377) <= 0; flappy_W(44, 378) <= 0; flappy_W(44, 379) <= 0; flappy_W(44, 380) <= 0; flappy_W(44, 381) <= 0; flappy_W(44, 382) <= 0; flappy_W(44, 383) <= 0; flappy_W(44, 384) <= 0; flappy_W(44, 385) <= 0; flappy_W(44, 386) <= 0; flappy_W(44, 387) <= 0; flappy_W(44, 388) <= 0; flappy_W(44, 389) <= 0; flappy_W(44, 390) <= 0; flappy_W(44, 391) <= 0; flappy_W(44, 392) <= 0; flappy_W(44, 393) <= 0; flappy_W(44, 394) <= 0; flappy_W(44, 395) <= 0; flappy_W(44, 396) <= 0; flappy_W(44, 397) <= 0; flappy_W(44, 398) <= 0; flappy_W(44, 399) <= 0; flappy_W(44, 400) <= 0; flappy_W(44, 401) <= 0; flappy_W(44, 402) <= 1; flappy_W(44, 403) <= 1; flappy_W(44, 404) <= 1; flappy_W(44, 405) <= 1; flappy_W(44, 406) <= 1; flappy_W(44, 407) <= 1; flappy_W(44, 408) <= 1; flappy_W(44, 409) <= 1; flappy_W(44, 410) <= 1; flappy_W(44, 411) <= 1; flappy_W(44, 412) <= 1; flappy_W(44, 413) <= 1; flappy_W(44, 414) <= 0; flappy_W(44, 415) <= 0; flappy_W(44, 416) <= 0; flappy_W(44, 417) <= 0; flappy_W(44, 418) <= 0; flappy_W(44, 419) <= 0; flappy_W(44, 420) <= 0; flappy_W(44, 421) <= 0; flappy_W(44, 422) <= 0; flappy_W(44, 423) <= 0; flappy_W(44, 424) <= 0; flappy_W(44, 425) <= 0; flappy_W(44, 426) <= 1; flappy_W(44, 427) <= 1; flappy_W(44, 428) <= 1; flappy_W(44, 429) <= 1; flappy_W(44, 430) <= 1; flappy_W(44, 431) <= 1; flappy_W(44, 432) <= 1; flappy_W(44, 433) <= 1; flappy_W(44, 434) <= 1; flappy_W(44, 435) <= 1; flappy_W(44, 436) <= 1; flappy_W(44, 437) <= 1; flappy_W(44, 438) <= 0; flappy_W(44, 439) <= 0; flappy_W(44, 440) <= 0; flappy_W(44, 441) <= 0; flappy_W(44, 442) <= 0; flappy_W(44, 443) <= 0; flappy_W(44, 444) <= 0; flappy_W(44, 445) <= 0; flappy_W(44, 446) <= 0; flappy_W(44, 447) <= 0; flappy_W(44, 448) <= 0; flappy_W(44, 449) <= 0; flappy_W(44, 450) <= 0; flappy_W(44, 451) <= 0; flappy_W(44, 452) <= 0; flappy_W(44, 453) <= 0; flappy_W(44, 454) <= 0; flappy_W(44, 455) <= 0; flappy_W(44, 456) <= 0; flappy_W(44, 457) <= 0; flappy_W(44, 458) <= 0; flappy_W(44, 459) <= 0; flappy_W(44, 460) <= 0; flappy_W(44, 461) <= 0; flappy_W(44, 462) <= 0; flappy_W(44, 463) <= 0; flappy_W(44, 464) <= 0; flappy_W(44, 465) <= 0; flappy_W(44, 466) <= 0; flappy_W(44, 467) <= 0; flappy_W(44, 468) <= 1; flappy_W(44, 469) <= 1; flappy_W(44, 470) <= 1; flappy_W(44, 471) <= 1; flappy_W(44, 472) <= 1; flappy_W(44, 473) <= 1; flappy_W(44, 474) <= 1; flappy_W(44, 475) <= 1; flappy_W(44, 476) <= 1; flappy_W(44, 477) <= 1; flappy_W(44, 478) <= 1; flappy_W(44, 479) <= 1; flappy_W(44, 480) <= 0; flappy_W(44, 481) <= 0; flappy_W(44, 482) <= 0; flappy_W(44, 483) <= 0; flappy_W(44, 484) <= 0; flappy_W(44, 485) <= 0; flappy_W(44, 486) <= 0; flappy_W(44, 487) <= 0; flappy_W(44, 488) <= 0; flappy_W(44, 489) <= 0; flappy_W(44, 490) <= 0; flappy_W(44, 491) <= 0; flappy_W(44, 492) <= 0; flappy_W(44, 493) <= 0; flappy_W(44, 494) <= 0; flappy_W(44, 495) <= 0; flappy_W(44, 496) <= 0; flappy_W(44, 497) <= 0; flappy_W(44, 498) <= 0; flappy_W(44, 499) <= 0; flappy_W(44, 500) <= 0; flappy_W(44, 501) <= 0; flappy_W(44, 502) <= 0; flappy_W(44, 503) <= 0; flappy_W(44, 504) <= 0; flappy_W(44, 505) <= 0; flappy_W(44, 506) <= 0; flappy_W(44, 507) <= 0; flappy_W(44, 508) <= 0; flappy_W(44, 509) <= 0; flappy_W(44, 510) <= 1; flappy_W(44, 511) <= 1; flappy_W(44, 512) <= 1; flappy_W(44, 513) <= 1; flappy_W(44, 514) <= 1; flappy_W(44, 515) <= 1; flappy_W(44, 516) <= 1; flappy_W(44, 517) <= 1; flappy_W(44, 518) <= 1; flappy_W(44, 519) <= 1; flappy_W(44, 520) <= 1; flappy_W(44, 521) <= 1; flappy_W(44, 522) <= 0; flappy_W(44, 523) <= 0; flappy_W(44, 524) <= 0; flappy_W(44, 525) <= 0; flappy_W(44, 526) <= 0; flappy_W(44, 527) <= 0; flappy_W(44, 528) <= 0; flappy_W(44, 529) <= 0; flappy_W(44, 530) <= 0; flappy_W(44, 531) <= 0; flappy_W(44, 532) <= 0; flappy_W(44, 533) <= 0; flappy_W(44, 534) <= 1; flappy_W(44, 535) <= 1; flappy_W(44, 536) <= 1; flappy_W(44, 537) <= 1; flappy_W(44, 538) <= 1; flappy_W(44, 539) <= 1; flappy_W(44, 540) <= 1; flappy_W(44, 541) <= 1; flappy_W(44, 542) <= 1; flappy_W(44, 543) <= 1; flappy_W(44, 544) <= 1; flappy_W(44, 545) <= 1; flappy_W(44, 546) <= 0; flappy_W(44, 547) <= 0; flappy_W(44, 548) <= 0; flappy_W(44, 549) <= 0; flappy_W(44, 550) <= 0; flappy_W(44, 551) <= 0; flappy_W(44, 552) <= 0; flappy_W(44, 553) <= 0; flappy_W(44, 554) <= 0; flappy_W(44, 555) <= 0; flappy_W(44, 556) <= 0; flappy_W(44, 557) <= 0; flappy_W(44, 558) <= 0; flappy_W(44, 559) <= 0; flappy_W(44, 560) <= 0; flappy_W(44, 561) <= 0; flappy_W(44, 562) <= 0; flappy_W(44, 563) <= 0; flappy_W(44, 564) <= 1; flappy_W(44, 565) <= 1; flappy_W(44, 566) <= 1; flappy_W(44, 567) <= 1; flappy_W(44, 568) <= 1; flappy_W(44, 569) <= 1; flappy_W(44, 570) <= 1; flappy_W(44, 571) <= 1; flappy_W(44, 572) <= 1; flappy_W(44, 573) <= 1; flappy_W(44, 574) <= 1; flappy_W(44, 575) <= 1; flappy_W(44, 576) <= 0; flappy_W(44, 577) <= 0; flappy_W(44, 578) <= 0; flappy_W(44, 579) <= 0; flappy_W(44, 580) <= 0; flappy_W(44, 581) <= 0; flappy_W(44, 582) <= 0; flappy_W(44, 583) <= 0; flappy_W(44, 584) <= 0; flappy_W(44, 585) <= 0; flappy_W(44, 586) <= 0; flappy_W(44, 587) <= 0; flappy_W(44, 588) <= 1; flappy_W(44, 589) <= 1; flappy_W(44, 590) <= 1; flappy_W(44, 591) <= 1; flappy_W(44, 592) <= 1; flappy_W(44, 593) <= 1; 
flappy_W(45, 0) <= 0; flappy_W(45, 1) <= 0; flappy_W(45, 2) <= 0; flappy_W(45, 3) <= 0; flappy_W(45, 4) <= 0; flappy_W(45, 5) <= 0; flappy_W(45, 6) <= 1; flappy_W(45, 7) <= 1; flappy_W(45, 8) <= 1; flappy_W(45, 9) <= 1; flappy_W(45, 10) <= 1; flappy_W(45, 11) <= 1; flappy_W(45, 12) <= 1; flappy_W(45, 13) <= 1; flappy_W(45, 14) <= 1; flappy_W(45, 15) <= 1; flappy_W(45, 16) <= 1; flappy_W(45, 17) <= 1; flappy_W(45, 18) <= 0; flappy_W(45, 19) <= 0; flappy_W(45, 20) <= 0; flappy_W(45, 21) <= 0; flappy_W(45, 22) <= 0; flappy_W(45, 23) <= 0; flappy_W(45, 24) <= 0; flappy_W(45, 25) <= 0; flappy_W(45, 26) <= 0; flappy_W(45, 27) <= 0; flappy_W(45, 28) <= 0; flappy_W(45, 29) <= 0; flappy_W(45, 30) <= 0; flappy_W(45, 31) <= 0; flappy_W(45, 32) <= 0; flappy_W(45, 33) <= 0; flappy_W(45, 34) <= 0; flappy_W(45, 35) <= 0; flappy_W(45, 36) <= 0; flappy_W(45, 37) <= 0; flappy_W(45, 38) <= 0; flappy_W(45, 39) <= 0; flappy_W(45, 40) <= 0; flappy_W(45, 41) <= 0; flappy_W(45, 42) <= 0; flappy_W(45, 43) <= 0; flappy_W(45, 44) <= 0; flappy_W(45, 45) <= 0; flappy_W(45, 46) <= 0; flappy_W(45, 47) <= 0; flappy_W(45, 48) <= 0; flappy_W(45, 49) <= 0; flappy_W(45, 50) <= 0; flappy_W(45, 51) <= 0; flappy_W(45, 52) <= 0; flappy_W(45, 53) <= 0; flappy_W(45, 54) <= 0; flappy_W(45, 55) <= 0; flappy_W(45, 56) <= 0; flappy_W(45, 57) <= 0; flappy_W(45, 58) <= 0; flappy_W(45, 59) <= 0; flappy_W(45, 60) <= 1; flappy_W(45, 61) <= 1; flappy_W(45, 62) <= 1; flappy_W(45, 63) <= 1; flappy_W(45, 64) <= 1; flappy_W(45, 65) <= 1; flappy_W(45, 66) <= 1; flappy_W(45, 67) <= 1; flappy_W(45, 68) <= 1; flappy_W(45, 69) <= 1; flappy_W(45, 70) <= 1; flappy_W(45, 71) <= 1; flappy_W(45, 72) <= 0; flappy_W(45, 73) <= 0; flappy_W(45, 74) <= 0; flappy_W(45, 75) <= 0; flappy_W(45, 76) <= 0; flappy_W(45, 77) <= 0; flappy_W(45, 78) <= 0; flappy_W(45, 79) <= 0; flappy_W(45, 80) <= 0; flappy_W(45, 81) <= 0; flappy_W(45, 82) <= 0; flappy_W(45, 83) <= 0; flappy_W(45, 84) <= 0; flappy_W(45, 85) <= 0; flappy_W(45, 86) <= 0; flappy_W(45, 87) <= 0; flappy_W(45, 88) <= 0; flappy_W(45, 89) <= 0; flappy_W(45, 90) <= 1; flappy_W(45, 91) <= 1; flappy_W(45, 92) <= 1; flappy_W(45, 93) <= 1; flappy_W(45, 94) <= 1; flappy_W(45, 95) <= 1; flappy_W(45, 96) <= 0; flappy_W(45, 97) <= 0; flappy_W(45, 98) <= 0; flappy_W(45, 99) <= 0; flappy_W(45, 100) <= 0; flappy_W(45, 101) <= 0; flappy_W(45, 102) <= 0; flappy_W(45, 103) <= 0; flappy_W(45, 104) <= 0; flappy_W(45, 105) <= 0; flappy_W(45, 106) <= 0; flappy_W(45, 107) <= 0; flappy_W(45, 108) <= 1; flappy_W(45, 109) <= 1; flappy_W(45, 110) <= 1; flappy_W(45, 111) <= 1; flappy_W(45, 112) <= 1; flappy_W(45, 113) <= 1; flappy_W(45, 114) <= 1; flappy_W(45, 115) <= 1; flappy_W(45, 116) <= 1; flappy_W(45, 117) <= 1; flappy_W(45, 118) <= 1; flappy_W(45, 119) <= 1; flappy_W(45, 120) <= 0; flappy_W(45, 121) <= 0; flappy_W(45, 122) <= 0; flappy_W(45, 123) <= 0; flappy_W(45, 124) <= 0; flappy_W(45, 125) <= 0; flappy_W(45, 126) <= 0; flappy_W(45, 127) <= 0; flappy_W(45, 128) <= 0; flappy_W(45, 129) <= 0; flappy_W(45, 130) <= 0; flappy_W(45, 131) <= 0; flappy_W(45, 132) <= 0; flappy_W(45, 133) <= 0; flappy_W(45, 134) <= 0; flappy_W(45, 135) <= 0; flappy_W(45, 136) <= 0; flappy_W(45, 137) <= 0; flappy_W(45, 138) <= 1; flappy_W(45, 139) <= 1; flappy_W(45, 140) <= 1; flappy_W(45, 141) <= 1; flappy_W(45, 142) <= 1; flappy_W(45, 143) <= 1; flappy_W(45, 144) <= 1; flappy_W(45, 145) <= 1; flappy_W(45, 146) <= 1; flappy_W(45, 147) <= 1; flappy_W(45, 148) <= 1; flappy_W(45, 149) <= 1; flappy_W(45, 150) <= 0; flappy_W(45, 151) <= 0; flappy_W(45, 152) <= 0; flappy_W(45, 153) <= 0; flappy_W(45, 154) <= 0; flappy_W(45, 155) <= 0; flappy_W(45, 156) <= 0; flappy_W(45, 157) <= 0; flappy_W(45, 158) <= 0; flappy_W(45, 159) <= 0; flappy_W(45, 160) <= 0; flappy_W(45, 161) <= 0; flappy_W(45, 162) <= 0; flappy_W(45, 163) <= 0; flappy_W(45, 164) <= 0; flappy_W(45, 165) <= 0; flappy_W(45, 166) <= 0; flappy_W(45, 167) <= 0; flappy_W(45, 168) <= 1; flappy_W(45, 169) <= 1; flappy_W(45, 170) <= 1; flappy_W(45, 171) <= 1; flappy_W(45, 172) <= 1; flappy_W(45, 173) <= 1; flappy_W(45, 174) <= 1; flappy_W(45, 175) <= 1; flappy_W(45, 176) <= 1; flappy_W(45, 177) <= 1; flappy_W(45, 178) <= 1; flappy_W(45, 179) <= 1; flappy_W(45, 180) <= 0; flappy_W(45, 181) <= 0; flappy_W(45, 182) <= 0; flappy_W(45, 183) <= 0; flappy_W(45, 184) <= 0; flappy_W(45, 185) <= 0; flappy_W(45, 186) <= 0; flappy_W(45, 187) <= 0; flappy_W(45, 188) <= 0; flappy_W(45, 189) <= 0; flappy_W(45, 190) <= 0; flappy_W(45, 191) <= 0; flappy_W(45, 192) <= 0; flappy_W(45, 193) <= 0; flappy_W(45, 194) <= 0; flappy_W(45, 195) <= 0; flappy_W(45, 196) <= 0; flappy_W(45, 197) <= 0; flappy_W(45, 198) <= 0; flappy_W(45, 199) <= 0; flappy_W(45, 200) <= 0; flappy_W(45, 201) <= 0; flappy_W(45, 202) <= 0; flappy_W(45, 203) <= 0; flappy_W(45, 204) <= 0; flappy_W(45, 205) <= 0; flappy_W(45, 206) <= 0; flappy_W(45, 207) <= 0; flappy_W(45, 208) <= 0; flappy_W(45, 209) <= 0; flappy_W(45, 210) <= 0; flappy_W(45, 211) <= 0; flappy_W(45, 212) <= 0; flappy_W(45, 213) <= 0; flappy_W(45, 214) <= 0; flappy_W(45, 215) <= 0; flappy_W(45, 216) <= 0; flappy_W(45, 217) <= 0; flappy_W(45, 218) <= 0; flappy_W(45, 219) <= 0; flappy_W(45, 220) <= 0; flappy_W(45, 221) <= 0; flappy_W(45, 222) <= 1; flappy_W(45, 223) <= 1; flappy_W(45, 224) <= 1; flappy_W(45, 225) <= 1; flappy_W(45, 226) <= 1; flappy_W(45, 227) <= 1; flappy_W(45, 228) <= 1; flappy_W(45, 229) <= 1; flappy_W(45, 230) <= 1; flappy_W(45, 231) <= 1; flappy_W(45, 232) <= 1; flappy_W(45, 233) <= 1; flappy_W(45, 234) <= 0; flappy_W(45, 235) <= 0; flappy_W(45, 236) <= 0; flappy_W(45, 237) <= 0; flappy_W(45, 238) <= 0; flappy_W(45, 239) <= 0; flappy_W(45, 240) <= 0; flappy_W(45, 241) <= 0; flappy_W(45, 242) <= 0; flappy_W(45, 243) <= 0; flappy_W(45, 244) <= 0; flappy_W(45, 245) <= 0; flappy_W(45, 246) <= 0; flappy_W(45, 247) <= 0; flappy_W(45, 248) <= 0; flappy_W(45, 249) <= 0; flappy_W(45, 250) <= 0; flappy_W(45, 251) <= 0; flappy_W(45, 252) <= 0; flappy_W(45, 253) <= 0; flappy_W(45, 254) <= 0; flappy_W(45, 255) <= 0; flappy_W(45, 256) <= 0; flappy_W(45, 257) <= 0; flappy_W(45, 258) <= 0; flappy_W(45, 259) <= 0; flappy_W(45, 260) <= 0; flappy_W(45, 261) <= 0; flappy_W(45, 262) <= 0; flappy_W(45, 263) <= 0; flappy_W(45, 264) <= 0; flappy_W(45, 265) <= 0; flappy_W(45, 266) <= 0; flappy_W(45, 267) <= 0; flappy_W(45, 268) <= 0; flappy_W(45, 269) <= 0; flappy_W(45, 270) <= 0; flappy_W(45, 271) <= 0; flappy_W(45, 272) <= 0; flappy_W(45, 273) <= 0; flappy_W(45, 274) <= 0; flappy_W(45, 275) <= 0; flappy_W(45, 276) <= 0; flappy_W(45, 277) <= 0; flappy_W(45, 278) <= 0; flappy_W(45, 279) <= 0; flappy_W(45, 280) <= 0; flappy_W(45, 281) <= 0; flappy_W(45, 282) <= 0; flappy_W(45, 283) <= 0; flappy_W(45, 284) <= 0; flappy_W(45, 285) <= 0; flappy_W(45, 286) <= 0; flappy_W(45, 287) <= 0; flappy_W(45, 288) <= 1; flappy_W(45, 289) <= 1; flappy_W(45, 290) <= 1; flappy_W(45, 291) <= 1; flappy_W(45, 292) <= 1; flappy_W(45, 293) <= 1; flappy_W(45, 294) <= 1; flappy_W(45, 295) <= 1; flappy_W(45, 296) <= 1; flappy_W(45, 297) <= 1; flappy_W(45, 298) <= 1; flappy_W(45, 299) <= 1; flappy_W(45, 300) <= 0; flappy_W(45, 301) <= 0; flappy_W(45, 302) <= 0; flappy_W(45, 303) <= 0; flappy_W(45, 304) <= 0; flappy_W(45, 305) <= 0; flappy_W(45, 306) <= 0; flappy_W(45, 307) <= 0; flappy_W(45, 308) <= 0; flappy_W(45, 309) <= 0; flappy_W(45, 310) <= 0; flappy_W(45, 311) <= 0; flappy_W(45, 312) <= 0; flappy_W(45, 313) <= 0; flappy_W(45, 314) <= 0; flappy_W(45, 315) <= 0; flappy_W(45, 316) <= 0; flappy_W(45, 317) <= 0; flappy_W(45, 318) <= 0; flappy_W(45, 319) <= 0; flappy_W(45, 320) <= 0; flappy_W(45, 321) <= 0; flappy_W(45, 322) <= 0; flappy_W(45, 323) <= 0; flappy_W(45, 324) <= 0; flappy_W(45, 325) <= 0; flappy_W(45, 326) <= 0; flappy_W(45, 327) <= 0; flappy_W(45, 328) <= 0; flappy_W(45, 329) <= 0; flappy_W(45, 330) <= 0; flappy_W(45, 331) <= 0; flappy_W(45, 332) <= 0; flappy_W(45, 333) <= 0; flappy_W(45, 334) <= 0; flappy_W(45, 335) <= 0; flappy_W(45, 336) <= 0; flappy_W(45, 337) <= 0; flappy_W(45, 338) <= 0; flappy_W(45, 339) <= 0; flappy_W(45, 340) <= 0; flappy_W(45, 341) <= 0; flappy_W(45, 342) <= 0; flappy_W(45, 343) <= 0; flappy_W(45, 344) <= 0; flappy_W(45, 345) <= 0; flappy_W(45, 346) <= 0; flappy_W(45, 347) <= 0; flappy_W(45, 348) <= 0; flappy_W(45, 349) <= 0; flappy_W(45, 350) <= 0; flappy_W(45, 351) <= 0; flappy_W(45, 352) <= 0; flappy_W(45, 353) <= 0; flappy_W(45, 354) <= 0; flappy_W(45, 355) <= 0; flappy_W(45, 356) <= 0; flappy_W(45, 357) <= 0; flappy_W(45, 358) <= 0; flappy_W(45, 359) <= 0; flappy_W(45, 360) <= 0; flappy_W(45, 361) <= 0; flappy_W(45, 362) <= 0; flappy_W(45, 363) <= 0; flappy_W(45, 364) <= 0; flappy_W(45, 365) <= 0; flappy_W(45, 366) <= 0; flappy_W(45, 367) <= 0; flappy_W(45, 368) <= 0; flappy_W(45, 369) <= 0; flappy_W(45, 370) <= 0; flappy_W(45, 371) <= 0; flappy_W(45, 372) <= 0; flappy_W(45, 373) <= 0; flappy_W(45, 374) <= 0; flappy_W(45, 375) <= 0; flappy_W(45, 376) <= 0; flappy_W(45, 377) <= 0; flappy_W(45, 378) <= 0; flappy_W(45, 379) <= 0; flappy_W(45, 380) <= 0; flappy_W(45, 381) <= 0; flappy_W(45, 382) <= 0; flappy_W(45, 383) <= 0; flappy_W(45, 384) <= 0; flappy_W(45, 385) <= 0; flappy_W(45, 386) <= 0; flappy_W(45, 387) <= 0; flappy_W(45, 388) <= 0; flappy_W(45, 389) <= 0; flappy_W(45, 390) <= 0; flappy_W(45, 391) <= 0; flappy_W(45, 392) <= 0; flappy_W(45, 393) <= 0; flappy_W(45, 394) <= 0; flappy_W(45, 395) <= 0; flappy_W(45, 396) <= 0; flappy_W(45, 397) <= 0; flappy_W(45, 398) <= 0; flappy_W(45, 399) <= 0; flappy_W(45, 400) <= 0; flappy_W(45, 401) <= 0; flappy_W(45, 402) <= 1; flappy_W(45, 403) <= 1; flappy_W(45, 404) <= 1; flappy_W(45, 405) <= 1; flappy_W(45, 406) <= 1; flappy_W(45, 407) <= 1; flappy_W(45, 408) <= 1; flappy_W(45, 409) <= 1; flappy_W(45, 410) <= 1; flappy_W(45, 411) <= 1; flappy_W(45, 412) <= 1; flappy_W(45, 413) <= 1; flappy_W(45, 414) <= 0; flappy_W(45, 415) <= 0; flappy_W(45, 416) <= 0; flappy_W(45, 417) <= 0; flappy_W(45, 418) <= 0; flappy_W(45, 419) <= 0; flappy_W(45, 420) <= 0; flappy_W(45, 421) <= 0; flappy_W(45, 422) <= 0; flappy_W(45, 423) <= 0; flappy_W(45, 424) <= 0; flappy_W(45, 425) <= 0; flappy_W(45, 426) <= 1; flappy_W(45, 427) <= 1; flappy_W(45, 428) <= 1; flappy_W(45, 429) <= 1; flappy_W(45, 430) <= 1; flappy_W(45, 431) <= 1; flappy_W(45, 432) <= 1; flappy_W(45, 433) <= 1; flappy_W(45, 434) <= 1; flappy_W(45, 435) <= 1; flappy_W(45, 436) <= 1; flappy_W(45, 437) <= 1; flappy_W(45, 438) <= 0; flappy_W(45, 439) <= 0; flappy_W(45, 440) <= 0; flappy_W(45, 441) <= 0; flappy_W(45, 442) <= 0; flappy_W(45, 443) <= 0; flappy_W(45, 444) <= 0; flappy_W(45, 445) <= 0; flappy_W(45, 446) <= 0; flappy_W(45, 447) <= 0; flappy_W(45, 448) <= 0; flappy_W(45, 449) <= 0; flappy_W(45, 450) <= 0; flappy_W(45, 451) <= 0; flappy_W(45, 452) <= 0; flappy_W(45, 453) <= 0; flappy_W(45, 454) <= 0; flappy_W(45, 455) <= 0; flappy_W(45, 456) <= 0; flappy_W(45, 457) <= 0; flappy_W(45, 458) <= 0; flappy_W(45, 459) <= 0; flappy_W(45, 460) <= 0; flappy_W(45, 461) <= 0; flappy_W(45, 462) <= 0; flappy_W(45, 463) <= 0; flappy_W(45, 464) <= 0; flappy_W(45, 465) <= 0; flappy_W(45, 466) <= 0; flappy_W(45, 467) <= 0; flappy_W(45, 468) <= 1; flappy_W(45, 469) <= 1; flappy_W(45, 470) <= 1; flappy_W(45, 471) <= 1; flappy_W(45, 472) <= 1; flappy_W(45, 473) <= 1; flappy_W(45, 474) <= 1; flappy_W(45, 475) <= 1; flappy_W(45, 476) <= 1; flappy_W(45, 477) <= 1; flappy_W(45, 478) <= 1; flappy_W(45, 479) <= 1; flappy_W(45, 480) <= 0; flappy_W(45, 481) <= 0; flappy_W(45, 482) <= 0; flappy_W(45, 483) <= 0; flappy_W(45, 484) <= 0; flappy_W(45, 485) <= 0; flappy_W(45, 486) <= 0; flappy_W(45, 487) <= 0; flappy_W(45, 488) <= 0; flappy_W(45, 489) <= 0; flappy_W(45, 490) <= 0; flappy_W(45, 491) <= 0; flappy_W(45, 492) <= 0; flappy_W(45, 493) <= 0; flappy_W(45, 494) <= 0; flappy_W(45, 495) <= 0; flappy_W(45, 496) <= 0; flappy_W(45, 497) <= 0; flappy_W(45, 498) <= 0; flappy_W(45, 499) <= 0; flappy_W(45, 500) <= 0; flappy_W(45, 501) <= 0; flappy_W(45, 502) <= 0; flappy_W(45, 503) <= 0; flappy_W(45, 504) <= 0; flappy_W(45, 505) <= 0; flappy_W(45, 506) <= 0; flappy_W(45, 507) <= 0; flappy_W(45, 508) <= 0; flappy_W(45, 509) <= 0; flappy_W(45, 510) <= 1; flappy_W(45, 511) <= 1; flappy_W(45, 512) <= 1; flappy_W(45, 513) <= 1; flappy_W(45, 514) <= 1; flappy_W(45, 515) <= 1; flappy_W(45, 516) <= 1; flappy_W(45, 517) <= 1; flappy_W(45, 518) <= 1; flappy_W(45, 519) <= 1; flappy_W(45, 520) <= 1; flappy_W(45, 521) <= 1; flappy_W(45, 522) <= 0; flappy_W(45, 523) <= 0; flappy_W(45, 524) <= 0; flappy_W(45, 525) <= 0; flappy_W(45, 526) <= 0; flappy_W(45, 527) <= 0; flappy_W(45, 528) <= 0; flappy_W(45, 529) <= 0; flappy_W(45, 530) <= 0; flappy_W(45, 531) <= 0; flappy_W(45, 532) <= 0; flappy_W(45, 533) <= 0; flappy_W(45, 534) <= 1; flappy_W(45, 535) <= 1; flappy_W(45, 536) <= 1; flappy_W(45, 537) <= 1; flappy_W(45, 538) <= 1; flappy_W(45, 539) <= 1; flappy_W(45, 540) <= 1; flappy_W(45, 541) <= 1; flappy_W(45, 542) <= 1; flappy_W(45, 543) <= 1; flappy_W(45, 544) <= 1; flappy_W(45, 545) <= 1; flappy_W(45, 546) <= 0; flappy_W(45, 547) <= 0; flappy_W(45, 548) <= 0; flappy_W(45, 549) <= 0; flappy_W(45, 550) <= 0; flappy_W(45, 551) <= 0; flappy_W(45, 552) <= 0; flappy_W(45, 553) <= 0; flappy_W(45, 554) <= 0; flappy_W(45, 555) <= 0; flappy_W(45, 556) <= 0; flappy_W(45, 557) <= 0; flappy_W(45, 558) <= 0; flappy_W(45, 559) <= 0; flappy_W(45, 560) <= 0; flappy_W(45, 561) <= 0; flappy_W(45, 562) <= 0; flappy_W(45, 563) <= 0; flappy_W(45, 564) <= 1; flappy_W(45, 565) <= 1; flappy_W(45, 566) <= 1; flappy_W(45, 567) <= 1; flappy_W(45, 568) <= 1; flappy_W(45, 569) <= 1; flappy_W(45, 570) <= 1; flappy_W(45, 571) <= 1; flappy_W(45, 572) <= 1; flappy_W(45, 573) <= 1; flappy_W(45, 574) <= 1; flappy_W(45, 575) <= 1; flappy_W(45, 576) <= 0; flappy_W(45, 577) <= 0; flappy_W(45, 578) <= 0; flappy_W(45, 579) <= 0; flappy_W(45, 580) <= 0; flappy_W(45, 581) <= 0; flappy_W(45, 582) <= 0; flappy_W(45, 583) <= 0; flappy_W(45, 584) <= 0; flappy_W(45, 585) <= 0; flappy_W(45, 586) <= 0; flappy_W(45, 587) <= 0; flappy_W(45, 588) <= 1; flappy_W(45, 589) <= 1; flappy_W(45, 590) <= 1; flappy_W(45, 591) <= 1; flappy_W(45, 592) <= 1; flappy_W(45, 593) <= 1; 
flappy_W(46, 0) <= 0; flappy_W(46, 1) <= 0; flappy_W(46, 2) <= 0; flappy_W(46, 3) <= 0; flappy_W(46, 4) <= 0; flappy_W(46, 5) <= 0; flappy_W(46, 6) <= 1; flappy_W(46, 7) <= 1; flappy_W(46, 8) <= 1; flappy_W(46, 9) <= 1; flappy_W(46, 10) <= 1; flappy_W(46, 11) <= 1; flappy_W(46, 12) <= 1; flappy_W(46, 13) <= 1; flappy_W(46, 14) <= 1; flappy_W(46, 15) <= 1; flappy_W(46, 16) <= 1; flappy_W(46, 17) <= 1; flappy_W(46, 18) <= 0; flappy_W(46, 19) <= 0; flappy_W(46, 20) <= 0; flappy_W(46, 21) <= 0; flappy_W(46, 22) <= 0; flappy_W(46, 23) <= 0; flappy_W(46, 24) <= 0; flappy_W(46, 25) <= 0; flappy_W(46, 26) <= 0; flappy_W(46, 27) <= 0; flappy_W(46, 28) <= 0; flappy_W(46, 29) <= 0; flappy_W(46, 30) <= 0; flappy_W(46, 31) <= 0; flappy_W(46, 32) <= 0; flappy_W(46, 33) <= 0; flappy_W(46, 34) <= 0; flappy_W(46, 35) <= 0; flappy_W(46, 36) <= 0; flappy_W(46, 37) <= 0; flappy_W(46, 38) <= 0; flappy_W(46, 39) <= 0; flappy_W(46, 40) <= 0; flappy_W(46, 41) <= 0; flappy_W(46, 42) <= 0; flappy_W(46, 43) <= 0; flappy_W(46, 44) <= 0; flappy_W(46, 45) <= 0; flappy_W(46, 46) <= 0; flappy_W(46, 47) <= 0; flappy_W(46, 48) <= 0; flappy_W(46, 49) <= 0; flappy_W(46, 50) <= 0; flappy_W(46, 51) <= 0; flappy_W(46, 52) <= 0; flappy_W(46, 53) <= 0; flappy_W(46, 54) <= 0; flappy_W(46, 55) <= 0; flappy_W(46, 56) <= 0; flappy_W(46, 57) <= 0; flappy_W(46, 58) <= 0; flappy_W(46, 59) <= 0; flappy_W(46, 60) <= 1; flappy_W(46, 61) <= 1; flappy_W(46, 62) <= 1; flappy_W(46, 63) <= 1; flappy_W(46, 64) <= 1; flappy_W(46, 65) <= 1; flappy_W(46, 66) <= 1; flappy_W(46, 67) <= 1; flappy_W(46, 68) <= 1; flappy_W(46, 69) <= 1; flappy_W(46, 70) <= 1; flappy_W(46, 71) <= 1; flappy_W(46, 72) <= 0; flappy_W(46, 73) <= 0; flappy_W(46, 74) <= 0; flappy_W(46, 75) <= 0; flappy_W(46, 76) <= 0; flappy_W(46, 77) <= 0; flappy_W(46, 78) <= 0; flappy_W(46, 79) <= 0; flappy_W(46, 80) <= 0; flappy_W(46, 81) <= 0; flappy_W(46, 82) <= 0; flappy_W(46, 83) <= 0; flappy_W(46, 84) <= 0; flappy_W(46, 85) <= 0; flappy_W(46, 86) <= 0; flappy_W(46, 87) <= 0; flappy_W(46, 88) <= 0; flappy_W(46, 89) <= 0; flappy_W(46, 90) <= 1; flappy_W(46, 91) <= 1; flappy_W(46, 92) <= 1; flappy_W(46, 93) <= 1; flappy_W(46, 94) <= 1; flappy_W(46, 95) <= 1; flappy_W(46, 96) <= 0; flappy_W(46, 97) <= 0; flappy_W(46, 98) <= 0; flappy_W(46, 99) <= 0; flappy_W(46, 100) <= 0; flappy_W(46, 101) <= 0; flappy_W(46, 102) <= 0; flappy_W(46, 103) <= 0; flappy_W(46, 104) <= 0; flappy_W(46, 105) <= 0; flappy_W(46, 106) <= 0; flappy_W(46, 107) <= 0; flappy_W(46, 108) <= 1; flappy_W(46, 109) <= 1; flappy_W(46, 110) <= 1; flappy_W(46, 111) <= 1; flappy_W(46, 112) <= 1; flappy_W(46, 113) <= 1; flappy_W(46, 114) <= 1; flappy_W(46, 115) <= 1; flappy_W(46, 116) <= 1; flappy_W(46, 117) <= 1; flappy_W(46, 118) <= 1; flappy_W(46, 119) <= 1; flappy_W(46, 120) <= 0; flappy_W(46, 121) <= 0; flappy_W(46, 122) <= 0; flappy_W(46, 123) <= 0; flappy_W(46, 124) <= 0; flappy_W(46, 125) <= 0; flappy_W(46, 126) <= 0; flappy_W(46, 127) <= 0; flappy_W(46, 128) <= 0; flappy_W(46, 129) <= 0; flappy_W(46, 130) <= 0; flappy_W(46, 131) <= 0; flappy_W(46, 132) <= 0; flappy_W(46, 133) <= 0; flappy_W(46, 134) <= 0; flappy_W(46, 135) <= 0; flappy_W(46, 136) <= 0; flappy_W(46, 137) <= 0; flappy_W(46, 138) <= 1; flappy_W(46, 139) <= 1; flappy_W(46, 140) <= 1; flappy_W(46, 141) <= 1; flappy_W(46, 142) <= 1; flappy_W(46, 143) <= 1; flappy_W(46, 144) <= 1; flappy_W(46, 145) <= 1; flappy_W(46, 146) <= 1; flappy_W(46, 147) <= 1; flappy_W(46, 148) <= 1; flappy_W(46, 149) <= 1; flappy_W(46, 150) <= 0; flappy_W(46, 151) <= 0; flappy_W(46, 152) <= 0; flappy_W(46, 153) <= 0; flappy_W(46, 154) <= 0; flappy_W(46, 155) <= 0; flappy_W(46, 156) <= 0; flappy_W(46, 157) <= 0; flappy_W(46, 158) <= 0; flappy_W(46, 159) <= 0; flappy_W(46, 160) <= 0; flappy_W(46, 161) <= 0; flappy_W(46, 162) <= 0; flappy_W(46, 163) <= 0; flappy_W(46, 164) <= 0; flappy_W(46, 165) <= 0; flappy_W(46, 166) <= 0; flappy_W(46, 167) <= 0; flappy_W(46, 168) <= 1; flappy_W(46, 169) <= 1; flappy_W(46, 170) <= 1; flappy_W(46, 171) <= 1; flappy_W(46, 172) <= 1; flappy_W(46, 173) <= 1; flappy_W(46, 174) <= 1; flappy_W(46, 175) <= 1; flappy_W(46, 176) <= 1; flappy_W(46, 177) <= 1; flappy_W(46, 178) <= 1; flappy_W(46, 179) <= 1; flappy_W(46, 180) <= 0; flappy_W(46, 181) <= 0; flappy_W(46, 182) <= 0; flappy_W(46, 183) <= 0; flappy_W(46, 184) <= 0; flappy_W(46, 185) <= 0; flappy_W(46, 186) <= 0; flappy_W(46, 187) <= 0; flappy_W(46, 188) <= 0; flappy_W(46, 189) <= 0; flappy_W(46, 190) <= 0; flappy_W(46, 191) <= 0; flappy_W(46, 192) <= 0; flappy_W(46, 193) <= 0; flappy_W(46, 194) <= 0; flappy_W(46, 195) <= 0; flappy_W(46, 196) <= 0; flappy_W(46, 197) <= 0; flappy_W(46, 198) <= 0; flappy_W(46, 199) <= 0; flappy_W(46, 200) <= 0; flappy_W(46, 201) <= 0; flappy_W(46, 202) <= 0; flappy_W(46, 203) <= 0; flappy_W(46, 204) <= 0; flappy_W(46, 205) <= 0; flappy_W(46, 206) <= 0; flappy_W(46, 207) <= 0; flappy_W(46, 208) <= 0; flappy_W(46, 209) <= 0; flappy_W(46, 210) <= 0; flappy_W(46, 211) <= 0; flappy_W(46, 212) <= 0; flappy_W(46, 213) <= 0; flappy_W(46, 214) <= 0; flappy_W(46, 215) <= 0; flappy_W(46, 216) <= 0; flappy_W(46, 217) <= 0; flappy_W(46, 218) <= 0; flappy_W(46, 219) <= 0; flappy_W(46, 220) <= 0; flappy_W(46, 221) <= 0; flappy_W(46, 222) <= 1; flappy_W(46, 223) <= 1; flappy_W(46, 224) <= 1; flappy_W(46, 225) <= 1; flappy_W(46, 226) <= 1; flappy_W(46, 227) <= 1; flappy_W(46, 228) <= 1; flappy_W(46, 229) <= 1; flappy_W(46, 230) <= 1; flappy_W(46, 231) <= 1; flappy_W(46, 232) <= 1; flappy_W(46, 233) <= 1; flappy_W(46, 234) <= 0; flappy_W(46, 235) <= 0; flappy_W(46, 236) <= 0; flappy_W(46, 237) <= 0; flappy_W(46, 238) <= 0; flappy_W(46, 239) <= 0; flappy_W(46, 240) <= 0; flappy_W(46, 241) <= 0; flappy_W(46, 242) <= 0; flappy_W(46, 243) <= 0; flappy_W(46, 244) <= 0; flappy_W(46, 245) <= 0; flappy_W(46, 246) <= 0; flappy_W(46, 247) <= 0; flappy_W(46, 248) <= 0; flappy_W(46, 249) <= 0; flappy_W(46, 250) <= 0; flappy_W(46, 251) <= 0; flappy_W(46, 252) <= 0; flappy_W(46, 253) <= 0; flappy_W(46, 254) <= 0; flappy_W(46, 255) <= 0; flappy_W(46, 256) <= 0; flappy_W(46, 257) <= 0; flappy_W(46, 258) <= 0; flappy_W(46, 259) <= 0; flappy_W(46, 260) <= 0; flappy_W(46, 261) <= 0; flappy_W(46, 262) <= 0; flappy_W(46, 263) <= 0; flappy_W(46, 264) <= 0; flappy_W(46, 265) <= 0; flappy_W(46, 266) <= 0; flappy_W(46, 267) <= 0; flappy_W(46, 268) <= 0; flappy_W(46, 269) <= 0; flappy_W(46, 270) <= 0; flappy_W(46, 271) <= 0; flappy_W(46, 272) <= 0; flappy_W(46, 273) <= 0; flappy_W(46, 274) <= 0; flappy_W(46, 275) <= 0; flappy_W(46, 276) <= 0; flappy_W(46, 277) <= 0; flappy_W(46, 278) <= 0; flappy_W(46, 279) <= 0; flappy_W(46, 280) <= 0; flappy_W(46, 281) <= 0; flappy_W(46, 282) <= 0; flappy_W(46, 283) <= 0; flappy_W(46, 284) <= 0; flappy_W(46, 285) <= 0; flappy_W(46, 286) <= 0; flappy_W(46, 287) <= 0; flappy_W(46, 288) <= 1; flappy_W(46, 289) <= 1; flappy_W(46, 290) <= 1; flappy_W(46, 291) <= 1; flappy_W(46, 292) <= 1; flappy_W(46, 293) <= 1; flappy_W(46, 294) <= 1; flappy_W(46, 295) <= 1; flappy_W(46, 296) <= 1; flappy_W(46, 297) <= 1; flappy_W(46, 298) <= 1; flappy_W(46, 299) <= 1; flappy_W(46, 300) <= 0; flappy_W(46, 301) <= 0; flappy_W(46, 302) <= 0; flappy_W(46, 303) <= 0; flappy_W(46, 304) <= 0; flappy_W(46, 305) <= 0; flappy_W(46, 306) <= 0; flappy_W(46, 307) <= 0; flappy_W(46, 308) <= 0; flappy_W(46, 309) <= 0; flappy_W(46, 310) <= 0; flappy_W(46, 311) <= 0; flappy_W(46, 312) <= 0; flappy_W(46, 313) <= 0; flappy_W(46, 314) <= 0; flappy_W(46, 315) <= 0; flappy_W(46, 316) <= 0; flappy_W(46, 317) <= 0; flappy_W(46, 318) <= 0; flappy_W(46, 319) <= 0; flappy_W(46, 320) <= 0; flappy_W(46, 321) <= 0; flappy_W(46, 322) <= 0; flappy_W(46, 323) <= 0; flappy_W(46, 324) <= 0; flappy_W(46, 325) <= 0; flappy_W(46, 326) <= 0; flappy_W(46, 327) <= 0; flappy_W(46, 328) <= 0; flappy_W(46, 329) <= 0; flappy_W(46, 330) <= 0; flappy_W(46, 331) <= 0; flappy_W(46, 332) <= 0; flappy_W(46, 333) <= 0; flappy_W(46, 334) <= 0; flappy_W(46, 335) <= 0; flappy_W(46, 336) <= 0; flappy_W(46, 337) <= 0; flappy_W(46, 338) <= 0; flappy_W(46, 339) <= 0; flappy_W(46, 340) <= 0; flappy_W(46, 341) <= 0; flappy_W(46, 342) <= 0; flappy_W(46, 343) <= 0; flappy_W(46, 344) <= 0; flappy_W(46, 345) <= 0; flappy_W(46, 346) <= 0; flappy_W(46, 347) <= 0; flappy_W(46, 348) <= 0; flappy_W(46, 349) <= 0; flappy_W(46, 350) <= 0; flappy_W(46, 351) <= 0; flappy_W(46, 352) <= 0; flappy_W(46, 353) <= 0; flappy_W(46, 354) <= 0; flappy_W(46, 355) <= 0; flappy_W(46, 356) <= 0; flappy_W(46, 357) <= 0; flappy_W(46, 358) <= 0; flappy_W(46, 359) <= 0; flappy_W(46, 360) <= 0; flappy_W(46, 361) <= 0; flappy_W(46, 362) <= 0; flappy_W(46, 363) <= 0; flappy_W(46, 364) <= 0; flappy_W(46, 365) <= 0; flappy_W(46, 366) <= 0; flappy_W(46, 367) <= 0; flappy_W(46, 368) <= 0; flappy_W(46, 369) <= 0; flappy_W(46, 370) <= 0; flappy_W(46, 371) <= 0; flappy_W(46, 372) <= 0; flappy_W(46, 373) <= 0; flappy_W(46, 374) <= 0; flappy_W(46, 375) <= 0; flappy_W(46, 376) <= 0; flappy_W(46, 377) <= 0; flappy_W(46, 378) <= 0; flappy_W(46, 379) <= 0; flappy_W(46, 380) <= 0; flappy_W(46, 381) <= 0; flappy_W(46, 382) <= 0; flappy_W(46, 383) <= 0; flappy_W(46, 384) <= 0; flappy_W(46, 385) <= 0; flappy_W(46, 386) <= 0; flappy_W(46, 387) <= 0; flappy_W(46, 388) <= 0; flappy_W(46, 389) <= 0; flappy_W(46, 390) <= 0; flappy_W(46, 391) <= 0; flappy_W(46, 392) <= 0; flappy_W(46, 393) <= 0; flappy_W(46, 394) <= 0; flappy_W(46, 395) <= 0; flappy_W(46, 396) <= 0; flappy_W(46, 397) <= 0; flappy_W(46, 398) <= 0; flappy_W(46, 399) <= 0; flappy_W(46, 400) <= 0; flappy_W(46, 401) <= 0; flappy_W(46, 402) <= 1; flappy_W(46, 403) <= 1; flappy_W(46, 404) <= 1; flappy_W(46, 405) <= 1; flappy_W(46, 406) <= 1; flappy_W(46, 407) <= 1; flappy_W(46, 408) <= 1; flappy_W(46, 409) <= 1; flappy_W(46, 410) <= 1; flappy_W(46, 411) <= 1; flappy_W(46, 412) <= 1; flappy_W(46, 413) <= 1; flappy_W(46, 414) <= 0; flappy_W(46, 415) <= 0; flappy_W(46, 416) <= 0; flappy_W(46, 417) <= 0; flappy_W(46, 418) <= 0; flappy_W(46, 419) <= 0; flappy_W(46, 420) <= 0; flappy_W(46, 421) <= 0; flappy_W(46, 422) <= 0; flappy_W(46, 423) <= 0; flappy_W(46, 424) <= 0; flappy_W(46, 425) <= 0; flappy_W(46, 426) <= 1; flappy_W(46, 427) <= 1; flappy_W(46, 428) <= 1; flappy_W(46, 429) <= 1; flappy_W(46, 430) <= 1; flappy_W(46, 431) <= 1; flappy_W(46, 432) <= 1; flappy_W(46, 433) <= 1; flappy_W(46, 434) <= 1; flappy_W(46, 435) <= 1; flappy_W(46, 436) <= 1; flappy_W(46, 437) <= 1; flappy_W(46, 438) <= 0; flappy_W(46, 439) <= 0; flappy_W(46, 440) <= 0; flappy_W(46, 441) <= 0; flappy_W(46, 442) <= 0; flappy_W(46, 443) <= 0; flappy_W(46, 444) <= 0; flappy_W(46, 445) <= 0; flappy_W(46, 446) <= 0; flappy_W(46, 447) <= 0; flappy_W(46, 448) <= 0; flappy_W(46, 449) <= 0; flappy_W(46, 450) <= 0; flappy_W(46, 451) <= 0; flappy_W(46, 452) <= 0; flappy_W(46, 453) <= 0; flappy_W(46, 454) <= 0; flappy_W(46, 455) <= 0; flappy_W(46, 456) <= 0; flappy_W(46, 457) <= 0; flappy_W(46, 458) <= 0; flappy_W(46, 459) <= 0; flappy_W(46, 460) <= 0; flappy_W(46, 461) <= 0; flappy_W(46, 462) <= 0; flappy_W(46, 463) <= 0; flappy_W(46, 464) <= 0; flappy_W(46, 465) <= 0; flappy_W(46, 466) <= 0; flappy_W(46, 467) <= 0; flappy_W(46, 468) <= 1; flappy_W(46, 469) <= 1; flappy_W(46, 470) <= 1; flappy_W(46, 471) <= 1; flappy_W(46, 472) <= 1; flappy_W(46, 473) <= 1; flappy_W(46, 474) <= 1; flappy_W(46, 475) <= 1; flappy_W(46, 476) <= 1; flappy_W(46, 477) <= 1; flappy_W(46, 478) <= 1; flappy_W(46, 479) <= 1; flappy_W(46, 480) <= 0; flappy_W(46, 481) <= 0; flappy_W(46, 482) <= 0; flappy_W(46, 483) <= 0; flappy_W(46, 484) <= 0; flappy_W(46, 485) <= 0; flappy_W(46, 486) <= 0; flappy_W(46, 487) <= 0; flappy_W(46, 488) <= 0; flappy_W(46, 489) <= 0; flappy_W(46, 490) <= 0; flappy_W(46, 491) <= 0; flappy_W(46, 492) <= 0; flappy_W(46, 493) <= 0; flappy_W(46, 494) <= 0; flappy_W(46, 495) <= 0; flappy_W(46, 496) <= 0; flappy_W(46, 497) <= 0; flappy_W(46, 498) <= 0; flappy_W(46, 499) <= 0; flappy_W(46, 500) <= 0; flappy_W(46, 501) <= 0; flappy_W(46, 502) <= 0; flappy_W(46, 503) <= 0; flappy_W(46, 504) <= 0; flappy_W(46, 505) <= 0; flappy_W(46, 506) <= 0; flappy_W(46, 507) <= 0; flappy_W(46, 508) <= 0; flappy_W(46, 509) <= 0; flappy_W(46, 510) <= 1; flappy_W(46, 511) <= 1; flappy_W(46, 512) <= 1; flappy_W(46, 513) <= 1; flappy_W(46, 514) <= 1; flappy_W(46, 515) <= 1; flappy_W(46, 516) <= 1; flappy_W(46, 517) <= 1; flappy_W(46, 518) <= 1; flappy_W(46, 519) <= 1; flappy_W(46, 520) <= 1; flappy_W(46, 521) <= 1; flappy_W(46, 522) <= 0; flappy_W(46, 523) <= 0; flappy_W(46, 524) <= 0; flappy_W(46, 525) <= 0; flappy_W(46, 526) <= 0; flappy_W(46, 527) <= 0; flappy_W(46, 528) <= 0; flappy_W(46, 529) <= 0; flappy_W(46, 530) <= 0; flappy_W(46, 531) <= 0; flappy_W(46, 532) <= 0; flappy_W(46, 533) <= 0; flappy_W(46, 534) <= 1; flappy_W(46, 535) <= 1; flappy_W(46, 536) <= 1; flappy_W(46, 537) <= 1; flappy_W(46, 538) <= 1; flappy_W(46, 539) <= 1; flappy_W(46, 540) <= 1; flappy_W(46, 541) <= 1; flappy_W(46, 542) <= 1; flappy_W(46, 543) <= 1; flappy_W(46, 544) <= 1; flappy_W(46, 545) <= 1; flappy_W(46, 546) <= 0; flappy_W(46, 547) <= 0; flappy_W(46, 548) <= 0; flappy_W(46, 549) <= 0; flappy_W(46, 550) <= 0; flappy_W(46, 551) <= 0; flappy_W(46, 552) <= 0; flappy_W(46, 553) <= 0; flappy_W(46, 554) <= 0; flappy_W(46, 555) <= 0; flappy_W(46, 556) <= 0; flappy_W(46, 557) <= 0; flappy_W(46, 558) <= 0; flappy_W(46, 559) <= 0; flappy_W(46, 560) <= 0; flappy_W(46, 561) <= 0; flappy_W(46, 562) <= 0; flappy_W(46, 563) <= 0; flappy_W(46, 564) <= 1; flappy_W(46, 565) <= 1; flappy_W(46, 566) <= 1; flappy_W(46, 567) <= 1; flappy_W(46, 568) <= 1; flappy_W(46, 569) <= 1; flappy_W(46, 570) <= 1; flappy_W(46, 571) <= 1; flappy_W(46, 572) <= 1; flappy_W(46, 573) <= 1; flappy_W(46, 574) <= 1; flappy_W(46, 575) <= 1; flappy_W(46, 576) <= 0; flappy_W(46, 577) <= 0; flappy_W(46, 578) <= 0; flappy_W(46, 579) <= 0; flappy_W(46, 580) <= 0; flappy_W(46, 581) <= 0; flappy_W(46, 582) <= 0; flappy_W(46, 583) <= 0; flappy_W(46, 584) <= 0; flappy_W(46, 585) <= 0; flappy_W(46, 586) <= 0; flappy_W(46, 587) <= 0; flappy_W(46, 588) <= 1; flappy_W(46, 589) <= 1; flappy_W(46, 590) <= 1; flappy_W(46, 591) <= 1; flappy_W(46, 592) <= 1; flappy_W(46, 593) <= 1; 
flappy_W(47, 0) <= 0; flappy_W(47, 1) <= 0; flappy_W(47, 2) <= 0; flappy_W(47, 3) <= 0; flappy_W(47, 4) <= 0; flappy_W(47, 5) <= 0; flappy_W(47, 6) <= 1; flappy_W(47, 7) <= 1; flappy_W(47, 8) <= 1; flappy_W(47, 9) <= 1; flappy_W(47, 10) <= 1; flappy_W(47, 11) <= 1; flappy_W(47, 12) <= 1; flappy_W(47, 13) <= 1; flappy_W(47, 14) <= 1; flappy_W(47, 15) <= 1; flappy_W(47, 16) <= 1; flappy_W(47, 17) <= 1; flappy_W(47, 18) <= 0; flappy_W(47, 19) <= 0; flappy_W(47, 20) <= 0; flappy_W(47, 21) <= 0; flappy_W(47, 22) <= 0; flappy_W(47, 23) <= 0; flappy_W(47, 24) <= 0; flappy_W(47, 25) <= 0; flappy_W(47, 26) <= 0; flappy_W(47, 27) <= 0; flappy_W(47, 28) <= 0; flappy_W(47, 29) <= 0; flappy_W(47, 30) <= 0; flappy_W(47, 31) <= 0; flappy_W(47, 32) <= 0; flappy_W(47, 33) <= 0; flappy_W(47, 34) <= 0; flappy_W(47, 35) <= 0; flappy_W(47, 36) <= 0; flappy_W(47, 37) <= 0; flappy_W(47, 38) <= 0; flappy_W(47, 39) <= 0; flappy_W(47, 40) <= 0; flappy_W(47, 41) <= 0; flappy_W(47, 42) <= 0; flappy_W(47, 43) <= 0; flappy_W(47, 44) <= 0; flappy_W(47, 45) <= 0; flappy_W(47, 46) <= 0; flappy_W(47, 47) <= 0; flappy_W(47, 48) <= 0; flappy_W(47, 49) <= 0; flappy_W(47, 50) <= 0; flappy_W(47, 51) <= 0; flappy_W(47, 52) <= 0; flappy_W(47, 53) <= 0; flappy_W(47, 54) <= 0; flappy_W(47, 55) <= 0; flappy_W(47, 56) <= 0; flappy_W(47, 57) <= 0; flappy_W(47, 58) <= 0; flappy_W(47, 59) <= 0; flappy_W(47, 60) <= 1; flappy_W(47, 61) <= 1; flappy_W(47, 62) <= 1; flappy_W(47, 63) <= 1; flappy_W(47, 64) <= 1; flappy_W(47, 65) <= 1; flappy_W(47, 66) <= 1; flappy_W(47, 67) <= 1; flappy_W(47, 68) <= 1; flappy_W(47, 69) <= 1; flappy_W(47, 70) <= 1; flappy_W(47, 71) <= 1; flappy_W(47, 72) <= 0; flappy_W(47, 73) <= 0; flappy_W(47, 74) <= 0; flappy_W(47, 75) <= 0; flappy_W(47, 76) <= 0; flappy_W(47, 77) <= 0; flappy_W(47, 78) <= 0; flappy_W(47, 79) <= 0; flappy_W(47, 80) <= 0; flappy_W(47, 81) <= 0; flappy_W(47, 82) <= 0; flappy_W(47, 83) <= 0; flappy_W(47, 84) <= 0; flappy_W(47, 85) <= 0; flappy_W(47, 86) <= 0; flappy_W(47, 87) <= 0; flappy_W(47, 88) <= 0; flappy_W(47, 89) <= 0; flappy_W(47, 90) <= 1; flappy_W(47, 91) <= 1; flappy_W(47, 92) <= 1; flappy_W(47, 93) <= 1; flappy_W(47, 94) <= 1; flappy_W(47, 95) <= 1; flappy_W(47, 96) <= 0; flappy_W(47, 97) <= 0; flappy_W(47, 98) <= 0; flappy_W(47, 99) <= 0; flappy_W(47, 100) <= 0; flappy_W(47, 101) <= 0; flappy_W(47, 102) <= 0; flappy_W(47, 103) <= 0; flappy_W(47, 104) <= 0; flappy_W(47, 105) <= 0; flappy_W(47, 106) <= 0; flappy_W(47, 107) <= 0; flappy_W(47, 108) <= 1; flappy_W(47, 109) <= 1; flappy_W(47, 110) <= 1; flappy_W(47, 111) <= 1; flappy_W(47, 112) <= 1; flappy_W(47, 113) <= 1; flappy_W(47, 114) <= 1; flappy_W(47, 115) <= 1; flappy_W(47, 116) <= 1; flappy_W(47, 117) <= 1; flappy_W(47, 118) <= 1; flappy_W(47, 119) <= 1; flappy_W(47, 120) <= 0; flappy_W(47, 121) <= 0; flappy_W(47, 122) <= 0; flappy_W(47, 123) <= 0; flappy_W(47, 124) <= 0; flappy_W(47, 125) <= 0; flappy_W(47, 126) <= 0; flappy_W(47, 127) <= 0; flappy_W(47, 128) <= 0; flappy_W(47, 129) <= 0; flappy_W(47, 130) <= 0; flappy_W(47, 131) <= 0; flappy_W(47, 132) <= 0; flappy_W(47, 133) <= 0; flappy_W(47, 134) <= 0; flappy_W(47, 135) <= 0; flappy_W(47, 136) <= 0; flappy_W(47, 137) <= 0; flappy_W(47, 138) <= 1; flappy_W(47, 139) <= 1; flappy_W(47, 140) <= 1; flappy_W(47, 141) <= 1; flappy_W(47, 142) <= 1; flappy_W(47, 143) <= 1; flappy_W(47, 144) <= 1; flappy_W(47, 145) <= 1; flappy_W(47, 146) <= 1; flappy_W(47, 147) <= 1; flappy_W(47, 148) <= 1; flappy_W(47, 149) <= 1; flappy_W(47, 150) <= 0; flappy_W(47, 151) <= 0; flappy_W(47, 152) <= 0; flappy_W(47, 153) <= 0; flappy_W(47, 154) <= 0; flappy_W(47, 155) <= 0; flappy_W(47, 156) <= 0; flappy_W(47, 157) <= 0; flappy_W(47, 158) <= 0; flappy_W(47, 159) <= 0; flappy_W(47, 160) <= 0; flappy_W(47, 161) <= 0; flappy_W(47, 162) <= 0; flappy_W(47, 163) <= 0; flappy_W(47, 164) <= 0; flappy_W(47, 165) <= 0; flappy_W(47, 166) <= 0; flappy_W(47, 167) <= 0; flappy_W(47, 168) <= 1; flappy_W(47, 169) <= 1; flappy_W(47, 170) <= 1; flappy_W(47, 171) <= 1; flappy_W(47, 172) <= 1; flappy_W(47, 173) <= 1; flappy_W(47, 174) <= 1; flappy_W(47, 175) <= 1; flappy_W(47, 176) <= 1; flappy_W(47, 177) <= 1; flappy_W(47, 178) <= 1; flappy_W(47, 179) <= 1; flappy_W(47, 180) <= 0; flappy_W(47, 181) <= 0; flappy_W(47, 182) <= 0; flappy_W(47, 183) <= 0; flappy_W(47, 184) <= 0; flappy_W(47, 185) <= 0; flappy_W(47, 186) <= 0; flappy_W(47, 187) <= 0; flappy_W(47, 188) <= 0; flappy_W(47, 189) <= 0; flappy_W(47, 190) <= 0; flappy_W(47, 191) <= 0; flappy_W(47, 192) <= 0; flappy_W(47, 193) <= 0; flappy_W(47, 194) <= 0; flappy_W(47, 195) <= 0; flappy_W(47, 196) <= 0; flappy_W(47, 197) <= 0; flappy_W(47, 198) <= 0; flappy_W(47, 199) <= 0; flappy_W(47, 200) <= 0; flappy_W(47, 201) <= 0; flappy_W(47, 202) <= 0; flappy_W(47, 203) <= 0; flappy_W(47, 204) <= 0; flappy_W(47, 205) <= 0; flappy_W(47, 206) <= 0; flappy_W(47, 207) <= 0; flappy_W(47, 208) <= 0; flappy_W(47, 209) <= 0; flappy_W(47, 210) <= 0; flappy_W(47, 211) <= 0; flappy_W(47, 212) <= 0; flappy_W(47, 213) <= 0; flappy_W(47, 214) <= 0; flappy_W(47, 215) <= 0; flappy_W(47, 216) <= 0; flappy_W(47, 217) <= 0; flappy_W(47, 218) <= 0; flappy_W(47, 219) <= 0; flappy_W(47, 220) <= 0; flappy_W(47, 221) <= 0; flappy_W(47, 222) <= 1; flappy_W(47, 223) <= 1; flappy_W(47, 224) <= 1; flappy_W(47, 225) <= 1; flappy_W(47, 226) <= 1; flappy_W(47, 227) <= 1; flappy_W(47, 228) <= 1; flappy_W(47, 229) <= 1; flappy_W(47, 230) <= 1; flappy_W(47, 231) <= 1; flappy_W(47, 232) <= 1; flappy_W(47, 233) <= 1; flappy_W(47, 234) <= 0; flappy_W(47, 235) <= 0; flappy_W(47, 236) <= 0; flappy_W(47, 237) <= 0; flappy_W(47, 238) <= 0; flappy_W(47, 239) <= 0; flappy_W(47, 240) <= 0; flappy_W(47, 241) <= 0; flappy_W(47, 242) <= 0; flappy_W(47, 243) <= 0; flappy_W(47, 244) <= 0; flappy_W(47, 245) <= 0; flappy_W(47, 246) <= 0; flappy_W(47, 247) <= 0; flappy_W(47, 248) <= 0; flappy_W(47, 249) <= 0; flappy_W(47, 250) <= 0; flappy_W(47, 251) <= 0; flappy_W(47, 252) <= 0; flappy_W(47, 253) <= 0; flappy_W(47, 254) <= 0; flappy_W(47, 255) <= 0; flappy_W(47, 256) <= 0; flappy_W(47, 257) <= 0; flappy_W(47, 258) <= 0; flappy_W(47, 259) <= 0; flappy_W(47, 260) <= 0; flappy_W(47, 261) <= 0; flappy_W(47, 262) <= 0; flappy_W(47, 263) <= 0; flappy_W(47, 264) <= 0; flappy_W(47, 265) <= 0; flappy_W(47, 266) <= 0; flappy_W(47, 267) <= 0; flappy_W(47, 268) <= 0; flappy_W(47, 269) <= 0; flappy_W(47, 270) <= 0; flappy_W(47, 271) <= 0; flappy_W(47, 272) <= 0; flappy_W(47, 273) <= 0; flappy_W(47, 274) <= 0; flappy_W(47, 275) <= 0; flappy_W(47, 276) <= 0; flappy_W(47, 277) <= 0; flappy_W(47, 278) <= 0; flappy_W(47, 279) <= 0; flappy_W(47, 280) <= 0; flappy_W(47, 281) <= 0; flappy_W(47, 282) <= 0; flappy_W(47, 283) <= 0; flappy_W(47, 284) <= 0; flappy_W(47, 285) <= 0; flappy_W(47, 286) <= 0; flappy_W(47, 287) <= 0; flappy_W(47, 288) <= 1; flappy_W(47, 289) <= 1; flappy_W(47, 290) <= 1; flappy_W(47, 291) <= 1; flappy_W(47, 292) <= 1; flappy_W(47, 293) <= 1; flappy_W(47, 294) <= 1; flappy_W(47, 295) <= 1; flappy_W(47, 296) <= 1; flappy_W(47, 297) <= 1; flappy_W(47, 298) <= 1; flappy_W(47, 299) <= 1; flappy_W(47, 300) <= 0; flappy_W(47, 301) <= 0; flappy_W(47, 302) <= 0; flappy_W(47, 303) <= 0; flappy_W(47, 304) <= 0; flappy_W(47, 305) <= 0; flappy_W(47, 306) <= 0; flappy_W(47, 307) <= 0; flappy_W(47, 308) <= 0; flappy_W(47, 309) <= 0; flappy_W(47, 310) <= 0; flappy_W(47, 311) <= 0; flappy_W(47, 312) <= 0; flappy_W(47, 313) <= 0; flappy_W(47, 314) <= 0; flappy_W(47, 315) <= 0; flappy_W(47, 316) <= 0; flappy_W(47, 317) <= 0; flappy_W(47, 318) <= 0; flappy_W(47, 319) <= 0; flappy_W(47, 320) <= 0; flappy_W(47, 321) <= 0; flappy_W(47, 322) <= 0; flappy_W(47, 323) <= 0; flappy_W(47, 324) <= 0; flappy_W(47, 325) <= 0; flappy_W(47, 326) <= 0; flappy_W(47, 327) <= 0; flappy_W(47, 328) <= 0; flappy_W(47, 329) <= 0; flappy_W(47, 330) <= 0; flappy_W(47, 331) <= 0; flappy_W(47, 332) <= 0; flappy_W(47, 333) <= 0; flappy_W(47, 334) <= 0; flappy_W(47, 335) <= 0; flappy_W(47, 336) <= 0; flappy_W(47, 337) <= 0; flappy_W(47, 338) <= 0; flappy_W(47, 339) <= 0; flappy_W(47, 340) <= 0; flappy_W(47, 341) <= 0; flappy_W(47, 342) <= 0; flappy_W(47, 343) <= 0; flappy_W(47, 344) <= 0; flappy_W(47, 345) <= 0; flappy_W(47, 346) <= 0; flappy_W(47, 347) <= 0; flappy_W(47, 348) <= 0; flappy_W(47, 349) <= 0; flappy_W(47, 350) <= 0; flappy_W(47, 351) <= 0; flappy_W(47, 352) <= 0; flappy_W(47, 353) <= 0; flappy_W(47, 354) <= 0; flappy_W(47, 355) <= 0; flappy_W(47, 356) <= 0; flappy_W(47, 357) <= 0; flappy_W(47, 358) <= 0; flappy_W(47, 359) <= 0; flappy_W(47, 360) <= 0; flappy_W(47, 361) <= 0; flappy_W(47, 362) <= 0; flappy_W(47, 363) <= 0; flappy_W(47, 364) <= 0; flappy_W(47, 365) <= 0; flappy_W(47, 366) <= 0; flappy_W(47, 367) <= 0; flappy_W(47, 368) <= 0; flappy_W(47, 369) <= 0; flappy_W(47, 370) <= 0; flappy_W(47, 371) <= 0; flappy_W(47, 372) <= 0; flappy_W(47, 373) <= 0; flappy_W(47, 374) <= 0; flappy_W(47, 375) <= 0; flappy_W(47, 376) <= 0; flappy_W(47, 377) <= 0; flappy_W(47, 378) <= 0; flappy_W(47, 379) <= 0; flappy_W(47, 380) <= 0; flappy_W(47, 381) <= 0; flappy_W(47, 382) <= 0; flappy_W(47, 383) <= 0; flappy_W(47, 384) <= 0; flappy_W(47, 385) <= 0; flappy_W(47, 386) <= 0; flappy_W(47, 387) <= 0; flappy_W(47, 388) <= 0; flappy_W(47, 389) <= 0; flappy_W(47, 390) <= 0; flappy_W(47, 391) <= 0; flappy_W(47, 392) <= 0; flappy_W(47, 393) <= 0; flappy_W(47, 394) <= 0; flappy_W(47, 395) <= 0; flappy_W(47, 396) <= 0; flappy_W(47, 397) <= 0; flappy_W(47, 398) <= 0; flappy_W(47, 399) <= 0; flappy_W(47, 400) <= 0; flappy_W(47, 401) <= 0; flappy_W(47, 402) <= 1; flappy_W(47, 403) <= 1; flappy_W(47, 404) <= 1; flappy_W(47, 405) <= 1; flappy_W(47, 406) <= 1; flappy_W(47, 407) <= 1; flappy_W(47, 408) <= 1; flappy_W(47, 409) <= 1; flappy_W(47, 410) <= 1; flappy_W(47, 411) <= 1; flappy_W(47, 412) <= 1; flappy_W(47, 413) <= 1; flappy_W(47, 414) <= 0; flappy_W(47, 415) <= 0; flappy_W(47, 416) <= 0; flappy_W(47, 417) <= 0; flappy_W(47, 418) <= 0; flappy_W(47, 419) <= 0; flappy_W(47, 420) <= 0; flappy_W(47, 421) <= 0; flappy_W(47, 422) <= 0; flappy_W(47, 423) <= 0; flappy_W(47, 424) <= 0; flappy_W(47, 425) <= 0; flappy_W(47, 426) <= 1; flappy_W(47, 427) <= 1; flappy_W(47, 428) <= 1; flappy_W(47, 429) <= 1; flappy_W(47, 430) <= 1; flappy_W(47, 431) <= 1; flappy_W(47, 432) <= 1; flappy_W(47, 433) <= 1; flappy_W(47, 434) <= 1; flappy_W(47, 435) <= 1; flappy_W(47, 436) <= 1; flappy_W(47, 437) <= 1; flappy_W(47, 438) <= 0; flappy_W(47, 439) <= 0; flappy_W(47, 440) <= 0; flappy_W(47, 441) <= 0; flappy_W(47, 442) <= 0; flappy_W(47, 443) <= 0; flappy_W(47, 444) <= 0; flappy_W(47, 445) <= 0; flappy_W(47, 446) <= 0; flappy_W(47, 447) <= 0; flappy_W(47, 448) <= 0; flappy_W(47, 449) <= 0; flappy_W(47, 450) <= 0; flappy_W(47, 451) <= 0; flappy_W(47, 452) <= 0; flappy_W(47, 453) <= 0; flappy_W(47, 454) <= 0; flappy_W(47, 455) <= 0; flappy_W(47, 456) <= 0; flappy_W(47, 457) <= 0; flappy_W(47, 458) <= 0; flappy_W(47, 459) <= 0; flappy_W(47, 460) <= 0; flappy_W(47, 461) <= 0; flappy_W(47, 462) <= 0; flappy_W(47, 463) <= 0; flappy_W(47, 464) <= 0; flappy_W(47, 465) <= 0; flappy_W(47, 466) <= 0; flappy_W(47, 467) <= 0; flappy_W(47, 468) <= 1; flappy_W(47, 469) <= 1; flappy_W(47, 470) <= 1; flappy_W(47, 471) <= 1; flappy_W(47, 472) <= 1; flappy_W(47, 473) <= 1; flappy_W(47, 474) <= 1; flappy_W(47, 475) <= 1; flappy_W(47, 476) <= 1; flappy_W(47, 477) <= 1; flappy_W(47, 478) <= 1; flappy_W(47, 479) <= 1; flappy_W(47, 480) <= 0; flappy_W(47, 481) <= 0; flappy_W(47, 482) <= 0; flappy_W(47, 483) <= 0; flappy_W(47, 484) <= 0; flappy_W(47, 485) <= 0; flappy_W(47, 486) <= 0; flappy_W(47, 487) <= 0; flappy_W(47, 488) <= 0; flappy_W(47, 489) <= 0; flappy_W(47, 490) <= 0; flappy_W(47, 491) <= 0; flappy_W(47, 492) <= 0; flappy_W(47, 493) <= 0; flappy_W(47, 494) <= 0; flappy_W(47, 495) <= 0; flappy_W(47, 496) <= 0; flappy_W(47, 497) <= 0; flappy_W(47, 498) <= 0; flappy_W(47, 499) <= 0; flappy_W(47, 500) <= 0; flappy_W(47, 501) <= 0; flappy_W(47, 502) <= 0; flappy_W(47, 503) <= 0; flappy_W(47, 504) <= 0; flappy_W(47, 505) <= 0; flappy_W(47, 506) <= 0; flappy_W(47, 507) <= 0; flappy_W(47, 508) <= 0; flappy_W(47, 509) <= 0; flappy_W(47, 510) <= 1; flappy_W(47, 511) <= 1; flappy_W(47, 512) <= 1; flappy_W(47, 513) <= 1; flappy_W(47, 514) <= 1; flappy_W(47, 515) <= 1; flappy_W(47, 516) <= 1; flappy_W(47, 517) <= 1; flappy_W(47, 518) <= 1; flappy_W(47, 519) <= 1; flappy_W(47, 520) <= 1; flappy_W(47, 521) <= 1; flappy_W(47, 522) <= 0; flappy_W(47, 523) <= 0; flappy_W(47, 524) <= 0; flappy_W(47, 525) <= 0; flappy_W(47, 526) <= 0; flappy_W(47, 527) <= 0; flappy_W(47, 528) <= 0; flappy_W(47, 529) <= 0; flappy_W(47, 530) <= 0; flappy_W(47, 531) <= 0; flappy_W(47, 532) <= 0; flappy_W(47, 533) <= 0; flappy_W(47, 534) <= 1; flappy_W(47, 535) <= 1; flappy_W(47, 536) <= 1; flappy_W(47, 537) <= 1; flappy_W(47, 538) <= 1; flappy_W(47, 539) <= 1; flappy_W(47, 540) <= 1; flappy_W(47, 541) <= 1; flappy_W(47, 542) <= 1; flappy_W(47, 543) <= 1; flappy_W(47, 544) <= 1; flappy_W(47, 545) <= 1; flappy_W(47, 546) <= 0; flappy_W(47, 547) <= 0; flappy_W(47, 548) <= 0; flappy_W(47, 549) <= 0; flappy_W(47, 550) <= 0; flappy_W(47, 551) <= 0; flappy_W(47, 552) <= 0; flappy_W(47, 553) <= 0; flappy_W(47, 554) <= 0; flappy_W(47, 555) <= 0; flappy_W(47, 556) <= 0; flappy_W(47, 557) <= 0; flappy_W(47, 558) <= 0; flappy_W(47, 559) <= 0; flappy_W(47, 560) <= 0; flappy_W(47, 561) <= 0; flappy_W(47, 562) <= 0; flappy_W(47, 563) <= 0; flappy_W(47, 564) <= 1; flappy_W(47, 565) <= 1; flappy_W(47, 566) <= 1; flappy_W(47, 567) <= 1; flappy_W(47, 568) <= 1; flappy_W(47, 569) <= 1; flappy_W(47, 570) <= 1; flappy_W(47, 571) <= 1; flappy_W(47, 572) <= 1; flappy_W(47, 573) <= 1; flappy_W(47, 574) <= 1; flappy_W(47, 575) <= 1; flappy_W(47, 576) <= 0; flappy_W(47, 577) <= 0; flappy_W(47, 578) <= 0; flappy_W(47, 579) <= 0; flappy_W(47, 580) <= 0; flappy_W(47, 581) <= 0; flappy_W(47, 582) <= 0; flappy_W(47, 583) <= 0; flappy_W(47, 584) <= 0; flappy_W(47, 585) <= 0; flappy_W(47, 586) <= 0; flappy_W(47, 587) <= 0; flappy_W(47, 588) <= 1; flappy_W(47, 589) <= 1; flappy_W(47, 590) <= 1; flappy_W(47, 591) <= 1; flappy_W(47, 592) <= 1; flappy_W(47, 593) <= 1; 
flappy_W(48, 0) <= 0; flappy_W(48, 1) <= 0; flappy_W(48, 2) <= 0; flappy_W(48, 3) <= 0; flappy_W(48, 4) <= 0; flappy_W(48, 5) <= 0; flappy_W(48, 6) <= 1; flappy_W(48, 7) <= 1; flappy_W(48, 8) <= 1; flappy_W(48, 9) <= 1; flappy_W(48, 10) <= 1; flappy_W(48, 11) <= 1; flappy_W(48, 12) <= 1; flappy_W(48, 13) <= 1; flappy_W(48, 14) <= 1; flappy_W(48, 15) <= 1; flappy_W(48, 16) <= 1; flappy_W(48, 17) <= 1; flappy_W(48, 18) <= 0; flappy_W(48, 19) <= 0; flappy_W(48, 20) <= 0; flappy_W(48, 21) <= 0; flappy_W(48, 22) <= 0; flappy_W(48, 23) <= 0; flappy_W(48, 24) <= 0; flappy_W(48, 25) <= 0; flappy_W(48, 26) <= 0; flappy_W(48, 27) <= 0; flappy_W(48, 28) <= 0; flappy_W(48, 29) <= 0; flappy_W(48, 30) <= 0; flappy_W(48, 31) <= 0; flappy_W(48, 32) <= 0; flappy_W(48, 33) <= 0; flappy_W(48, 34) <= 0; flappy_W(48, 35) <= 0; flappy_W(48, 36) <= 0; flappy_W(48, 37) <= 0; flappy_W(48, 38) <= 0; flappy_W(48, 39) <= 0; flappy_W(48, 40) <= 0; flappy_W(48, 41) <= 0; flappy_W(48, 42) <= 0; flappy_W(48, 43) <= 0; flappy_W(48, 44) <= 0; flappy_W(48, 45) <= 0; flappy_W(48, 46) <= 0; flappy_W(48, 47) <= 0; flappy_W(48, 48) <= 0; flappy_W(48, 49) <= 0; flappy_W(48, 50) <= 0; flappy_W(48, 51) <= 0; flappy_W(48, 52) <= 0; flappy_W(48, 53) <= 0; flappy_W(48, 54) <= 0; flappy_W(48, 55) <= 0; flappy_W(48, 56) <= 0; flappy_W(48, 57) <= 0; flappy_W(48, 58) <= 0; flappy_W(48, 59) <= 0; flappy_W(48, 60) <= 1; flappy_W(48, 61) <= 1; flappy_W(48, 62) <= 1; flappy_W(48, 63) <= 1; flappy_W(48, 64) <= 1; flappy_W(48, 65) <= 1; flappy_W(48, 66) <= 1; flappy_W(48, 67) <= 1; flappy_W(48, 68) <= 1; flappy_W(48, 69) <= 1; flappy_W(48, 70) <= 1; flappy_W(48, 71) <= 1; flappy_W(48, 72) <= 0; flappy_W(48, 73) <= 0; flappy_W(48, 74) <= 0; flappy_W(48, 75) <= 0; flappy_W(48, 76) <= 0; flappy_W(48, 77) <= 0; flappy_W(48, 78) <= 0; flappy_W(48, 79) <= 0; flappy_W(48, 80) <= 0; flappy_W(48, 81) <= 0; flappy_W(48, 82) <= 0; flappy_W(48, 83) <= 0; flappy_W(48, 84) <= 1; flappy_W(48, 85) <= 1; flappy_W(48, 86) <= 1; flappy_W(48, 87) <= 1; flappy_W(48, 88) <= 1; flappy_W(48, 89) <= 1; flappy_W(48, 90) <= 1; flappy_W(48, 91) <= 1; flappy_W(48, 92) <= 1; flappy_W(48, 93) <= 1; flappy_W(48, 94) <= 1; flappy_W(48, 95) <= 1; flappy_W(48, 96) <= 0; flappy_W(48, 97) <= 0; flappy_W(48, 98) <= 0; flappy_W(48, 99) <= 0; flappy_W(48, 100) <= 0; flappy_W(48, 101) <= 0; flappy_W(48, 102) <= 0; flappy_W(48, 103) <= 0; flappy_W(48, 104) <= 0; flappy_W(48, 105) <= 0; flappy_W(48, 106) <= 0; flappy_W(48, 107) <= 0; flappy_W(48, 108) <= 1; flappy_W(48, 109) <= 1; flappy_W(48, 110) <= 1; flappy_W(48, 111) <= 1; flappy_W(48, 112) <= 1; flappy_W(48, 113) <= 1; flappy_W(48, 114) <= 1; flappy_W(48, 115) <= 1; flappy_W(48, 116) <= 1; flappy_W(48, 117) <= 1; flappy_W(48, 118) <= 1; flappy_W(48, 119) <= 1; flappy_W(48, 120) <= 0; flappy_W(48, 121) <= 0; flappy_W(48, 122) <= 0; flappy_W(48, 123) <= 0; flappy_W(48, 124) <= 0; flappy_W(48, 125) <= 0; flappy_W(48, 126) <= 0; flappy_W(48, 127) <= 0; flappy_W(48, 128) <= 0; flappy_W(48, 129) <= 0; flappy_W(48, 130) <= 0; flappy_W(48, 131) <= 0; flappy_W(48, 132) <= 0; flappy_W(48, 133) <= 0; flappy_W(48, 134) <= 0; flappy_W(48, 135) <= 0; flappy_W(48, 136) <= 0; flappy_W(48, 137) <= 0; flappy_W(48, 138) <= 1; flappy_W(48, 139) <= 1; flappy_W(48, 140) <= 1; flappy_W(48, 141) <= 1; flappy_W(48, 142) <= 1; flappy_W(48, 143) <= 1; flappy_W(48, 144) <= 1; flappy_W(48, 145) <= 1; flappy_W(48, 146) <= 1; flappy_W(48, 147) <= 1; flappy_W(48, 148) <= 1; flappy_W(48, 149) <= 1; flappy_W(48, 150) <= 0; flappy_W(48, 151) <= 0; flappy_W(48, 152) <= 0; flappy_W(48, 153) <= 0; flappy_W(48, 154) <= 0; flappy_W(48, 155) <= 0; flappy_W(48, 156) <= 0; flappy_W(48, 157) <= 0; flappy_W(48, 158) <= 0; flappy_W(48, 159) <= 0; flappy_W(48, 160) <= 0; flappy_W(48, 161) <= 0; flappy_W(48, 162) <= 0; flappy_W(48, 163) <= 0; flappy_W(48, 164) <= 0; flappy_W(48, 165) <= 0; flappy_W(48, 166) <= 0; flappy_W(48, 167) <= 0; flappy_W(48, 168) <= 1; flappy_W(48, 169) <= 1; flappy_W(48, 170) <= 1; flappy_W(48, 171) <= 1; flappy_W(48, 172) <= 1; flappy_W(48, 173) <= 1; flappy_W(48, 174) <= 1; flappy_W(48, 175) <= 1; flappy_W(48, 176) <= 1; flappy_W(48, 177) <= 1; flappy_W(48, 178) <= 1; flappy_W(48, 179) <= 1; flappy_W(48, 180) <= 0; flappy_W(48, 181) <= 0; flappy_W(48, 182) <= 0; flappy_W(48, 183) <= 0; flappy_W(48, 184) <= 0; flappy_W(48, 185) <= 0; flappy_W(48, 186) <= 0; flappy_W(48, 187) <= 0; flappy_W(48, 188) <= 0; flappy_W(48, 189) <= 0; flappy_W(48, 190) <= 0; flappy_W(48, 191) <= 0; flappy_W(48, 192) <= 0; flappy_W(48, 193) <= 0; flappy_W(48, 194) <= 0; flappy_W(48, 195) <= 0; flappy_W(48, 196) <= 0; flappy_W(48, 197) <= 0; flappy_W(48, 198) <= 0; flappy_W(48, 199) <= 0; flappy_W(48, 200) <= 0; flappy_W(48, 201) <= 0; flappy_W(48, 202) <= 0; flappy_W(48, 203) <= 0; flappy_W(48, 204) <= 0; flappy_W(48, 205) <= 0; flappy_W(48, 206) <= 0; flappy_W(48, 207) <= 0; flappy_W(48, 208) <= 0; flappy_W(48, 209) <= 0; flappy_W(48, 210) <= 0; flappy_W(48, 211) <= 0; flappy_W(48, 212) <= 0; flappy_W(48, 213) <= 0; flappy_W(48, 214) <= 0; flappy_W(48, 215) <= 0; flappy_W(48, 216) <= 0; flappy_W(48, 217) <= 0; flappy_W(48, 218) <= 0; flappy_W(48, 219) <= 0; flappy_W(48, 220) <= 0; flappy_W(48, 221) <= 0; flappy_W(48, 222) <= 1; flappy_W(48, 223) <= 1; flappy_W(48, 224) <= 1; flappy_W(48, 225) <= 1; flappy_W(48, 226) <= 1; flappy_W(48, 227) <= 1; flappy_W(48, 228) <= 1; flappy_W(48, 229) <= 1; flappy_W(48, 230) <= 1; flappy_W(48, 231) <= 1; flappy_W(48, 232) <= 1; flappy_W(48, 233) <= 1; flappy_W(48, 234) <= 0; flappy_W(48, 235) <= 0; flappy_W(48, 236) <= 0; flappy_W(48, 237) <= 0; flappy_W(48, 238) <= 0; flappy_W(48, 239) <= 0; flappy_W(48, 240) <= 0; flappy_W(48, 241) <= 0; flappy_W(48, 242) <= 0; flappy_W(48, 243) <= 0; flappy_W(48, 244) <= 0; flappy_W(48, 245) <= 0; flappy_W(48, 246) <= 0; flappy_W(48, 247) <= 0; flappy_W(48, 248) <= 0; flappy_W(48, 249) <= 0; flappy_W(48, 250) <= 0; flappy_W(48, 251) <= 0; flappy_W(48, 252) <= 0; flappy_W(48, 253) <= 0; flappy_W(48, 254) <= 0; flappy_W(48, 255) <= 0; flappy_W(48, 256) <= 0; flappy_W(48, 257) <= 0; flappy_W(48, 258) <= 0; flappy_W(48, 259) <= 0; flappy_W(48, 260) <= 0; flappy_W(48, 261) <= 0; flappy_W(48, 262) <= 0; flappy_W(48, 263) <= 0; flappy_W(48, 264) <= 0; flappy_W(48, 265) <= 0; flappy_W(48, 266) <= 0; flappy_W(48, 267) <= 0; flappy_W(48, 268) <= 0; flappy_W(48, 269) <= 0; flappy_W(48, 270) <= 0; flappy_W(48, 271) <= 0; flappy_W(48, 272) <= 0; flappy_W(48, 273) <= 0; flappy_W(48, 274) <= 0; flappy_W(48, 275) <= 0; flappy_W(48, 276) <= 0; flappy_W(48, 277) <= 0; flappy_W(48, 278) <= 0; flappy_W(48, 279) <= 0; flappy_W(48, 280) <= 0; flappy_W(48, 281) <= 0; flappy_W(48, 282) <= 0; flappy_W(48, 283) <= 0; flappy_W(48, 284) <= 0; flappy_W(48, 285) <= 0; flappy_W(48, 286) <= 0; flappy_W(48, 287) <= 0; flappy_W(48, 288) <= 1; flappy_W(48, 289) <= 1; flappy_W(48, 290) <= 1; flappy_W(48, 291) <= 1; flappy_W(48, 292) <= 1; flappy_W(48, 293) <= 1; flappy_W(48, 294) <= 1; flappy_W(48, 295) <= 1; flappy_W(48, 296) <= 1; flappy_W(48, 297) <= 1; flappy_W(48, 298) <= 1; flappy_W(48, 299) <= 1; flappy_W(48, 300) <= 0; flappy_W(48, 301) <= 0; flappy_W(48, 302) <= 0; flappy_W(48, 303) <= 0; flappy_W(48, 304) <= 0; flappy_W(48, 305) <= 0; flappy_W(48, 306) <= 0; flappy_W(48, 307) <= 0; flappy_W(48, 308) <= 0; flappy_W(48, 309) <= 0; flappy_W(48, 310) <= 0; flappy_W(48, 311) <= 0; flappy_W(48, 312) <= 0; flappy_W(48, 313) <= 0; flappy_W(48, 314) <= 0; flappy_W(48, 315) <= 0; flappy_W(48, 316) <= 0; flappy_W(48, 317) <= 0; flappy_W(48, 318) <= 0; flappy_W(48, 319) <= 0; flappy_W(48, 320) <= 0; flappy_W(48, 321) <= 0; flappy_W(48, 322) <= 0; flappy_W(48, 323) <= 0; flappy_W(48, 324) <= 0; flappy_W(48, 325) <= 0; flappy_W(48, 326) <= 0; flappy_W(48, 327) <= 0; flappy_W(48, 328) <= 0; flappy_W(48, 329) <= 0; flappy_W(48, 330) <= 0; flappy_W(48, 331) <= 0; flappy_W(48, 332) <= 0; flappy_W(48, 333) <= 0; flappy_W(48, 334) <= 0; flappy_W(48, 335) <= 0; flappy_W(48, 336) <= 0; flappy_W(48, 337) <= 0; flappy_W(48, 338) <= 0; flappy_W(48, 339) <= 0; flappy_W(48, 340) <= 0; flappy_W(48, 341) <= 0; flappy_W(48, 342) <= 0; flappy_W(48, 343) <= 0; flappy_W(48, 344) <= 0; flappy_W(48, 345) <= 0; flappy_W(48, 346) <= 0; flappy_W(48, 347) <= 0; flappy_W(48, 348) <= 0; flappy_W(48, 349) <= 0; flappy_W(48, 350) <= 0; flappy_W(48, 351) <= 0; flappy_W(48, 352) <= 0; flappy_W(48, 353) <= 0; flappy_W(48, 354) <= 0; flappy_W(48, 355) <= 0; flappy_W(48, 356) <= 0; flappy_W(48, 357) <= 0; flappy_W(48, 358) <= 0; flappy_W(48, 359) <= 0; flappy_W(48, 360) <= 0; flappy_W(48, 361) <= 0; flappy_W(48, 362) <= 0; flappy_W(48, 363) <= 0; flappy_W(48, 364) <= 0; flappy_W(48, 365) <= 0; flappy_W(48, 366) <= 0; flappy_W(48, 367) <= 0; flappy_W(48, 368) <= 0; flappy_W(48, 369) <= 0; flappy_W(48, 370) <= 0; flappy_W(48, 371) <= 0; flappy_W(48, 372) <= 0; flappy_W(48, 373) <= 0; flappy_W(48, 374) <= 0; flappy_W(48, 375) <= 0; flappy_W(48, 376) <= 0; flappy_W(48, 377) <= 0; flappy_W(48, 378) <= 0; flappy_W(48, 379) <= 0; flappy_W(48, 380) <= 0; flappy_W(48, 381) <= 0; flappy_W(48, 382) <= 0; flappy_W(48, 383) <= 0; flappy_W(48, 384) <= 0; flappy_W(48, 385) <= 0; flappy_W(48, 386) <= 0; flappy_W(48, 387) <= 0; flappy_W(48, 388) <= 0; flappy_W(48, 389) <= 0; flappy_W(48, 390) <= 0; flappy_W(48, 391) <= 0; flappy_W(48, 392) <= 0; flappy_W(48, 393) <= 0; flappy_W(48, 394) <= 0; flappy_W(48, 395) <= 0; flappy_W(48, 396) <= 0; flappy_W(48, 397) <= 0; flappy_W(48, 398) <= 0; flappy_W(48, 399) <= 0; flappy_W(48, 400) <= 0; flappy_W(48, 401) <= 0; flappy_W(48, 402) <= 1; flappy_W(48, 403) <= 1; flappy_W(48, 404) <= 1; flappy_W(48, 405) <= 1; flappy_W(48, 406) <= 1; flappy_W(48, 407) <= 1; flappy_W(48, 408) <= 1; flappy_W(48, 409) <= 1; flappy_W(48, 410) <= 1; flappy_W(48, 411) <= 1; flappy_W(48, 412) <= 1; flappy_W(48, 413) <= 1; flappy_W(48, 414) <= 0; flappy_W(48, 415) <= 0; flappy_W(48, 416) <= 0; flappy_W(48, 417) <= 0; flappy_W(48, 418) <= 0; flappy_W(48, 419) <= 0; flappy_W(48, 420) <= 0; flappy_W(48, 421) <= 0; flappy_W(48, 422) <= 0; flappy_W(48, 423) <= 0; flappy_W(48, 424) <= 0; flappy_W(48, 425) <= 0; flappy_W(48, 426) <= 1; flappy_W(48, 427) <= 1; flappy_W(48, 428) <= 1; flappy_W(48, 429) <= 1; flappy_W(48, 430) <= 1; flappy_W(48, 431) <= 1; flappy_W(48, 432) <= 1; flappy_W(48, 433) <= 1; flappy_W(48, 434) <= 1; flappy_W(48, 435) <= 1; flappy_W(48, 436) <= 1; flappy_W(48, 437) <= 1; flappy_W(48, 438) <= 0; flappy_W(48, 439) <= 0; flappy_W(48, 440) <= 0; flappy_W(48, 441) <= 0; flappy_W(48, 442) <= 0; flappy_W(48, 443) <= 0; flappy_W(48, 444) <= 0; flappy_W(48, 445) <= 0; flappy_W(48, 446) <= 0; flappy_W(48, 447) <= 0; flappy_W(48, 448) <= 0; flappy_W(48, 449) <= 0; flappy_W(48, 450) <= 0; flappy_W(48, 451) <= 0; flappy_W(48, 452) <= 0; flappy_W(48, 453) <= 0; flappy_W(48, 454) <= 0; flappy_W(48, 455) <= 0; flappy_W(48, 456) <= 0; flappy_W(48, 457) <= 0; flappy_W(48, 458) <= 0; flappy_W(48, 459) <= 0; flappy_W(48, 460) <= 0; flappy_W(48, 461) <= 0; flappy_W(48, 462) <= 0; flappy_W(48, 463) <= 0; flappy_W(48, 464) <= 0; flappy_W(48, 465) <= 0; flappy_W(48, 466) <= 0; flappy_W(48, 467) <= 0; flappy_W(48, 468) <= 1; flappy_W(48, 469) <= 1; flappy_W(48, 470) <= 1; flappy_W(48, 471) <= 1; flappy_W(48, 472) <= 1; flappy_W(48, 473) <= 1; flappy_W(48, 474) <= 1; flappy_W(48, 475) <= 1; flappy_W(48, 476) <= 1; flappy_W(48, 477) <= 1; flappy_W(48, 478) <= 1; flappy_W(48, 479) <= 1; flappy_W(48, 480) <= 0; flappy_W(48, 481) <= 0; flappy_W(48, 482) <= 0; flappy_W(48, 483) <= 0; flappy_W(48, 484) <= 0; flappy_W(48, 485) <= 0; flappy_W(48, 486) <= 0; flappy_W(48, 487) <= 0; flappy_W(48, 488) <= 0; flappy_W(48, 489) <= 0; flappy_W(48, 490) <= 0; flappy_W(48, 491) <= 0; flappy_W(48, 492) <= 0; flappy_W(48, 493) <= 0; flappy_W(48, 494) <= 0; flappy_W(48, 495) <= 0; flappy_W(48, 496) <= 0; flappy_W(48, 497) <= 0; flappy_W(48, 498) <= 0; flappy_W(48, 499) <= 0; flappy_W(48, 500) <= 0; flappy_W(48, 501) <= 0; flappy_W(48, 502) <= 0; flappy_W(48, 503) <= 0; flappy_W(48, 504) <= 0; flappy_W(48, 505) <= 0; flappy_W(48, 506) <= 0; flappy_W(48, 507) <= 0; flappy_W(48, 508) <= 0; flappy_W(48, 509) <= 0; flappy_W(48, 510) <= 1; flappy_W(48, 511) <= 1; flappy_W(48, 512) <= 1; flappy_W(48, 513) <= 1; flappy_W(48, 514) <= 1; flappy_W(48, 515) <= 1; flappy_W(48, 516) <= 1; flappy_W(48, 517) <= 1; flappy_W(48, 518) <= 1; flappy_W(48, 519) <= 1; flappy_W(48, 520) <= 1; flappy_W(48, 521) <= 1; flappy_W(48, 522) <= 0; flappy_W(48, 523) <= 0; flappy_W(48, 524) <= 0; flappy_W(48, 525) <= 0; flappy_W(48, 526) <= 0; flappy_W(48, 527) <= 0; flappy_W(48, 528) <= 0; flappy_W(48, 529) <= 0; flappy_W(48, 530) <= 0; flappy_W(48, 531) <= 0; flappy_W(48, 532) <= 0; flappy_W(48, 533) <= 0; flappy_W(48, 534) <= 1; flappy_W(48, 535) <= 1; flappy_W(48, 536) <= 1; flappy_W(48, 537) <= 1; flappy_W(48, 538) <= 1; flappy_W(48, 539) <= 1; flappy_W(48, 540) <= 1; flappy_W(48, 541) <= 1; flappy_W(48, 542) <= 1; flappy_W(48, 543) <= 1; flappy_W(48, 544) <= 1; flappy_W(48, 545) <= 1; flappy_W(48, 546) <= 0; flappy_W(48, 547) <= 0; flappy_W(48, 548) <= 0; flappy_W(48, 549) <= 0; flappy_W(48, 550) <= 0; flappy_W(48, 551) <= 0; flappy_W(48, 552) <= 0; flappy_W(48, 553) <= 0; flappy_W(48, 554) <= 0; flappy_W(48, 555) <= 0; flappy_W(48, 556) <= 0; flappy_W(48, 557) <= 0; flappy_W(48, 558) <= 0; flappy_W(48, 559) <= 0; flappy_W(48, 560) <= 0; flappy_W(48, 561) <= 0; flappy_W(48, 562) <= 0; flappy_W(48, 563) <= 0; flappy_W(48, 564) <= 1; flappy_W(48, 565) <= 1; flappy_W(48, 566) <= 1; flappy_W(48, 567) <= 1; flappy_W(48, 568) <= 1; flappy_W(48, 569) <= 1; flappy_W(48, 570) <= 1; flappy_W(48, 571) <= 1; flappy_W(48, 572) <= 1; flappy_W(48, 573) <= 1; flappy_W(48, 574) <= 1; flappy_W(48, 575) <= 1; flappy_W(48, 576) <= 0; flappy_W(48, 577) <= 0; flappy_W(48, 578) <= 0; flappy_W(48, 579) <= 0; flappy_W(48, 580) <= 0; flappy_W(48, 581) <= 0; flappy_W(48, 582) <= 1; flappy_W(48, 583) <= 1; flappy_W(48, 584) <= 1; flappy_W(48, 585) <= 1; flappy_W(48, 586) <= 1; flappy_W(48, 587) <= 1; flappy_W(48, 588) <= 1; flappy_W(48, 589) <= 1; flappy_W(48, 590) <= 1; flappy_W(48, 591) <= 1; flappy_W(48, 592) <= 1; flappy_W(48, 593) <= 1; 
flappy_W(49, 0) <= 0; flappy_W(49, 1) <= 0; flappy_W(49, 2) <= 0; flappy_W(49, 3) <= 0; flappy_W(49, 4) <= 0; flappy_W(49, 5) <= 0; flappy_W(49, 6) <= 1; flappy_W(49, 7) <= 1; flappy_W(49, 8) <= 1; flappy_W(49, 9) <= 1; flappy_W(49, 10) <= 1; flappy_W(49, 11) <= 1; flappy_W(49, 12) <= 1; flappy_W(49, 13) <= 1; flappy_W(49, 14) <= 1; flappy_W(49, 15) <= 1; flappy_W(49, 16) <= 1; flappy_W(49, 17) <= 1; flappy_W(49, 18) <= 0; flappy_W(49, 19) <= 0; flappy_W(49, 20) <= 0; flappy_W(49, 21) <= 0; flappy_W(49, 22) <= 0; flappy_W(49, 23) <= 0; flappy_W(49, 24) <= 0; flappy_W(49, 25) <= 0; flappy_W(49, 26) <= 0; flappy_W(49, 27) <= 0; flappy_W(49, 28) <= 0; flappy_W(49, 29) <= 0; flappy_W(49, 30) <= 0; flappy_W(49, 31) <= 0; flappy_W(49, 32) <= 0; flappy_W(49, 33) <= 0; flappy_W(49, 34) <= 0; flappy_W(49, 35) <= 0; flappy_W(49, 36) <= 0; flappy_W(49, 37) <= 0; flappy_W(49, 38) <= 0; flappy_W(49, 39) <= 0; flappy_W(49, 40) <= 0; flappy_W(49, 41) <= 0; flappy_W(49, 42) <= 0; flappy_W(49, 43) <= 0; flappy_W(49, 44) <= 0; flappy_W(49, 45) <= 0; flappy_W(49, 46) <= 0; flappy_W(49, 47) <= 0; flappy_W(49, 48) <= 0; flappy_W(49, 49) <= 0; flappy_W(49, 50) <= 0; flappy_W(49, 51) <= 0; flappy_W(49, 52) <= 0; flappy_W(49, 53) <= 0; flappy_W(49, 54) <= 0; flappy_W(49, 55) <= 0; flappy_W(49, 56) <= 0; flappy_W(49, 57) <= 0; flappy_W(49, 58) <= 0; flappy_W(49, 59) <= 0; flappy_W(49, 60) <= 1; flappy_W(49, 61) <= 1; flappy_W(49, 62) <= 1; flappy_W(49, 63) <= 1; flappy_W(49, 64) <= 1; flappy_W(49, 65) <= 1; flappy_W(49, 66) <= 1; flappy_W(49, 67) <= 1; flappy_W(49, 68) <= 1; flappy_W(49, 69) <= 1; flappy_W(49, 70) <= 1; flappy_W(49, 71) <= 1; flappy_W(49, 72) <= 0; flappy_W(49, 73) <= 0; flappy_W(49, 74) <= 0; flappy_W(49, 75) <= 0; flappy_W(49, 76) <= 0; flappy_W(49, 77) <= 0; flappy_W(49, 78) <= 0; flappy_W(49, 79) <= 0; flappy_W(49, 80) <= 0; flappy_W(49, 81) <= 0; flappy_W(49, 82) <= 0; flappy_W(49, 83) <= 0; flappy_W(49, 84) <= 1; flappy_W(49, 85) <= 1; flappy_W(49, 86) <= 1; flappy_W(49, 87) <= 1; flappy_W(49, 88) <= 1; flappy_W(49, 89) <= 1; flappy_W(49, 90) <= 1; flappy_W(49, 91) <= 1; flappy_W(49, 92) <= 1; flappy_W(49, 93) <= 1; flappy_W(49, 94) <= 1; flappy_W(49, 95) <= 1; flappy_W(49, 96) <= 0; flappy_W(49, 97) <= 0; flappy_W(49, 98) <= 0; flappy_W(49, 99) <= 0; flappy_W(49, 100) <= 0; flappy_W(49, 101) <= 0; flappy_W(49, 102) <= 0; flappy_W(49, 103) <= 0; flappy_W(49, 104) <= 0; flappy_W(49, 105) <= 0; flappy_W(49, 106) <= 0; flappy_W(49, 107) <= 0; flappy_W(49, 108) <= 1; flappy_W(49, 109) <= 1; flappy_W(49, 110) <= 1; flappy_W(49, 111) <= 1; flappy_W(49, 112) <= 1; flappy_W(49, 113) <= 1; flappy_W(49, 114) <= 1; flappy_W(49, 115) <= 1; flappy_W(49, 116) <= 1; flappy_W(49, 117) <= 1; flappy_W(49, 118) <= 1; flappy_W(49, 119) <= 1; flappy_W(49, 120) <= 0; flappy_W(49, 121) <= 0; flappy_W(49, 122) <= 0; flappy_W(49, 123) <= 0; flappy_W(49, 124) <= 0; flappy_W(49, 125) <= 0; flappy_W(49, 126) <= 0; flappy_W(49, 127) <= 0; flappy_W(49, 128) <= 0; flappy_W(49, 129) <= 0; flappy_W(49, 130) <= 0; flappy_W(49, 131) <= 0; flappy_W(49, 132) <= 0; flappy_W(49, 133) <= 0; flappy_W(49, 134) <= 0; flappy_W(49, 135) <= 0; flappy_W(49, 136) <= 0; flappy_W(49, 137) <= 0; flappy_W(49, 138) <= 1; flappy_W(49, 139) <= 1; flappy_W(49, 140) <= 1; flappy_W(49, 141) <= 1; flappy_W(49, 142) <= 1; flappy_W(49, 143) <= 1; flappy_W(49, 144) <= 1; flappy_W(49, 145) <= 1; flappy_W(49, 146) <= 1; flappy_W(49, 147) <= 1; flappy_W(49, 148) <= 1; flappy_W(49, 149) <= 1; flappy_W(49, 150) <= 0; flappy_W(49, 151) <= 0; flappy_W(49, 152) <= 0; flappy_W(49, 153) <= 0; flappy_W(49, 154) <= 0; flappy_W(49, 155) <= 0; flappy_W(49, 156) <= 0; flappy_W(49, 157) <= 0; flappy_W(49, 158) <= 0; flappy_W(49, 159) <= 0; flappy_W(49, 160) <= 0; flappy_W(49, 161) <= 0; flappy_W(49, 162) <= 0; flappy_W(49, 163) <= 0; flappy_W(49, 164) <= 0; flappy_W(49, 165) <= 0; flappy_W(49, 166) <= 0; flappy_W(49, 167) <= 0; flappy_W(49, 168) <= 1; flappy_W(49, 169) <= 1; flappy_W(49, 170) <= 1; flappy_W(49, 171) <= 1; flappy_W(49, 172) <= 1; flappy_W(49, 173) <= 1; flappy_W(49, 174) <= 1; flappy_W(49, 175) <= 1; flappy_W(49, 176) <= 1; flappy_W(49, 177) <= 1; flappy_W(49, 178) <= 1; flappy_W(49, 179) <= 1; flappy_W(49, 180) <= 0; flappy_W(49, 181) <= 0; flappy_W(49, 182) <= 0; flappy_W(49, 183) <= 0; flappy_W(49, 184) <= 0; flappy_W(49, 185) <= 0; flappy_W(49, 186) <= 0; flappy_W(49, 187) <= 0; flappy_W(49, 188) <= 0; flappy_W(49, 189) <= 0; flappy_W(49, 190) <= 0; flappy_W(49, 191) <= 0; flappy_W(49, 192) <= 0; flappy_W(49, 193) <= 0; flappy_W(49, 194) <= 0; flappy_W(49, 195) <= 0; flappy_W(49, 196) <= 0; flappy_W(49, 197) <= 0; flappy_W(49, 198) <= 0; flappy_W(49, 199) <= 0; flappy_W(49, 200) <= 0; flappy_W(49, 201) <= 0; flappy_W(49, 202) <= 0; flappy_W(49, 203) <= 0; flappy_W(49, 204) <= 0; flappy_W(49, 205) <= 0; flappy_W(49, 206) <= 0; flappy_W(49, 207) <= 0; flappy_W(49, 208) <= 0; flappy_W(49, 209) <= 0; flappy_W(49, 210) <= 0; flappy_W(49, 211) <= 0; flappy_W(49, 212) <= 0; flappy_W(49, 213) <= 0; flappy_W(49, 214) <= 0; flappy_W(49, 215) <= 0; flappy_W(49, 216) <= 0; flappy_W(49, 217) <= 0; flappy_W(49, 218) <= 0; flappy_W(49, 219) <= 0; flappy_W(49, 220) <= 0; flappy_W(49, 221) <= 0; flappy_W(49, 222) <= 1; flappy_W(49, 223) <= 1; flappy_W(49, 224) <= 1; flappy_W(49, 225) <= 1; flappy_W(49, 226) <= 1; flappy_W(49, 227) <= 1; flappy_W(49, 228) <= 1; flappy_W(49, 229) <= 1; flappy_W(49, 230) <= 1; flappy_W(49, 231) <= 1; flappy_W(49, 232) <= 1; flappy_W(49, 233) <= 1; flappy_W(49, 234) <= 0; flappy_W(49, 235) <= 0; flappy_W(49, 236) <= 0; flappy_W(49, 237) <= 0; flappy_W(49, 238) <= 0; flappy_W(49, 239) <= 0; flappy_W(49, 240) <= 0; flappy_W(49, 241) <= 0; flappy_W(49, 242) <= 0; flappy_W(49, 243) <= 0; flappy_W(49, 244) <= 0; flappy_W(49, 245) <= 0; flappy_W(49, 246) <= 0; flappy_W(49, 247) <= 0; flappy_W(49, 248) <= 0; flappy_W(49, 249) <= 0; flappy_W(49, 250) <= 0; flappy_W(49, 251) <= 0; flappy_W(49, 252) <= 0; flappy_W(49, 253) <= 0; flappy_W(49, 254) <= 0; flappy_W(49, 255) <= 0; flappy_W(49, 256) <= 0; flappy_W(49, 257) <= 0; flappy_W(49, 258) <= 0; flappy_W(49, 259) <= 0; flappy_W(49, 260) <= 0; flappy_W(49, 261) <= 0; flappy_W(49, 262) <= 0; flappy_W(49, 263) <= 0; flappy_W(49, 264) <= 0; flappy_W(49, 265) <= 0; flappy_W(49, 266) <= 0; flappy_W(49, 267) <= 0; flappy_W(49, 268) <= 0; flappy_W(49, 269) <= 0; flappy_W(49, 270) <= 0; flappy_W(49, 271) <= 0; flappy_W(49, 272) <= 0; flappy_W(49, 273) <= 0; flappy_W(49, 274) <= 0; flappy_W(49, 275) <= 0; flappy_W(49, 276) <= 0; flappy_W(49, 277) <= 0; flappy_W(49, 278) <= 0; flappy_W(49, 279) <= 0; flappy_W(49, 280) <= 0; flappy_W(49, 281) <= 0; flappy_W(49, 282) <= 0; flappy_W(49, 283) <= 0; flappy_W(49, 284) <= 0; flappy_W(49, 285) <= 0; flappy_W(49, 286) <= 0; flappy_W(49, 287) <= 0; flappy_W(49, 288) <= 1; flappy_W(49, 289) <= 1; flappy_W(49, 290) <= 1; flappy_W(49, 291) <= 1; flappy_W(49, 292) <= 1; flappy_W(49, 293) <= 1; flappy_W(49, 294) <= 1; flappy_W(49, 295) <= 1; flappy_W(49, 296) <= 1; flappy_W(49, 297) <= 1; flappy_W(49, 298) <= 1; flappy_W(49, 299) <= 1; flappy_W(49, 300) <= 0; flappy_W(49, 301) <= 0; flappy_W(49, 302) <= 0; flappy_W(49, 303) <= 0; flappy_W(49, 304) <= 0; flappy_W(49, 305) <= 0; flappy_W(49, 306) <= 0; flappy_W(49, 307) <= 0; flappy_W(49, 308) <= 0; flappy_W(49, 309) <= 0; flappy_W(49, 310) <= 0; flappy_W(49, 311) <= 0; flappy_W(49, 312) <= 0; flappy_W(49, 313) <= 0; flappy_W(49, 314) <= 0; flappy_W(49, 315) <= 0; flappy_W(49, 316) <= 0; flappy_W(49, 317) <= 0; flappy_W(49, 318) <= 0; flappy_W(49, 319) <= 0; flappy_W(49, 320) <= 0; flappy_W(49, 321) <= 0; flappy_W(49, 322) <= 0; flappy_W(49, 323) <= 0; flappy_W(49, 324) <= 0; flappy_W(49, 325) <= 0; flappy_W(49, 326) <= 0; flappy_W(49, 327) <= 0; flappy_W(49, 328) <= 0; flappy_W(49, 329) <= 0; flappy_W(49, 330) <= 0; flappy_W(49, 331) <= 0; flappy_W(49, 332) <= 0; flappy_W(49, 333) <= 0; flappy_W(49, 334) <= 0; flappy_W(49, 335) <= 0; flappy_W(49, 336) <= 0; flappy_W(49, 337) <= 0; flappy_W(49, 338) <= 0; flappy_W(49, 339) <= 0; flappy_W(49, 340) <= 0; flappy_W(49, 341) <= 0; flappy_W(49, 342) <= 0; flappy_W(49, 343) <= 0; flappy_W(49, 344) <= 0; flappy_W(49, 345) <= 0; flappy_W(49, 346) <= 0; flappy_W(49, 347) <= 0; flappy_W(49, 348) <= 0; flappy_W(49, 349) <= 0; flappy_W(49, 350) <= 0; flappy_W(49, 351) <= 0; flappy_W(49, 352) <= 0; flappy_W(49, 353) <= 0; flappy_W(49, 354) <= 0; flappy_W(49, 355) <= 0; flappy_W(49, 356) <= 0; flappy_W(49, 357) <= 0; flappy_W(49, 358) <= 0; flappy_W(49, 359) <= 0; flappy_W(49, 360) <= 0; flappy_W(49, 361) <= 0; flappy_W(49, 362) <= 0; flappy_W(49, 363) <= 0; flappy_W(49, 364) <= 0; flappy_W(49, 365) <= 0; flappy_W(49, 366) <= 0; flappy_W(49, 367) <= 0; flappy_W(49, 368) <= 0; flappy_W(49, 369) <= 0; flappy_W(49, 370) <= 0; flappy_W(49, 371) <= 0; flappy_W(49, 372) <= 0; flappy_W(49, 373) <= 0; flappy_W(49, 374) <= 0; flappy_W(49, 375) <= 0; flappy_W(49, 376) <= 0; flappy_W(49, 377) <= 0; flappy_W(49, 378) <= 0; flappy_W(49, 379) <= 0; flappy_W(49, 380) <= 0; flappy_W(49, 381) <= 0; flappy_W(49, 382) <= 0; flappy_W(49, 383) <= 0; flappy_W(49, 384) <= 0; flappy_W(49, 385) <= 0; flappy_W(49, 386) <= 0; flappy_W(49, 387) <= 0; flappy_W(49, 388) <= 0; flappy_W(49, 389) <= 0; flappy_W(49, 390) <= 0; flappy_W(49, 391) <= 0; flappy_W(49, 392) <= 0; flappy_W(49, 393) <= 0; flappy_W(49, 394) <= 0; flappy_W(49, 395) <= 0; flappy_W(49, 396) <= 0; flappy_W(49, 397) <= 0; flappy_W(49, 398) <= 0; flappy_W(49, 399) <= 0; flappy_W(49, 400) <= 0; flappy_W(49, 401) <= 0; flappy_W(49, 402) <= 1; flappy_W(49, 403) <= 1; flappy_W(49, 404) <= 1; flappy_W(49, 405) <= 1; flappy_W(49, 406) <= 1; flappy_W(49, 407) <= 1; flappy_W(49, 408) <= 1; flappy_W(49, 409) <= 1; flappy_W(49, 410) <= 1; flappy_W(49, 411) <= 1; flappy_W(49, 412) <= 1; flappy_W(49, 413) <= 1; flappy_W(49, 414) <= 0; flappy_W(49, 415) <= 0; flappy_W(49, 416) <= 0; flappy_W(49, 417) <= 0; flappy_W(49, 418) <= 0; flappy_W(49, 419) <= 0; flappy_W(49, 420) <= 0; flappy_W(49, 421) <= 0; flappy_W(49, 422) <= 0; flappy_W(49, 423) <= 0; flappy_W(49, 424) <= 0; flappy_W(49, 425) <= 0; flappy_W(49, 426) <= 1; flappy_W(49, 427) <= 1; flappy_W(49, 428) <= 1; flappy_W(49, 429) <= 1; flappy_W(49, 430) <= 1; flappy_W(49, 431) <= 1; flappy_W(49, 432) <= 1; flappy_W(49, 433) <= 1; flappy_W(49, 434) <= 1; flappy_W(49, 435) <= 1; flappy_W(49, 436) <= 1; flappy_W(49, 437) <= 1; flappy_W(49, 438) <= 0; flappy_W(49, 439) <= 0; flappy_W(49, 440) <= 0; flappy_W(49, 441) <= 0; flappy_W(49, 442) <= 0; flappy_W(49, 443) <= 0; flappy_W(49, 444) <= 0; flappy_W(49, 445) <= 0; flappy_W(49, 446) <= 0; flappy_W(49, 447) <= 0; flappy_W(49, 448) <= 0; flappy_W(49, 449) <= 0; flappy_W(49, 450) <= 0; flappy_W(49, 451) <= 0; flappy_W(49, 452) <= 0; flappy_W(49, 453) <= 0; flappy_W(49, 454) <= 0; flappy_W(49, 455) <= 0; flappy_W(49, 456) <= 0; flappy_W(49, 457) <= 0; flappy_W(49, 458) <= 0; flappy_W(49, 459) <= 0; flappy_W(49, 460) <= 0; flappy_W(49, 461) <= 0; flappy_W(49, 462) <= 0; flappy_W(49, 463) <= 0; flappy_W(49, 464) <= 0; flappy_W(49, 465) <= 0; flappy_W(49, 466) <= 0; flappy_W(49, 467) <= 0; flappy_W(49, 468) <= 1; flappy_W(49, 469) <= 1; flappy_W(49, 470) <= 1; flappy_W(49, 471) <= 1; flappy_W(49, 472) <= 1; flappy_W(49, 473) <= 1; flappy_W(49, 474) <= 1; flappy_W(49, 475) <= 1; flappy_W(49, 476) <= 1; flappy_W(49, 477) <= 1; flappy_W(49, 478) <= 1; flappy_W(49, 479) <= 1; flappy_W(49, 480) <= 0; flappy_W(49, 481) <= 0; flappy_W(49, 482) <= 0; flappy_W(49, 483) <= 0; flappy_W(49, 484) <= 0; flappy_W(49, 485) <= 0; flappy_W(49, 486) <= 0; flappy_W(49, 487) <= 0; flappy_W(49, 488) <= 0; flappy_W(49, 489) <= 0; flappy_W(49, 490) <= 0; flappy_W(49, 491) <= 0; flappy_W(49, 492) <= 0; flappy_W(49, 493) <= 0; flappy_W(49, 494) <= 0; flappy_W(49, 495) <= 0; flappy_W(49, 496) <= 0; flappy_W(49, 497) <= 0; flappy_W(49, 498) <= 0; flappy_W(49, 499) <= 0; flappy_W(49, 500) <= 0; flappy_W(49, 501) <= 0; flappy_W(49, 502) <= 0; flappy_W(49, 503) <= 0; flappy_W(49, 504) <= 0; flappy_W(49, 505) <= 0; flappy_W(49, 506) <= 0; flappy_W(49, 507) <= 0; flappy_W(49, 508) <= 0; flappy_W(49, 509) <= 0; flappy_W(49, 510) <= 1; flappy_W(49, 511) <= 1; flappy_W(49, 512) <= 1; flappy_W(49, 513) <= 1; flappy_W(49, 514) <= 1; flappy_W(49, 515) <= 1; flappy_W(49, 516) <= 1; flappy_W(49, 517) <= 1; flappy_W(49, 518) <= 1; flappy_W(49, 519) <= 1; flappy_W(49, 520) <= 1; flappy_W(49, 521) <= 1; flappy_W(49, 522) <= 0; flappy_W(49, 523) <= 0; flappy_W(49, 524) <= 0; flappy_W(49, 525) <= 0; flappy_W(49, 526) <= 0; flappy_W(49, 527) <= 0; flappy_W(49, 528) <= 0; flappy_W(49, 529) <= 0; flappy_W(49, 530) <= 0; flappy_W(49, 531) <= 0; flappy_W(49, 532) <= 0; flappy_W(49, 533) <= 0; flappy_W(49, 534) <= 1; flappy_W(49, 535) <= 1; flappy_W(49, 536) <= 1; flappy_W(49, 537) <= 1; flappy_W(49, 538) <= 1; flappy_W(49, 539) <= 1; flappy_W(49, 540) <= 1; flappy_W(49, 541) <= 1; flappy_W(49, 542) <= 1; flappy_W(49, 543) <= 1; flappy_W(49, 544) <= 1; flappy_W(49, 545) <= 1; flappy_W(49, 546) <= 0; flappy_W(49, 547) <= 0; flappy_W(49, 548) <= 0; flappy_W(49, 549) <= 0; flappy_W(49, 550) <= 0; flappy_W(49, 551) <= 0; flappy_W(49, 552) <= 0; flappy_W(49, 553) <= 0; flappy_W(49, 554) <= 0; flappy_W(49, 555) <= 0; flappy_W(49, 556) <= 0; flappy_W(49, 557) <= 0; flappy_W(49, 558) <= 0; flappy_W(49, 559) <= 0; flappy_W(49, 560) <= 0; flappy_W(49, 561) <= 0; flappy_W(49, 562) <= 0; flappy_W(49, 563) <= 0; flappy_W(49, 564) <= 1; flappy_W(49, 565) <= 1; flappy_W(49, 566) <= 1; flappy_W(49, 567) <= 1; flappy_W(49, 568) <= 1; flappy_W(49, 569) <= 1; flappy_W(49, 570) <= 1; flappy_W(49, 571) <= 1; flappy_W(49, 572) <= 1; flappy_W(49, 573) <= 1; flappy_W(49, 574) <= 1; flappy_W(49, 575) <= 1; flappy_W(49, 576) <= 0; flappy_W(49, 577) <= 0; flappy_W(49, 578) <= 0; flappy_W(49, 579) <= 0; flappy_W(49, 580) <= 0; flappy_W(49, 581) <= 0; flappy_W(49, 582) <= 1; flappy_W(49, 583) <= 1; flappy_W(49, 584) <= 1; flappy_W(49, 585) <= 1; flappy_W(49, 586) <= 1; flappy_W(49, 587) <= 1; flappy_W(49, 588) <= 1; flappy_W(49, 589) <= 1; flappy_W(49, 590) <= 1; flappy_W(49, 591) <= 1; flappy_W(49, 592) <= 1; flappy_W(49, 593) <= 1; 
flappy_W(50, 0) <= 0; flappy_W(50, 1) <= 0; flappy_W(50, 2) <= 0; flappy_W(50, 3) <= 0; flappy_W(50, 4) <= 0; flappy_W(50, 5) <= 0; flappy_W(50, 6) <= 1; flappy_W(50, 7) <= 1; flappy_W(50, 8) <= 1; flappy_W(50, 9) <= 1; flappy_W(50, 10) <= 1; flappy_W(50, 11) <= 1; flappy_W(50, 12) <= 1; flappy_W(50, 13) <= 1; flappy_W(50, 14) <= 1; flappy_W(50, 15) <= 1; flappy_W(50, 16) <= 1; flappy_W(50, 17) <= 1; flappy_W(50, 18) <= 0; flappy_W(50, 19) <= 0; flappy_W(50, 20) <= 0; flappy_W(50, 21) <= 0; flappy_W(50, 22) <= 0; flappy_W(50, 23) <= 0; flappy_W(50, 24) <= 0; flappy_W(50, 25) <= 0; flappy_W(50, 26) <= 0; flappy_W(50, 27) <= 0; flappy_W(50, 28) <= 0; flappy_W(50, 29) <= 0; flappy_W(50, 30) <= 0; flappy_W(50, 31) <= 0; flappy_W(50, 32) <= 0; flappy_W(50, 33) <= 0; flappy_W(50, 34) <= 0; flappy_W(50, 35) <= 0; flappy_W(50, 36) <= 0; flappy_W(50, 37) <= 0; flappy_W(50, 38) <= 0; flappy_W(50, 39) <= 0; flappy_W(50, 40) <= 0; flappy_W(50, 41) <= 0; flappy_W(50, 42) <= 0; flappy_W(50, 43) <= 0; flappy_W(50, 44) <= 0; flappy_W(50, 45) <= 0; flappy_W(50, 46) <= 0; flappy_W(50, 47) <= 0; flappy_W(50, 48) <= 0; flappy_W(50, 49) <= 0; flappy_W(50, 50) <= 0; flappy_W(50, 51) <= 0; flappy_W(50, 52) <= 0; flappy_W(50, 53) <= 0; flappy_W(50, 54) <= 0; flappy_W(50, 55) <= 0; flappy_W(50, 56) <= 0; flappy_W(50, 57) <= 0; flappy_W(50, 58) <= 0; flappy_W(50, 59) <= 0; flappy_W(50, 60) <= 1; flappy_W(50, 61) <= 1; flappy_W(50, 62) <= 1; flappy_W(50, 63) <= 1; flappy_W(50, 64) <= 1; flappy_W(50, 65) <= 1; flappy_W(50, 66) <= 1; flappy_W(50, 67) <= 1; flappy_W(50, 68) <= 1; flappy_W(50, 69) <= 1; flappy_W(50, 70) <= 1; flappy_W(50, 71) <= 1; flappy_W(50, 72) <= 0; flappy_W(50, 73) <= 0; flappy_W(50, 74) <= 0; flappy_W(50, 75) <= 0; flappy_W(50, 76) <= 0; flappy_W(50, 77) <= 0; flappy_W(50, 78) <= 0; flappy_W(50, 79) <= 0; flappy_W(50, 80) <= 0; flappy_W(50, 81) <= 0; flappy_W(50, 82) <= 0; flappy_W(50, 83) <= 0; flappy_W(50, 84) <= 1; flappy_W(50, 85) <= 1; flappy_W(50, 86) <= 1; flappy_W(50, 87) <= 1; flappy_W(50, 88) <= 1; flappy_W(50, 89) <= 1; flappy_W(50, 90) <= 1; flappy_W(50, 91) <= 1; flappy_W(50, 92) <= 1; flappy_W(50, 93) <= 1; flappy_W(50, 94) <= 1; flappy_W(50, 95) <= 1; flappy_W(50, 96) <= 0; flappy_W(50, 97) <= 0; flappy_W(50, 98) <= 0; flappy_W(50, 99) <= 0; flappy_W(50, 100) <= 0; flappy_W(50, 101) <= 0; flappy_W(50, 102) <= 0; flappy_W(50, 103) <= 0; flappy_W(50, 104) <= 0; flappy_W(50, 105) <= 0; flappy_W(50, 106) <= 0; flappy_W(50, 107) <= 0; flappy_W(50, 108) <= 1; flappy_W(50, 109) <= 1; flappy_W(50, 110) <= 1; flappy_W(50, 111) <= 1; flappy_W(50, 112) <= 1; flappy_W(50, 113) <= 1; flappy_W(50, 114) <= 1; flappy_W(50, 115) <= 1; flappy_W(50, 116) <= 1; flappy_W(50, 117) <= 1; flappy_W(50, 118) <= 1; flappy_W(50, 119) <= 1; flappy_W(50, 120) <= 0; flappy_W(50, 121) <= 0; flappy_W(50, 122) <= 0; flappy_W(50, 123) <= 0; flappy_W(50, 124) <= 0; flappy_W(50, 125) <= 0; flappy_W(50, 126) <= 0; flappy_W(50, 127) <= 0; flappy_W(50, 128) <= 0; flappy_W(50, 129) <= 0; flappy_W(50, 130) <= 0; flappy_W(50, 131) <= 0; flappy_W(50, 132) <= 0; flappy_W(50, 133) <= 0; flappy_W(50, 134) <= 0; flappy_W(50, 135) <= 0; flappy_W(50, 136) <= 0; flappy_W(50, 137) <= 0; flappy_W(50, 138) <= 1; flappy_W(50, 139) <= 1; flappy_W(50, 140) <= 1; flappy_W(50, 141) <= 1; flappy_W(50, 142) <= 1; flappy_W(50, 143) <= 1; flappy_W(50, 144) <= 1; flappy_W(50, 145) <= 1; flappy_W(50, 146) <= 1; flappy_W(50, 147) <= 1; flappy_W(50, 148) <= 1; flappy_W(50, 149) <= 1; flappy_W(50, 150) <= 0; flappy_W(50, 151) <= 0; flappy_W(50, 152) <= 0; flappy_W(50, 153) <= 0; flappy_W(50, 154) <= 0; flappy_W(50, 155) <= 0; flappy_W(50, 156) <= 0; flappy_W(50, 157) <= 0; flappy_W(50, 158) <= 0; flappy_W(50, 159) <= 0; flappy_W(50, 160) <= 0; flappy_W(50, 161) <= 0; flappy_W(50, 162) <= 0; flappy_W(50, 163) <= 0; flappy_W(50, 164) <= 0; flappy_W(50, 165) <= 0; flappy_W(50, 166) <= 0; flappy_W(50, 167) <= 0; flappy_W(50, 168) <= 1; flappy_W(50, 169) <= 1; flappy_W(50, 170) <= 1; flappy_W(50, 171) <= 1; flappy_W(50, 172) <= 1; flappy_W(50, 173) <= 1; flappy_W(50, 174) <= 1; flappy_W(50, 175) <= 1; flappy_W(50, 176) <= 1; flappy_W(50, 177) <= 1; flappy_W(50, 178) <= 1; flappy_W(50, 179) <= 1; flappy_W(50, 180) <= 0; flappy_W(50, 181) <= 0; flappy_W(50, 182) <= 0; flappy_W(50, 183) <= 0; flappy_W(50, 184) <= 0; flappy_W(50, 185) <= 0; flappy_W(50, 186) <= 0; flappy_W(50, 187) <= 0; flappy_W(50, 188) <= 0; flappy_W(50, 189) <= 0; flappy_W(50, 190) <= 0; flappy_W(50, 191) <= 0; flappy_W(50, 192) <= 0; flappy_W(50, 193) <= 0; flappy_W(50, 194) <= 0; flappy_W(50, 195) <= 0; flappy_W(50, 196) <= 0; flappy_W(50, 197) <= 0; flappy_W(50, 198) <= 0; flappy_W(50, 199) <= 0; flappy_W(50, 200) <= 0; flappy_W(50, 201) <= 0; flappy_W(50, 202) <= 0; flappy_W(50, 203) <= 0; flappy_W(50, 204) <= 0; flappy_W(50, 205) <= 0; flappy_W(50, 206) <= 0; flappy_W(50, 207) <= 0; flappy_W(50, 208) <= 0; flappy_W(50, 209) <= 0; flappy_W(50, 210) <= 0; flappy_W(50, 211) <= 0; flappy_W(50, 212) <= 0; flappy_W(50, 213) <= 0; flappy_W(50, 214) <= 0; flappy_W(50, 215) <= 0; flappy_W(50, 216) <= 0; flappy_W(50, 217) <= 0; flappy_W(50, 218) <= 0; flappy_W(50, 219) <= 0; flappy_W(50, 220) <= 0; flappy_W(50, 221) <= 0; flappy_W(50, 222) <= 1; flappy_W(50, 223) <= 1; flappy_W(50, 224) <= 1; flappy_W(50, 225) <= 1; flappy_W(50, 226) <= 1; flappy_W(50, 227) <= 1; flappy_W(50, 228) <= 1; flappy_W(50, 229) <= 1; flappy_W(50, 230) <= 1; flappy_W(50, 231) <= 1; flappy_W(50, 232) <= 1; flappy_W(50, 233) <= 1; flappy_W(50, 234) <= 0; flappy_W(50, 235) <= 0; flappy_W(50, 236) <= 0; flappy_W(50, 237) <= 0; flappy_W(50, 238) <= 0; flappy_W(50, 239) <= 0; flappy_W(50, 240) <= 0; flappy_W(50, 241) <= 0; flappy_W(50, 242) <= 0; flappy_W(50, 243) <= 0; flappy_W(50, 244) <= 0; flappy_W(50, 245) <= 0; flappy_W(50, 246) <= 0; flappy_W(50, 247) <= 0; flappy_W(50, 248) <= 0; flappy_W(50, 249) <= 0; flappy_W(50, 250) <= 0; flappy_W(50, 251) <= 0; flappy_W(50, 252) <= 0; flappy_W(50, 253) <= 0; flappy_W(50, 254) <= 0; flappy_W(50, 255) <= 0; flappy_W(50, 256) <= 0; flappy_W(50, 257) <= 0; flappy_W(50, 258) <= 0; flappy_W(50, 259) <= 0; flappy_W(50, 260) <= 0; flappy_W(50, 261) <= 0; flappy_W(50, 262) <= 0; flappy_W(50, 263) <= 0; flappy_W(50, 264) <= 0; flappy_W(50, 265) <= 0; flappy_W(50, 266) <= 0; flappy_W(50, 267) <= 0; flappy_W(50, 268) <= 0; flappy_W(50, 269) <= 0; flappy_W(50, 270) <= 0; flappy_W(50, 271) <= 0; flappy_W(50, 272) <= 0; flappy_W(50, 273) <= 0; flappy_W(50, 274) <= 0; flappy_W(50, 275) <= 0; flappy_W(50, 276) <= 0; flappy_W(50, 277) <= 0; flappy_W(50, 278) <= 0; flappy_W(50, 279) <= 0; flappy_W(50, 280) <= 0; flappy_W(50, 281) <= 0; flappy_W(50, 282) <= 0; flappy_W(50, 283) <= 0; flappy_W(50, 284) <= 0; flappy_W(50, 285) <= 0; flappy_W(50, 286) <= 0; flappy_W(50, 287) <= 0; flappy_W(50, 288) <= 1; flappy_W(50, 289) <= 1; flappy_W(50, 290) <= 1; flappy_W(50, 291) <= 1; flappy_W(50, 292) <= 1; flappy_W(50, 293) <= 1; flappy_W(50, 294) <= 1; flappy_W(50, 295) <= 1; flappy_W(50, 296) <= 1; flappy_W(50, 297) <= 1; flappy_W(50, 298) <= 1; flappy_W(50, 299) <= 1; flappy_W(50, 300) <= 0; flappy_W(50, 301) <= 0; flappy_W(50, 302) <= 0; flappy_W(50, 303) <= 0; flappy_W(50, 304) <= 0; flappy_W(50, 305) <= 0; flappy_W(50, 306) <= 0; flappy_W(50, 307) <= 0; flappy_W(50, 308) <= 0; flappy_W(50, 309) <= 0; flappy_W(50, 310) <= 0; flappy_W(50, 311) <= 0; flappy_W(50, 312) <= 0; flappy_W(50, 313) <= 0; flappy_W(50, 314) <= 0; flappy_W(50, 315) <= 0; flappy_W(50, 316) <= 0; flappy_W(50, 317) <= 0; flappy_W(50, 318) <= 0; flappy_W(50, 319) <= 0; flappy_W(50, 320) <= 0; flappy_W(50, 321) <= 0; flappy_W(50, 322) <= 0; flappy_W(50, 323) <= 0; flappy_W(50, 324) <= 0; flappy_W(50, 325) <= 0; flappy_W(50, 326) <= 0; flappy_W(50, 327) <= 0; flappy_W(50, 328) <= 0; flappy_W(50, 329) <= 0; flappy_W(50, 330) <= 0; flappy_W(50, 331) <= 0; flappy_W(50, 332) <= 0; flappy_W(50, 333) <= 0; flappy_W(50, 334) <= 0; flappy_W(50, 335) <= 0; flappy_W(50, 336) <= 0; flappy_W(50, 337) <= 0; flappy_W(50, 338) <= 0; flappy_W(50, 339) <= 0; flappy_W(50, 340) <= 0; flappy_W(50, 341) <= 0; flappy_W(50, 342) <= 0; flappy_W(50, 343) <= 0; flappy_W(50, 344) <= 0; flappy_W(50, 345) <= 0; flappy_W(50, 346) <= 0; flappy_W(50, 347) <= 0; flappy_W(50, 348) <= 0; flappy_W(50, 349) <= 0; flappy_W(50, 350) <= 0; flappy_W(50, 351) <= 0; flappy_W(50, 352) <= 0; flappy_W(50, 353) <= 0; flappy_W(50, 354) <= 0; flappy_W(50, 355) <= 0; flappy_W(50, 356) <= 0; flappy_W(50, 357) <= 0; flappy_W(50, 358) <= 0; flappy_W(50, 359) <= 0; flappy_W(50, 360) <= 0; flappy_W(50, 361) <= 0; flappy_W(50, 362) <= 0; flappy_W(50, 363) <= 0; flappy_W(50, 364) <= 0; flappy_W(50, 365) <= 0; flappy_W(50, 366) <= 0; flappy_W(50, 367) <= 0; flappy_W(50, 368) <= 0; flappy_W(50, 369) <= 0; flappy_W(50, 370) <= 0; flappy_W(50, 371) <= 0; flappy_W(50, 372) <= 0; flappy_W(50, 373) <= 0; flappy_W(50, 374) <= 0; flappy_W(50, 375) <= 0; flappy_W(50, 376) <= 0; flappy_W(50, 377) <= 0; flappy_W(50, 378) <= 0; flappy_W(50, 379) <= 0; flappy_W(50, 380) <= 0; flappy_W(50, 381) <= 0; flappy_W(50, 382) <= 0; flappy_W(50, 383) <= 0; flappy_W(50, 384) <= 0; flappy_W(50, 385) <= 0; flappy_W(50, 386) <= 0; flappy_W(50, 387) <= 0; flappy_W(50, 388) <= 0; flappy_W(50, 389) <= 0; flappy_W(50, 390) <= 0; flappy_W(50, 391) <= 0; flappy_W(50, 392) <= 0; flappy_W(50, 393) <= 0; flappy_W(50, 394) <= 0; flappy_W(50, 395) <= 0; flappy_W(50, 396) <= 0; flappy_W(50, 397) <= 0; flappy_W(50, 398) <= 0; flappy_W(50, 399) <= 0; flappy_W(50, 400) <= 0; flappy_W(50, 401) <= 0; flappy_W(50, 402) <= 1; flappy_W(50, 403) <= 1; flappy_W(50, 404) <= 1; flappy_W(50, 405) <= 1; flappy_W(50, 406) <= 1; flappy_W(50, 407) <= 1; flappy_W(50, 408) <= 1; flappy_W(50, 409) <= 1; flappy_W(50, 410) <= 1; flappy_W(50, 411) <= 1; flappy_W(50, 412) <= 1; flappy_W(50, 413) <= 1; flappy_W(50, 414) <= 0; flappy_W(50, 415) <= 0; flappy_W(50, 416) <= 0; flappy_W(50, 417) <= 0; flappy_W(50, 418) <= 0; flappy_W(50, 419) <= 0; flappy_W(50, 420) <= 0; flappy_W(50, 421) <= 0; flappy_W(50, 422) <= 0; flappy_W(50, 423) <= 0; flappy_W(50, 424) <= 0; flappy_W(50, 425) <= 0; flappy_W(50, 426) <= 1; flappy_W(50, 427) <= 1; flappy_W(50, 428) <= 1; flappy_W(50, 429) <= 1; flappy_W(50, 430) <= 1; flappy_W(50, 431) <= 1; flappy_W(50, 432) <= 1; flappy_W(50, 433) <= 1; flappy_W(50, 434) <= 1; flappy_W(50, 435) <= 1; flappy_W(50, 436) <= 1; flappy_W(50, 437) <= 1; flappy_W(50, 438) <= 0; flappy_W(50, 439) <= 0; flappy_W(50, 440) <= 0; flappy_W(50, 441) <= 0; flappy_W(50, 442) <= 0; flappy_W(50, 443) <= 0; flappy_W(50, 444) <= 0; flappy_W(50, 445) <= 0; flappy_W(50, 446) <= 0; flappy_W(50, 447) <= 0; flappy_W(50, 448) <= 0; flappy_W(50, 449) <= 0; flappy_W(50, 450) <= 0; flappy_W(50, 451) <= 0; flappy_W(50, 452) <= 0; flappy_W(50, 453) <= 0; flappy_W(50, 454) <= 0; flappy_W(50, 455) <= 0; flappy_W(50, 456) <= 0; flappy_W(50, 457) <= 0; flappy_W(50, 458) <= 0; flappy_W(50, 459) <= 0; flappy_W(50, 460) <= 0; flappy_W(50, 461) <= 0; flappy_W(50, 462) <= 0; flappy_W(50, 463) <= 0; flappy_W(50, 464) <= 0; flappy_W(50, 465) <= 0; flappy_W(50, 466) <= 0; flappy_W(50, 467) <= 0; flappy_W(50, 468) <= 1; flappy_W(50, 469) <= 1; flappy_W(50, 470) <= 1; flappy_W(50, 471) <= 1; flappy_W(50, 472) <= 1; flappy_W(50, 473) <= 1; flappy_W(50, 474) <= 1; flappy_W(50, 475) <= 1; flappy_W(50, 476) <= 1; flappy_W(50, 477) <= 1; flappy_W(50, 478) <= 1; flappy_W(50, 479) <= 1; flappy_W(50, 480) <= 0; flappy_W(50, 481) <= 0; flappy_W(50, 482) <= 0; flappy_W(50, 483) <= 0; flappy_W(50, 484) <= 0; flappy_W(50, 485) <= 0; flappy_W(50, 486) <= 0; flappy_W(50, 487) <= 0; flappy_W(50, 488) <= 0; flappy_W(50, 489) <= 0; flappy_W(50, 490) <= 0; flappy_W(50, 491) <= 0; flappy_W(50, 492) <= 0; flappy_W(50, 493) <= 0; flappy_W(50, 494) <= 0; flappy_W(50, 495) <= 0; flappy_W(50, 496) <= 0; flappy_W(50, 497) <= 0; flappy_W(50, 498) <= 0; flappy_W(50, 499) <= 0; flappy_W(50, 500) <= 0; flappy_W(50, 501) <= 0; flappy_W(50, 502) <= 0; flappy_W(50, 503) <= 0; flappy_W(50, 504) <= 0; flappy_W(50, 505) <= 0; flappy_W(50, 506) <= 0; flappy_W(50, 507) <= 0; flappy_W(50, 508) <= 0; flappy_W(50, 509) <= 0; flappy_W(50, 510) <= 1; flappy_W(50, 511) <= 1; flappy_W(50, 512) <= 1; flappy_W(50, 513) <= 1; flappy_W(50, 514) <= 1; flappy_W(50, 515) <= 1; flappy_W(50, 516) <= 1; flappy_W(50, 517) <= 1; flappy_W(50, 518) <= 1; flappy_W(50, 519) <= 1; flappy_W(50, 520) <= 1; flappy_W(50, 521) <= 1; flappy_W(50, 522) <= 0; flappy_W(50, 523) <= 0; flappy_W(50, 524) <= 0; flappy_W(50, 525) <= 0; flappy_W(50, 526) <= 0; flappy_W(50, 527) <= 0; flappy_W(50, 528) <= 0; flappy_W(50, 529) <= 0; flappy_W(50, 530) <= 0; flappy_W(50, 531) <= 0; flappy_W(50, 532) <= 0; flappy_W(50, 533) <= 0; flappy_W(50, 534) <= 1; flappy_W(50, 535) <= 1; flappy_W(50, 536) <= 1; flappy_W(50, 537) <= 1; flappy_W(50, 538) <= 1; flappy_W(50, 539) <= 1; flappy_W(50, 540) <= 1; flappy_W(50, 541) <= 1; flappy_W(50, 542) <= 1; flappy_W(50, 543) <= 1; flappy_W(50, 544) <= 1; flappy_W(50, 545) <= 1; flappy_W(50, 546) <= 0; flappy_W(50, 547) <= 0; flappy_W(50, 548) <= 0; flappy_W(50, 549) <= 0; flappy_W(50, 550) <= 0; flappy_W(50, 551) <= 0; flappy_W(50, 552) <= 0; flappy_W(50, 553) <= 0; flappy_W(50, 554) <= 0; flappy_W(50, 555) <= 0; flappy_W(50, 556) <= 0; flappy_W(50, 557) <= 0; flappy_W(50, 558) <= 0; flappy_W(50, 559) <= 0; flappy_W(50, 560) <= 0; flappy_W(50, 561) <= 0; flappy_W(50, 562) <= 0; flappy_W(50, 563) <= 0; flappy_W(50, 564) <= 1; flappy_W(50, 565) <= 1; flappy_W(50, 566) <= 1; flappy_W(50, 567) <= 1; flappy_W(50, 568) <= 1; flappy_W(50, 569) <= 1; flappy_W(50, 570) <= 1; flappy_W(50, 571) <= 1; flappy_W(50, 572) <= 1; flappy_W(50, 573) <= 1; flappy_W(50, 574) <= 1; flappy_W(50, 575) <= 1; flappy_W(50, 576) <= 0; flappy_W(50, 577) <= 0; flappy_W(50, 578) <= 0; flappy_W(50, 579) <= 0; flappy_W(50, 580) <= 0; flappy_W(50, 581) <= 0; flappy_W(50, 582) <= 1; flappy_W(50, 583) <= 1; flappy_W(50, 584) <= 1; flappy_W(50, 585) <= 1; flappy_W(50, 586) <= 1; flappy_W(50, 587) <= 1; flappy_W(50, 588) <= 1; flappy_W(50, 589) <= 1; flappy_W(50, 590) <= 1; flappy_W(50, 591) <= 1; flappy_W(50, 592) <= 1; flappy_W(50, 593) <= 1; 
flappy_W(51, 0) <= 0; flappy_W(51, 1) <= 0; flappy_W(51, 2) <= 0; flappy_W(51, 3) <= 0; flappy_W(51, 4) <= 0; flappy_W(51, 5) <= 0; flappy_W(51, 6) <= 1; flappy_W(51, 7) <= 1; flappy_W(51, 8) <= 1; flappy_W(51, 9) <= 1; flappy_W(51, 10) <= 1; flappy_W(51, 11) <= 1; flappy_W(51, 12) <= 1; flappy_W(51, 13) <= 1; flappy_W(51, 14) <= 1; flappy_W(51, 15) <= 1; flappy_W(51, 16) <= 1; flappy_W(51, 17) <= 1; flappy_W(51, 18) <= 0; flappy_W(51, 19) <= 0; flappy_W(51, 20) <= 0; flappy_W(51, 21) <= 0; flappy_W(51, 22) <= 0; flappy_W(51, 23) <= 0; flappy_W(51, 24) <= 0; flappy_W(51, 25) <= 0; flappy_W(51, 26) <= 0; flappy_W(51, 27) <= 0; flappy_W(51, 28) <= 0; flappy_W(51, 29) <= 0; flappy_W(51, 30) <= 0; flappy_W(51, 31) <= 0; flappy_W(51, 32) <= 0; flappy_W(51, 33) <= 0; flappy_W(51, 34) <= 0; flappy_W(51, 35) <= 0; flappy_W(51, 36) <= 0; flappy_W(51, 37) <= 0; flappy_W(51, 38) <= 0; flappy_W(51, 39) <= 0; flappy_W(51, 40) <= 0; flappy_W(51, 41) <= 0; flappy_W(51, 42) <= 0; flappy_W(51, 43) <= 0; flappy_W(51, 44) <= 0; flappy_W(51, 45) <= 0; flappy_W(51, 46) <= 0; flappy_W(51, 47) <= 0; flappy_W(51, 48) <= 0; flappy_W(51, 49) <= 0; flappy_W(51, 50) <= 0; flappy_W(51, 51) <= 0; flappy_W(51, 52) <= 0; flappy_W(51, 53) <= 0; flappy_W(51, 54) <= 0; flappy_W(51, 55) <= 0; flappy_W(51, 56) <= 0; flappy_W(51, 57) <= 0; flappy_W(51, 58) <= 0; flappy_W(51, 59) <= 0; flappy_W(51, 60) <= 1; flappy_W(51, 61) <= 1; flappy_W(51, 62) <= 1; flappy_W(51, 63) <= 1; flappy_W(51, 64) <= 1; flappy_W(51, 65) <= 1; flappy_W(51, 66) <= 1; flappy_W(51, 67) <= 1; flappy_W(51, 68) <= 1; flappy_W(51, 69) <= 1; flappy_W(51, 70) <= 1; flappy_W(51, 71) <= 1; flappy_W(51, 72) <= 0; flappy_W(51, 73) <= 0; flappy_W(51, 74) <= 0; flappy_W(51, 75) <= 0; flappy_W(51, 76) <= 0; flappy_W(51, 77) <= 0; flappy_W(51, 78) <= 0; flappy_W(51, 79) <= 0; flappy_W(51, 80) <= 0; flappy_W(51, 81) <= 0; flappy_W(51, 82) <= 0; flappy_W(51, 83) <= 0; flappy_W(51, 84) <= 1; flappy_W(51, 85) <= 1; flappy_W(51, 86) <= 1; flappy_W(51, 87) <= 1; flappy_W(51, 88) <= 1; flappy_W(51, 89) <= 1; flappy_W(51, 90) <= 1; flappy_W(51, 91) <= 1; flappy_W(51, 92) <= 1; flappy_W(51, 93) <= 1; flappy_W(51, 94) <= 1; flappy_W(51, 95) <= 1; flappy_W(51, 96) <= 0; flappy_W(51, 97) <= 0; flappy_W(51, 98) <= 0; flappy_W(51, 99) <= 0; flappy_W(51, 100) <= 0; flappy_W(51, 101) <= 0; flappy_W(51, 102) <= 0; flappy_W(51, 103) <= 0; flappy_W(51, 104) <= 0; flappy_W(51, 105) <= 0; flappy_W(51, 106) <= 0; flappy_W(51, 107) <= 0; flappy_W(51, 108) <= 1; flappy_W(51, 109) <= 1; flappy_W(51, 110) <= 1; flappy_W(51, 111) <= 1; flappy_W(51, 112) <= 1; flappy_W(51, 113) <= 1; flappy_W(51, 114) <= 1; flappy_W(51, 115) <= 1; flappy_W(51, 116) <= 1; flappy_W(51, 117) <= 1; flappy_W(51, 118) <= 1; flappy_W(51, 119) <= 1; flappy_W(51, 120) <= 0; flappy_W(51, 121) <= 0; flappy_W(51, 122) <= 0; flappy_W(51, 123) <= 0; flappy_W(51, 124) <= 0; flappy_W(51, 125) <= 0; flappy_W(51, 126) <= 0; flappy_W(51, 127) <= 0; flappy_W(51, 128) <= 0; flappy_W(51, 129) <= 0; flappy_W(51, 130) <= 0; flappy_W(51, 131) <= 0; flappy_W(51, 132) <= 0; flappy_W(51, 133) <= 0; flappy_W(51, 134) <= 0; flappy_W(51, 135) <= 0; flappy_W(51, 136) <= 0; flappy_W(51, 137) <= 0; flappy_W(51, 138) <= 1; flappy_W(51, 139) <= 1; flappy_W(51, 140) <= 1; flappy_W(51, 141) <= 1; flappy_W(51, 142) <= 1; flappy_W(51, 143) <= 1; flappy_W(51, 144) <= 1; flappy_W(51, 145) <= 1; flappy_W(51, 146) <= 1; flappy_W(51, 147) <= 1; flappy_W(51, 148) <= 1; flappy_W(51, 149) <= 1; flappy_W(51, 150) <= 0; flappy_W(51, 151) <= 0; flappy_W(51, 152) <= 0; flappy_W(51, 153) <= 0; flappy_W(51, 154) <= 0; flappy_W(51, 155) <= 0; flappy_W(51, 156) <= 0; flappy_W(51, 157) <= 0; flappy_W(51, 158) <= 0; flappy_W(51, 159) <= 0; flappy_W(51, 160) <= 0; flappy_W(51, 161) <= 0; flappy_W(51, 162) <= 0; flappy_W(51, 163) <= 0; flappy_W(51, 164) <= 0; flappy_W(51, 165) <= 0; flappy_W(51, 166) <= 0; flappy_W(51, 167) <= 0; flappy_W(51, 168) <= 1; flappy_W(51, 169) <= 1; flappy_W(51, 170) <= 1; flappy_W(51, 171) <= 1; flappy_W(51, 172) <= 1; flappy_W(51, 173) <= 1; flappy_W(51, 174) <= 1; flappy_W(51, 175) <= 1; flappy_W(51, 176) <= 1; flappy_W(51, 177) <= 1; flappy_W(51, 178) <= 1; flappy_W(51, 179) <= 1; flappy_W(51, 180) <= 0; flappy_W(51, 181) <= 0; flappy_W(51, 182) <= 0; flappy_W(51, 183) <= 0; flappy_W(51, 184) <= 0; flappy_W(51, 185) <= 0; flappy_W(51, 186) <= 0; flappy_W(51, 187) <= 0; flappy_W(51, 188) <= 0; flappy_W(51, 189) <= 0; flappy_W(51, 190) <= 0; flappy_W(51, 191) <= 0; flappy_W(51, 192) <= 0; flappy_W(51, 193) <= 0; flappy_W(51, 194) <= 0; flappy_W(51, 195) <= 0; flappy_W(51, 196) <= 0; flappy_W(51, 197) <= 0; flappy_W(51, 198) <= 0; flappy_W(51, 199) <= 0; flappy_W(51, 200) <= 0; flappy_W(51, 201) <= 0; flappy_W(51, 202) <= 0; flappy_W(51, 203) <= 0; flappy_W(51, 204) <= 0; flappy_W(51, 205) <= 0; flappy_W(51, 206) <= 0; flappy_W(51, 207) <= 0; flappy_W(51, 208) <= 0; flappy_W(51, 209) <= 0; flappy_W(51, 210) <= 0; flappy_W(51, 211) <= 0; flappy_W(51, 212) <= 0; flappy_W(51, 213) <= 0; flappy_W(51, 214) <= 0; flappy_W(51, 215) <= 0; flappy_W(51, 216) <= 0; flappy_W(51, 217) <= 0; flappy_W(51, 218) <= 0; flappy_W(51, 219) <= 0; flappy_W(51, 220) <= 0; flappy_W(51, 221) <= 0; flappy_W(51, 222) <= 1; flappy_W(51, 223) <= 1; flappy_W(51, 224) <= 1; flappy_W(51, 225) <= 1; flappy_W(51, 226) <= 1; flappy_W(51, 227) <= 1; flappy_W(51, 228) <= 1; flappy_W(51, 229) <= 1; flappy_W(51, 230) <= 1; flappy_W(51, 231) <= 1; flappy_W(51, 232) <= 1; flappy_W(51, 233) <= 1; flappy_W(51, 234) <= 0; flappy_W(51, 235) <= 0; flappy_W(51, 236) <= 0; flappy_W(51, 237) <= 0; flappy_W(51, 238) <= 0; flappy_W(51, 239) <= 0; flappy_W(51, 240) <= 0; flappy_W(51, 241) <= 0; flappy_W(51, 242) <= 0; flappy_W(51, 243) <= 0; flappy_W(51, 244) <= 0; flappy_W(51, 245) <= 0; flappy_W(51, 246) <= 0; flappy_W(51, 247) <= 0; flappy_W(51, 248) <= 0; flappy_W(51, 249) <= 0; flappy_W(51, 250) <= 0; flappy_W(51, 251) <= 0; flappy_W(51, 252) <= 0; flappy_W(51, 253) <= 0; flappy_W(51, 254) <= 0; flappy_W(51, 255) <= 0; flappy_W(51, 256) <= 0; flappy_W(51, 257) <= 0; flappy_W(51, 258) <= 0; flappy_W(51, 259) <= 0; flappy_W(51, 260) <= 0; flappy_W(51, 261) <= 0; flappy_W(51, 262) <= 0; flappy_W(51, 263) <= 0; flappy_W(51, 264) <= 0; flappy_W(51, 265) <= 0; flappy_W(51, 266) <= 0; flappy_W(51, 267) <= 0; flappy_W(51, 268) <= 0; flappy_W(51, 269) <= 0; flappy_W(51, 270) <= 0; flappy_W(51, 271) <= 0; flappy_W(51, 272) <= 0; flappy_W(51, 273) <= 0; flappy_W(51, 274) <= 0; flappy_W(51, 275) <= 0; flappy_W(51, 276) <= 0; flappy_W(51, 277) <= 0; flappy_W(51, 278) <= 0; flappy_W(51, 279) <= 0; flappy_W(51, 280) <= 0; flappy_W(51, 281) <= 0; flappy_W(51, 282) <= 0; flappy_W(51, 283) <= 0; flappy_W(51, 284) <= 0; flappy_W(51, 285) <= 0; flappy_W(51, 286) <= 0; flappy_W(51, 287) <= 0; flappy_W(51, 288) <= 1; flappy_W(51, 289) <= 1; flappy_W(51, 290) <= 1; flappy_W(51, 291) <= 1; flappy_W(51, 292) <= 1; flappy_W(51, 293) <= 1; flappy_W(51, 294) <= 1; flappy_W(51, 295) <= 1; flappy_W(51, 296) <= 1; flappy_W(51, 297) <= 1; flappy_W(51, 298) <= 1; flappy_W(51, 299) <= 1; flappy_W(51, 300) <= 0; flappy_W(51, 301) <= 0; flappy_W(51, 302) <= 0; flappy_W(51, 303) <= 0; flappy_W(51, 304) <= 0; flappy_W(51, 305) <= 0; flappy_W(51, 306) <= 0; flappy_W(51, 307) <= 0; flappy_W(51, 308) <= 0; flappy_W(51, 309) <= 0; flappy_W(51, 310) <= 0; flappy_W(51, 311) <= 0; flappy_W(51, 312) <= 0; flappy_W(51, 313) <= 0; flappy_W(51, 314) <= 0; flappy_W(51, 315) <= 0; flappy_W(51, 316) <= 0; flappy_W(51, 317) <= 0; flappy_W(51, 318) <= 0; flappy_W(51, 319) <= 0; flappy_W(51, 320) <= 0; flappy_W(51, 321) <= 0; flappy_W(51, 322) <= 0; flappy_W(51, 323) <= 0; flappy_W(51, 324) <= 0; flappy_W(51, 325) <= 0; flappy_W(51, 326) <= 0; flappy_W(51, 327) <= 0; flappy_W(51, 328) <= 0; flappy_W(51, 329) <= 0; flappy_W(51, 330) <= 0; flappy_W(51, 331) <= 0; flappy_W(51, 332) <= 0; flappy_W(51, 333) <= 0; flappy_W(51, 334) <= 0; flappy_W(51, 335) <= 0; flappy_W(51, 336) <= 0; flappy_W(51, 337) <= 0; flappy_W(51, 338) <= 0; flappy_W(51, 339) <= 0; flappy_W(51, 340) <= 0; flappy_W(51, 341) <= 0; flappy_W(51, 342) <= 0; flappy_W(51, 343) <= 0; flappy_W(51, 344) <= 0; flappy_W(51, 345) <= 0; flappy_W(51, 346) <= 0; flappy_W(51, 347) <= 0; flappy_W(51, 348) <= 0; flappy_W(51, 349) <= 0; flappy_W(51, 350) <= 0; flappy_W(51, 351) <= 0; flappy_W(51, 352) <= 0; flappy_W(51, 353) <= 0; flappy_W(51, 354) <= 0; flappy_W(51, 355) <= 0; flappy_W(51, 356) <= 0; flappy_W(51, 357) <= 0; flappy_W(51, 358) <= 0; flappy_W(51, 359) <= 0; flappy_W(51, 360) <= 0; flappy_W(51, 361) <= 0; flappy_W(51, 362) <= 0; flappy_W(51, 363) <= 0; flappy_W(51, 364) <= 0; flappy_W(51, 365) <= 0; flappy_W(51, 366) <= 0; flappy_W(51, 367) <= 0; flappy_W(51, 368) <= 0; flappy_W(51, 369) <= 0; flappy_W(51, 370) <= 0; flappy_W(51, 371) <= 0; flappy_W(51, 372) <= 0; flappy_W(51, 373) <= 0; flappy_W(51, 374) <= 0; flappy_W(51, 375) <= 0; flappy_W(51, 376) <= 0; flappy_W(51, 377) <= 0; flappy_W(51, 378) <= 0; flappy_W(51, 379) <= 0; flappy_W(51, 380) <= 0; flappy_W(51, 381) <= 0; flappy_W(51, 382) <= 0; flappy_W(51, 383) <= 0; flappy_W(51, 384) <= 0; flappy_W(51, 385) <= 0; flappy_W(51, 386) <= 0; flappy_W(51, 387) <= 0; flappy_W(51, 388) <= 0; flappy_W(51, 389) <= 0; flappy_W(51, 390) <= 0; flappy_W(51, 391) <= 0; flappy_W(51, 392) <= 0; flappy_W(51, 393) <= 0; flappy_W(51, 394) <= 0; flappy_W(51, 395) <= 0; flappy_W(51, 396) <= 0; flappy_W(51, 397) <= 0; flappy_W(51, 398) <= 0; flappy_W(51, 399) <= 0; flappy_W(51, 400) <= 0; flappy_W(51, 401) <= 0; flappy_W(51, 402) <= 1; flappy_W(51, 403) <= 1; flappy_W(51, 404) <= 1; flappy_W(51, 405) <= 1; flappy_W(51, 406) <= 1; flappy_W(51, 407) <= 1; flappy_W(51, 408) <= 1; flappy_W(51, 409) <= 1; flappy_W(51, 410) <= 1; flappy_W(51, 411) <= 1; flappy_W(51, 412) <= 1; flappy_W(51, 413) <= 1; flappy_W(51, 414) <= 0; flappy_W(51, 415) <= 0; flappy_W(51, 416) <= 0; flappy_W(51, 417) <= 0; flappy_W(51, 418) <= 0; flappy_W(51, 419) <= 0; flappy_W(51, 420) <= 0; flappy_W(51, 421) <= 0; flappy_W(51, 422) <= 0; flappy_W(51, 423) <= 0; flappy_W(51, 424) <= 0; flappy_W(51, 425) <= 0; flappy_W(51, 426) <= 1; flappy_W(51, 427) <= 1; flappy_W(51, 428) <= 1; flappy_W(51, 429) <= 1; flappy_W(51, 430) <= 1; flappy_W(51, 431) <= 1; flappy_W(51, 432) <= 1; flappy_W(51, 433) <= 1; flappy_W(51, 434) <= 1; flappy_W(51, 435) <= 1; flappy_W(51, 436) <= 1; flappy_W(51, 437) <= 1; flappy_W(51, 438) <= 0; flappy_W(51, 439) <= 0; flappy_W(51, 440) <= 0; flappy_W(51, 441) <= 0; flappy_W(51, 442) <= 0; flappy_W(51, 443) <= 0; flappy_W(51, 444) <= 0; flappy_W(51, 445) <= 0; flappy_W(51, 446) <= 0; flappy_W(51, 447) <= 0; flappy_W(51, 448) <= 0; flappy_W(51, 449) <= 0; flappy_W(51, 450) <= 0; flappy_W(51, 451) <= 0; flappy_W(51, 452) <= 0; flappy_W(51, 453) <= 0; flappy_W(51, 454) <= 0; flappy_W(51, 455) <= 0; flappy_W(51, 456) <= 0; flappy_W(51, 457) <= 0; flappy_W(51, 458) <= 0; flappy_W(51, 459) <= 0; flappy_W(51, 460) <= 0; flappy_W(51, 461) <= 0; flappy_W(51, 462) <= 0; flappy_W(51, 463) <= 0; flappy_W(51, 464) <= 0; flappy_W(51, 465) <= 0; flappy_W(51, 466) <= 0; flappy_W(51, 467) <= 0; flappy_W(51, 468) <= 1; flappy_W(51, 469) <= 1; flappy_W(51, 470) <= 1; flappy_W(51, 471) <= 1; flappy_W(51, 472) <= 1; flappy_W(51, 473) <= 1; flappy_W(51, 474) <= 1; flappy_W(51, 475) <= 1; flappy_W(51, 476) <= 1; flappy_W(51, 477) <= 1; flappy_W(51, 478) <= 1; flappy_W(51, 479) <= 1; flappy_W(51, 480) <= 0; flappy_W(51, 481) <= 0; flappy_W(51, 482) <= 0; flappy_W(51, 483) <= 0; flappy_W(51, 484) <= 0; flappy_W(51, 485) <= 0; flappy_W(51, 486) <= 0; flappy_W(51, 487) <= 0; flappy_W(51, 488) <= 0; flappy_W(51, 489) <= 0; flappy_W(51, 490) <= 0; flappy_W(51, 491) <= 0; flappy_W(51, 492) <= 0; flappy_W(51, 493) <= 0; flappy_W(51, 494) <= 0; flappy_W(51, 495) <= 0; flappy_W(51, 496) <= 0; flappy_W(51, 497) <= 0; flappy_W(51, 498) <= 0; flappy_W(51, 499) <= 0; flappy_W(51, 500) <= 0; flappy_W(51, 501) <= 0; flappy_W(51, 502) <= 0; flappy_W(51, 503) <= 0; flappy_W(51, 504) <= 0; flappy_W(51, 505) <= 0; flappy_W(51, 506) <= 0; flappy_W(51, 507) <= 0; flappy_W(51, 508) <= 0; flappy_W(51, 509) <= 0; flappy_W(51, 510) <= 1; flappy_W(51, 511) <= 1; flappy_W(51, 512) <= 1; flappy_W(51, 513) <= 1; flappy_W(51, 514) <= 1; flappy_W(51, 515) <= 1; flappy_W(51, 516) <= 1; flappy_W(51, 517) <= 1; flappy_W(51, 518) <= 1; flappy_W(51, 519) <= 1; flappy_W(51, 520) <= 1; flappy_W(51, 521) <= 1; flappy_W(51, 522) <= 0; flappy_W(51, 523) <= 0; flappy_W(51, 524) <= 0; flappy_W(51, 525) <= 0; flappy_W(51, 526) <= 0; flappy_W(51, 527) <= 0; flappy_W(51, 528) <= 0; flappy_W(51, 529) <= 0; flappy_W(51, 530) <= 0; flappy_W(51, 531) <= 0; flappy_W(51, 532) <= 0; flappy_W(51, 533) <= 0; flappy_W(51, 534) <= 1; flappy_W(51, 535) <= 1; flappy_W(51, 536) <= 1; flappy_W(51, 537) <= 1; flappy_W(51, 538) <= 1; flappy_W(51, 539) <= 1; flappy_W(51, 540) <= 1; flappy_W(51, 541) <= 1; flappy_W(51, 542) <= 1; flappy_W(51, 543) <= 1; flappy_W(51, 544) <= 1; flappy_W(51, 545) <= 1; flappy_W(51, 546) <= 0; flappy_W(51, 547) <= 0; flappy_W(51, 548) <= 0; flappy_W(51, 549) <= 0; flappy_W(51, 550) <= 0; flappy_W(51, 551) <= 0; flappy_W(51, 552) <= 0; flappy_W(51, 553) <= 0; flappy_W(51, 554) <= 0; flappy_W(51, 555) <= 0; flappy_W(51, 556) <= 0; flappy_W(51, 557) <= 0; flappy_W(51, 558) <= 0; flappy_W(51, 559) <= 0; flappy_W(51, 560) <= 0; flappy_W(51, 561) <= 0; flappy_W(51, 562) <= 0; flappy_W(51, 563) <= 0; flappy_W(51, 564) <= 1; flappy_W(51, 565) <= 1; flappy_W(51, 566) <= 1; flappy_W(51, 567) <= 1; flappy_W(51, 568) <= 1; flappy_W(51, 569) <= 1; flappy_W(51, 570) <= 1; flappy_W(51, 571) <= 1; flappy_W(51, 572) <= 1; flappy_W(51, 573) <= 1; flappy_W(51, 574) <= 1; flappy_W(51, 575) <= 1; flappy_W(51, 576) <= 0; flappy_W(51, 577) <= 0; flappy_W(51, 578) <= 0; flappy_W(51, 579) <= 0; flappy_W(51, 580) <= 0; flappy_W(51, 581) <= 0; flappy_W(51, 582) <= 1; flappy_W(51, 583) <= 1; flappy_W(51, 584) <= 1; flappy_W(51, 585) <= 1; flappy_W(51, 586) <= 1; flappy_W(51, 587) <= 1; flappy_W(51, 588) <= 1; flappy_W(51, 589) <= 1; flappy_W(51, 590) <= 1; flappy_W(51, 591) <= 1; flappy_W(51, 592) <= 1; flappy_W(51, 593) <= 1; 
flappy_W(52, 0) <= 0; flappy_W(52, 1) <= 0; flappy_W(52, 2) <= 0; flappy_W(52, 3) <= 0; flappy_W(52, 4) <= 0; flappy_W(52, 5) <= 0; flappy_W(52, 6) <= 1; flappy_W(52, 7) <= 1; flappy_W(52, 8) <= 1; flappy_W(52, 9) <= 1; flappy_W(52, 10) <= 1; flappy_W(52, 11) <= 1; flappy_W(52, 12) <= 1; flappy_W(52, 13) <= 1; flappy_W(52, 14) <= 1; flappy_W(52, 15) <= 1; flappy_W(52, 16) <= 1; flappy_W(52, 17) <= 1; flappy_W(52, 18) <= 0; flappy_W(52, 19) <= 0; flappy_W(52, 20) <= 0; flappy_W(52, 21) <= 0; flappy_W(52, 22) <= 0; flappy_W(52, 23) <= 0; flappy_W(52, 24) <= 0; flappy_W(52, 25) <= 0; flappy_W(52, 26) <= 0; flappy_W(52, 27) <= 0; flappy_W(52, 28) <= 0; flappy_W(52, 29) <= 0; flappy_W(52, 30) <= 0; flappy_W(52, 31) <= 0; flappy_W(52, 32) <= 0; flappy_W(52, 33) <= 0; flappy_W(52, 34) <= 0; flappy_W(52, 35) <= 0; flappy_W(52, 36) <= 0; flappy_W(52, 37) <= 0; flappy_W(52, 38) <= 0; flappy_W(52, 39) <= 0; flappy_W(52, 40) <= 0; flappy_W(52, 41) <= 0; flappy_W(52, 42) <= 0; flappy_W(52, 43) <= 0; flappy_W(52, 44) <= 0; flappy_W(52, 45) <= 0; flappy_W(52, 46) <= 0; flappy_W(52, 47) <= 0; flappy_W(52, 48) <= 0; flappy_W(52, 49) <= 0; flappy_W(52, 50) <= 0; flappy_W(52, 51) <= 0; flappy_W(52, 52) <= 0; flappy_W(52, 53) <= 0; flappy_W(52, 54) <= 0; flappy_W(52, 55) <= 0; flappy_W(52, 56) <= 0; flappy_W(52, 57) <= 0; flappy_W(52, 58) <= 0; flappy_W(52, 59) <= 0; flappy_W(52, 60) <= 1; flappy_W(52, 61) <= 1; flappy_W(52, 62) <= 1; flappy_W(52, 63) <= 1; flappy_W(52, 64) <= 1; flappy_W(52, 65) <= 1; flappy_W(52, 66) <= 1; flappy_W(52, 67) <= 1; flappy_W(52, 68) <= 1; flappy_W(52, 69) <= 1; flappy_W(52, 70) <= 1; flappy_W(52, 71) <= 1; flappy_W(52, 72) <= 0; flappy_W(52, 73) <= 0; flappy_W(52, 74) <= 0; flappy_W(52, 75) <= 0; flappy_W(52, 76) <= 0; flappy_W(52, 77) <= 0; flappy_W(52, 78) <= 0; flappy_W(52, 79) <= 0; flappy_W(52, 80) <= 0; flappy_W(52, 81) <= 0; flappy_W(52, 82) <= 0; flappy_W(52, 83) <= 0; flappy_W(52, 84) <= 1; flappy_W(52, 85) <= 1; flappy_W(52, 86) <= 1; flappy_W(52, 87) <= 1; flappy_W(52, 88) <= 1; flappy_W(52, 89) <= 1; flappy_W(52, 90) <= 1; flappy_W(52, 91) <= 1; flappy_W(52, 92) <= 1; flappy_W(52, 93) <= 1; flappy_W(52, 94) <= 1; flappy_W(52, 95) <= 1; flappy_W(52, 96) <= 0; flappy_W(52, 97) <= 0; flappy_W(52, 98) <= 0; flappy_W(52, 99) <= 0; flappy_W(52, 100) <= 0; flappy_W(52, 101) <= 0; flappy_W(52, 102) <= 0; flappy_W(52, 103) <= 0; flappy_W(52, 104) <= 0; flappy_W(52, 105) <= 0; flappy_W(52, 106) <= 0; flappy_W(52, 107) <= 0; flappy_W(52, 108) <= 1; flappy_W(52, 109) <= 1; flappy_W(52, 110) <= 1; flappy_W(52, 111) <= 1; flappy_W(52, 112) <= 1; flappy_W(52, 113) <= 1; flappy_W(52, 114) <= 1; flappy_W(52, 115) <= 1; flappy_W(52, 116) <= 1; flappy_W(52, 117) <= 1; flappy_W(52, 118) <= 1; flappy_W(52, 119) <= 1; flappy_W(52, 120) <= 0; flappy_W(52, 121) <= 0; flappy_W(52, 122) <= 0; flappy_W(52, 123) <= 0; flappy_W(52, 124) <= 0; flappy_W(52, 125) <= 0; flappy_W(52, 126) <= 0; flappy_W(52, 127) <= 0; flappy_W(52, 128) <= 0; flappy_W(52, 129) <= 0; flappy_W(52, 130) <= 0; flappy_W(52, 131) <= 0; flappy_W(52, 132) <= 0; flappy_W(52, 133) <= 0; flappy_W(52, 134) <= 0; flappy_W(52, 135) <= 0; flappy_W(52, 136) <= 0; flappy_W(52, 137) <= 0; flappy_W(52, 138) <= 1; flappy_W(52, 139) <= 1; flappy_W(52, 140) <= 1; flappy_W(52, 141) <= 1; flappy_W(52, 142) <= 1; flappy_W(52, 143) <= 1; flappy_W(52, 144) <= 1; flappy_W(52, 145) <= 1; flappy_W(52, 146) <= 1; flappy_W(52, 147) <= 1; flappy_W(52, 148) <= 1; flappy_W(52, 149) <= 1; flappy_W(52, 150) <= 0; flappy_W(52, 151) <= 0; flappy_W(52, 152) <= 0; flappy_W(52, 153) <= 0; flappy_W(52, 154) <= 0; flappy_W(52, 155) <= 0; flappy_W(52, 156) <= 0; flappy_W(52, 157) <= 0; flappy_W(52, 158) <= 0; flappy_W(52, 159) <= 0; flappy_W(52, 160) <= 0; flappy_W(52, 161) <= 0; flappy_W(52, 162) <= 0; flappy_W(52, 163) <= 0; flappy_W(52, 164) <= 0; flappy_W(52, 165) <= 0; flappy_W(52, 166) <= 0; flappy_W(52, 167) <= 0; flappy_W(52, 168) <= 1; flappy_W(52, 169) <= 1; flappy_W(52, 170) <= 1; flappy_W(52, 171) <= 1; flappy_W(52, 172) <= 1; flappy_W(52, 173) <= 1; flappy_W(52, 174) <= 1; flappy_W(52, 175) <= 1; flappy_W(52, 176) <= 1; flappy_W(52, 177) <= 1; flappy_W(52, 178) <= 1; flappy_W(52, 179) <= 1; flappy_W(52, 180) <= 0; flappy_W(52, 181) <= 0; flappy_W(52, 182) <= 0; flappy_W(52, 183) <= 0; flappy_W(52, 184) <= 0; flappy_W(52, 185) <= 0; flappy_W(52, 186) <= 0; flappy_W(52, 187) <= 0; flappy_W(52, 188) <= 0; flappy_W(52, 189) <= 0; flappy_W(52, 190) <= 0; flappy_W(52, 191) <= 0; flappy_W(52, 192) <= 0; flappy_W(52, 193) <= 0; flappy_W(52, 194) <= 0; flappy_W(52, 195) <= 0; flappy_W(52, 196) <= 0; flappy_W(52, 197) <= 0; flappy_W(52, 198) <= 0; flappy_W(52, 199) <= 0; flappy_W(52, 200) <= 0; flappy_W(52, 201) <= 0; flappy_W(52, 202) <= 0; flappy_W(52, 203) <= 0; flappy_W(52, 204) <= 0; flappy_W(52, 205) <= 0; flappy_W(52, 206) <= 0; flappy_W(52, 207) <= 0; flappy_W(52, 208) <= 0; flappy_W(52, 209) <= 0; flappy_W(52, 210) <= 0; flappy_W(52, 211) <= 0; flappy_W(52, 212) <= 0; flappy_W(52, 213) <= 0; flappy_W(52, 214) <= 0; flappy_W(52, 215) <= 0; flappy_W(52, 216) <= 0; flappy_W(52, 217) <= 0; flappy_W(52, 218) <= 0; flappy_W(52, 219) <= 0; flappy_W(52, 220) <= 0; flappy_W(52, 221) <= 0; flappy_W(52, 222) <= 1; flappy_W(52, 223) <= 1; flappy_W(52, 224) <= 1; flappy_W(52, 225) <= 1; flappy_W(52, 226) <= 1; flappy_W(52, 227) <= 1; flappy_W(52, 228) <= 1; flappy_W(52, 229) <= 1; flappy_W(52, 230) <= 1; flappy_W(52, 231) <= 1; flappy_W(52, 232) <= 1; flappy_W(52, 233) <= 1; flappy_W(52, 234) <= 0; flappy_W(52, 235) <= 0; flappy_W(52, 236) <= 0; flappy_W(52, 237) <= 0; flappy_W(52, 238) <= 0; flappy_W(52, 239) <= 0; flappy_W(52, 240) <= 0; flappy_W(52, 241) <= 0; flappy_W(52, 242) <= 0; flappy_W(52, 243) <= 0; flappy_W(52, 244) <= 0; flappy_W(52, 245) <= 0; flappy_W(52, 246) <= 0; flappy_W(52, 247) <= 0; flappy_W(52, 248) <= 0; flappy_W(52, 249) <= 0; flappy_W(52, 250) <= 0; flappy_W(52, 251) <= 0; flappy_W(52, 252) <= 0; flappy_W(52, 253) <= 0; flappy_W(52, 254) <= 0; flappy_W(52, 255) <= 0; flappy_W(52, 256) <= 0; flappy_W(52, 257) <= 0; flappy_W(52, 258) <= 0; flappy_W(52, 259) <= 0; flappy_W(52, 260) <= 0; flappy_W(52, 261) <= 0; flappy_W(52, 262) <= 0; flappy_W(52, 263) <= 0; flappy_W(52, 264) <= 0; flappy_W(52, 265) <= 0; flappy_W(52, 266) <= 0; flappy_W(52, 267) <= 0; flappy_W(52, 268) <= 0; flappy_W(52, 269) <= 0; flappy_W(52, 270) <= 0; flappy_W(52, 271) <= 0; flappy_W(52, 272) <= 0; flappy_W(52, 273) <= 0; flappy_W(52, 274) <= 0; flappy_W(52, 275) <= 0; flappy_W(52, 276) <= 0; flappy_W(52, 277) <= 0; flappy_W(52, 278) <= 0; flappy_W(52, 279) <= 0; flappy_W(52, 280) <= 0; flappy_W(52, 281) <= 0; flappy_W(52, 282) <= 0; flappy_W(52, 283) <= 0; flappy_W(52, 284) <= 0; flappy_W(52, 285) <= 0; flappy_W(52, 286) <= 0; flappy_W(52, 287) <= 0; flappy_W(52, 288) <= 1; flappy_W(52, 289) <= 1; flappy_W(52, 290) <= 1; flappy_W(52, 291) <= 1; flappy_W(52, 292) <= 1; flappy_W(52, 293) <= 1; flappy_W(52, 294) <= 1; flappy_W(52, 295) <= 1; flappy_W(52, 296) <= 1; flappy_W(52, 297) <= 1; flappy_W(52, 298) <= 1; flappy_W(52, 299) <= 1; flappy_W(52, 300) <= 0; flappy_W(52, 301) <= 0; flappy_W(52, 302) <= 0; flappy_W(52, 303) <= 0; flappy_W(52, 304) <= 0; flappy_W(52, 305) <= 0; flappy_W(52, 306) <= 0; flappy_W(52, 307) <= 0; flappy_W(52, 308) <= 0; flappy_W(52, 309) <= 0; flappy_W(52, 310) <= 0; flappy_W(52, 311) <= 0; flappy_W(52, 312) <= 0; flappy_W(52, 313) <= 0; flappy_W(52, 314) <= 0; flappy_W(52, 315) <= 0; flappy_W(52, 316) <= 0; flappy_W(52, 317) <= 0; flappy_W(52, 318) <= 0; flappy_W(52, 319) <= 0; flappy_W(52, 320) <= 0; flappy_W(52, 321) <= 0; flappy_W(52, 322) <= 0; flappy_W(52, 323) <= 0; flappy_W(52, 324) <= 0; flappy_W(52, 325) <= 0; flappy_W(52, 326) <= 0; flappy_W(52, 327) <= 0; flappy_W(52, 328) <= 0; flappy_W(52, 329) <= 0; flappy_W(52, 330) <= 0; flappy_W(52, 331) <= 0; flappy_W(52, 332) <= 0; flappy_W(52, 333) <= 0; flappy_W(52, 334) <= 0; flappy_W(52, 335) <= 0; flappy_W(52, 336) <= 0; flappy_W(52, 337) <= 0; flappy_W(52, 338) <= 0; flappy_W(52, 339) <= 0; flappy_W(52, 340) <= 0; flappy_W(52, 341) <= 0; flappy_W(52, 342) <= 0; flappy_W(52, 343) <= 0; flappy_W(52, 344) <= 0; flappy_W(52, 345) <= 0; flappy_W(52, 346) <= 0; flappy_W(52, 347) <= 0; flappy_W(52, 348) <= 0; flappy_W(52, 349) <= 0; flappy_W(52, 350) <= 0; flappy_W(52, 351) <= 0; flappy_W(52, 352) <= 0; flappy_W(52, 353) <= 0; flappy_W(52, 354) <= 0; flappy_W(52, 355) <= 0; flappy_W(52, 356) <= 0; flappy_W(52, 357) <= 0; flappy_W(52, 358) <= 0; flappy_W(52, 359) <= 0; flappy_W(52, 360) <= 0; flappy_W(52, 361) <= 0; flappy_W(52, 362) <= 0; flappy_W(52, 363) <= 0; flappy_W(52, 364) <= 0; flappy_W(52, 365) <= 0; flappy_W(52, 366) <= 0; flappy_W(52, 367) <= 0; flappy_W(52, 368) <= 0; flappy_W(52, 369) <= 0; flappy_W(52, 370) <= 0; flappy_W(52, 371) <= 0; flappy_W(52, 372) <= 0; flappy_W(52, 373) <= 0; flappy_W(52, 374) <= 0; flappy_W(52, 375) <= 0; flappy_W(52, 376) <= 0; flappy_W(52, 377) <= 0; flappy_W(52, 378) <= 0; flappy_W(52, 379) <= 0; flappy_W(52, 380) <= 0; flappy_W(52, 381) <= 0; flappy_W(52, 382) <= 0; flappy_W(52, 383) <= 0; flappy_W(52, 384) <= 0; flappy_W(52, 385) <= 0; flappy_W(52, 386) <= 0; flappy_W(52, 387) <= 0; flappy_W(52, 388) <= 0; flappy_W(52, 389) <= 0; flappy_W(52, 390) <= 0; flappy_W(52, 391) <= 0; flappy_W(52, 392) <= 0; flappy_W(52, 393) <= 0; flappy_W(52, 394) <= 0; flappy_W(52, 395) <= 0; flappy_W(52, 396) <= 0; flappy_W(52, 397) <= 0; flappy_W(52, 398) <= 0; flappy_W(52, 399) <= 0; flappy_W(52, 400) <= 0; flappy_W(52, 401) <= 0; flappy_W(52, 402) <= 1; flappy_W(52, 403) <= 1; flappy_W(52, 404) <= 1; flappy_W(52, 405) <= 1; flappy_W(52, 406) <= 1; flappy_W(52, 407) <= 1; flappy_W(52, 408) <= 1; flappy_W(52, 409) <= 1; flappy_W(52, 410) <= 1; flappy_W(52, 411) <= 1; flappy_W(52, 412) <= 1; flappy_W(52, 413) <= 1; flappy_W(52, 414) <= 0; flappy_W(52, 415) <= 0; flappy_W(52, 416) <= 0; flappy_W(52, 417) <= 0; flappy_W(52, 418) <= 0; flappy_W(52, 419) <= 0; flappy_W(52, 420) <= 0; flappy_W(52, 421) <= 0; flappy_W(52, 422) <= 0; flappy_W(52, 423) <= 0; flappy_W(52, 424) <= 0; flappy_W(52, 425) <= 0; flappy_W(52, 426) <= 1; flappy_W(52, 427) <= 1; flappy_W(52, 428) <= 1; flappy_W(52, 429) <= 1; flappy_W(52, 430) <= 1; flappy_W(52, 431) <= 1; flappy_W(52, 432) <= 1; flappy_W(52, 433) <= 1; flappy_W(52, 434) <= 1; flappy_W(52, 435) <= 1; flappy_W(52, 436) <= 1; flappy_W(52, 437) <= 1; flappy_W(52, 438) <= 0; flappy_W(52, 439) <= 0; flappy_W(52, 440) <= 0; flappy_W(52, 441) <= 0; flappy_W(52, 442) <= 0; flappy_W(52, 443) <= 0; flappy_W(52, 444) <= 0; flappy_W(52, 445) <= 0; flappy_W(52, 446) <= 0; flappy_W(52, 447) <= 0; flappy_W(52, 448) <= 0; flappy_W(52, 449) <= 0; flappy_W(52, 450) <= 0; flappy_W(52, 451) <= 0; flappy_W(52, 452) <= 0; flappy_W(52, 453) <= 0; flappy_W(52, 454) <= 0; flappy_W(52, 455) <= 0; flappy_W(52, 456) <= 0; flappy_W(52, 457) <= 0; flappy_W(52, 458) <= 0; flappy_W(52, 459) <= 0; flappy_W(52, 460) <= 0; flappy_W(52, 461) <= 0; flappy_W(52, 462) <= 0; flappy_W(52, 463) <= 0; flappy_W(52, 464) <= 0; flappy_W(52, 465) <= 0; flappy_W(52, 466) <= 0; flappy_W(52, 467) <= 0; flappy_W(52, 468) <= 1; flappy_W(52, 469) <= 1; flappy_W(52, 470) <= 1; flappy_W(52, 471) <= 1; flappy_W(52, 472) <= 1; flappy_W(52, 473) <= 1; flappy_W(52, 474) <= 1; flappy_W(52, 475) <= 1; flappy_W(52, 476) <= 1; flappy_W(52, 477) <= 1; flappy_W(52, 478) <= 1; flappy_W(52, 479) <= 1; flappy_W(52, 480) <= 0; flappy_W(52, 481) <= 0; flappy_W(52, 482) <= 0; flappy_W(52, 483) <= 0; flappy_W(52, 484) <= 0; flappy_W(52, 485) <= 0; flappy_W(52, 486) <= 0; flappy_W(52, 487) <= 0; flappy_W(52, 488) <= 0; flappy_W(52, 489) <= 0; flappy_W(52, 490) <= 0; flappy_W(52, 491) <= 0; flappy_W(52, 492) <= 0; flappy_W(52, 493) <= 0; flappy_W(52, 494) <= 0; flappy_W(52, 495) <= 0; flappy_W(52, 496) <= 0; flappy_W(52, 497) <= 0; flappy_W(52, 498) <= 0; flappy_W(52, 499) <= 0; flappy_W(52, 500) <= 0; flappy_W(52, 501) <= 0; flappy_W(52, 502) <= 0; flappy_W(52, 503) <= 0; flappy_W(52, 504) <= 0; flappy_W(52, 505) <= 0; flappy_W(52, 506) <= 0; flappy_W(52, 507) <= 0; flappy_W(52, 508) <= 0; flappy_W(52, 509) <= 0; flappy_W(52, 510) <= 1; flappy_W(52, 511) <= 1; flappy_W(52, 512) <= 1; flappy_W(52, 513) <= 1; flappy_W(52, 514) <= 1; flappy_W(52, 515) <= 1; flappy_W(52, 516) <= 1; flappy_W(52, 517) <= 1; flappy_W(52, 518) <= 1; flappy_W(52, 519) <= 1; flappy_W(52, 520) <= 1; flappy_W(52, 521) <= 1; flappy_W(52, 522) <= 0; flappy_W(52, 523) <= 0; flappy_W(52, 524) <= 0; flappy_W(52, 525) <= 0; flappy_W(52, 526) <= 0; flappy_W(52, 527) <= 0; flappy_W(52, 528) <= 0; flappy_W(52, 529) <= 0; flappy_W(52, 530) <= 0; flappy_W(52, 531) <= 0; flappy_W(52, 532) <= 0; flappy_W(52, 533) <= 0; flappy_W(52, 534) <= 1; flappy_W(52, 535) <= 1; flappy_W(52, 536) <= 1; flappy_W(52, 537) <= 1; flappy_W(52, 538) <= 1; flappy_W(52, 539) <= 1; flappy_W(52, 540) <= 1; flappy_W(52, 541) <= 1; flappy_W(52, 542) <= 1; flappy_W(52, 543) <= 1; flappy_W(52, 544) <= 1; flappy_W(52, 545) <= 1; flappy_W(52, 546) <= 0; flappy_W(52, 547) <= 0; flappy_W(52, 548) <= 0; flappy_W(52, 549) <= 0; flappy_W(52, 550) <= 0; flappy_W(52, 551) <= 0; flappy_W(52, 552) <= 0; flappy_W(52, 553) <= 0; flappy_W(52, 554) <= 0; flappy_W(52, 555) <= 0; flappy_W(52, 556) <= 0; flappy_W(52, 557) <= 0; flappy_W(52, 558) <= 0; flappy_W(52, 559) <= 0; flappy_W(52, 560) <= 0; flappy_W(52, 561) <= 0; flappy_W(52, 562) <= 0; flappy_W(52, 563) <= 0; flappy_W(52, 564) <= 1; flappy_W(52, 565) <= 1; flappy_W(52, 566) <= 1; flappy_W(52, 567) <= 1; flappy_W(52, 568) <= 1; flappy_W(52, 569) <= 1; flappy_W(52, 570) <= 1; flappy_W(52, 571) <= 1; flappy_W(52, 572) <= 1; flappy_W(52, 573) <= 1; flappy_W(52, 574) <= 1; flappy_W(52, 575) <= 1; flappy_W(52, 576) <= 0; flappy_W(52, 577) <= 0; flappy_W(52, 578) <= 0; flappy_W(52, 579) <= 0; flappy_W(52, 580) <= 0; flappy_W(52, 581) <= 0; flappy_W(52, 582) <= 1; flappy_W(52, 583) <= 1; flappy_W(52, 584) <= 1; flappy_W(52, 585) <= 1; flappy_W(52, 586) <= 1; flappy_W(52, 587) <= 1; flappy_W(52, 588) <= 1; flappy_W(52, 589) <= 1; flappy_W(52, 590) <= 1; flappy_W(52, 591) <= 1; flappy_W(52, 592) <= 1; flappy_W(52, 593) <= 1; 
flappy_W(53, 0) <= 0; flappy_W(53, 1) <= 0; flappy_W(53, 2) <= 0; flappy_W(53, 3) <= 0; flappy_W(53, 4) <= 0; flappy_W(53, 5) <= 0; flappy_W(53, 6) <= 1; flappy_W(53, 7) <= 1; flappy_W(53, 8) <= 1; flappy_W(53, 9) <= 1; flappy_W(53, 10) <= 1; flappy_W(53, 11) <= 1; flappy_W(53, 12) <= 1; flappy_W(53, 13) <= 1; flappy_W(53, 14) <= 1; flappy_W(53, 15) <= 1; flappy_W(53, 16) <= 1; flappy_W(53, 17) <= 1; flappy_W(53, 18) <= 0; flappy_W(53, 19) <= 0; flappy_W(53, 20) <= 0; flappy_W(53, 21) <= 0; flappy_W(53, 22) <= 0; flappy_W(53, 23) <= 0; flappy_W(53, 24) <= 0; flappy_W(53, 25) <= 0; flappy_W(53, 26) <= 0; flappy_W(53, 27) <= 0; flappy_W(53, 28) <= 0; flappy_W(53, 29) <= 0; flappy_W(53, 30) <= 0; flappy_W(53, 31) <= 0; flappy_W(53, 32) <= 0; flappy_W(53, 33) <= 0; flappy_W(53, 34) <= 0; flappy_W(53, 35) <= 0; flappy_W(53, 36) <= 0; flappy_W(53, 37) <= 0; flappy_W(53, 38) <= 0; flappy_W(53, 39) <= 0; flappy_W(53, 40) <= 0; flappy_W(53, 41) <= 0; flappy_W(53, 42) <= 0; flappy_W(53, 43) <= 0; flappy_W(53, 44) <= 0; flappy_W(53, 45) <= 0; flappy_W(53, 46) <= 0; flappy_W(53, 47) <= 0; flappy_W(53, 48) <= 0; flappy_W(53, 49) <= 0; flappy_W(53, 50) <= 0; flappy_W(53, 51) <= 0; flappy_W(53, 52) <= 0; flappy_W(53, 53) <= 0; flappy_W(53, 54) <= 0; flappy_W(53, 55) <= 0; flappy_W(53, 56) <= 0; flappy_W(53, 57) <= 0; flappy_W(53, 58) <= 0; flappy_W(53, 59) <= 0; flappy_W(53, 60) <= 1; flappy_W(53, 61) <= 1; flappy_W(53, 62) <= 1; flappy_W(53, 63) <= 1; flappy_W(53, 64) <= 1; flappy_W(53, 65) <= 1; flappy_W(53, 66) <= 1; flappy_W(53, 67) <= 1; flappy_W(53, 68) <= 1; flappy_W(53, 69) <= 1; flappy_W(53, 70) <= 1; flappy_W(53, 71) <= 1; flappy_W(53, 72) <= 0; flappy_W(53, 73) <= 0; flappy_W(53, 74) <= 0; flappy_W(53, 75) <= 0; flappy_W(53, 76) <= 0; flappy_W(53, 77) <= 0; flappy_W(53, 78) <= 0; flappy_W(53, 79) <= 0; flappy_W(53, 80) <= 0; flappy_W(53, 81) <= 0; flappy_W(53, 82) <= 0; flappy_W(53, 83) <= 0; flappy_W(53, 84) <= 1; flappy_W(53, 85) <= 1; flappy_W(53, 86) <= 1; flappy_W(53, 87) <= 1; flappy_W(53, 88) <= 1; flappy_W(53, 89) <= 1; flappy_W(53, 90) <= 1; flappy_W(53, 91) <= 1; flappy_W(53, 92) <= 1; flappy_W(53, 93) <= 1; flappy_W(53, 94) <= 1; flappy_W(53, 95) <= 1; flappy_W(53, 96) <= 0; flappy_W(53, 97) <= 0; flappy_W(53, 98) <= 0; flappy_W(53, 99) <= 0; flappy_W(53, 100) <= 0; flappy_W(53, 101) <= 0; flappy_W(53, 102) <= 0; flappy_W(53, 103) <= 0; flappy_W(53, 104) <= 0; flappy_W(53, 105) <= 0; flappy_W(53, 106) <= 0; flappy_W(53, 107) <= 0; flappy_W(53, 108) <= 1; flappy_W(53, 109) <= 1; flappy_W(53, 110) <= 1; flappy_W(53, 111) <= 1; flappy_W(53, 112) <= 1; flappy_W(53, 113) <= 1; flappy_W(53, 114) <= 1; flappy_W(53, 115) <= 1; flappy_W(53, 116) <= 1; flappy_W(53, 117) <= 1; flappy_W(53, 118) <= 1; flappy_W(53, 119) <= 1; flappy_W(53, 120) <= 0; flappy_W(53, 121) <= 0; flappy_W(53, 122) <= 0; flappy_W(53, 123) <= 0; flappy_W(53, 124) <= 0; flappy_W(53, 125) <= 0; flappy_W(53, 126) <= 0; flappy_W(53, 127) <= 0; flappy_W(53, 128) <= 0; flappy_W(53, 129) <= 0; flappy_W(53, 130) <= 0; flappy_W(53, 131) <= 0; flappy_W(53, 132) <= 0; flappy_W(53, 133) <= 0; flappy_W(53, 134) <= 0; flappy_W(53, 135) <= 0; flappy_W(53, 136) <= 0; flappy_W(53, 137) <= 0; flappy_W(53, 138) <= 1; flappy_W(53, 139) <= 1; flappy_W(53, 140) <= 1; flappy_W(53, 141) <= 1; flappy_W(53, 142) <= 1; flappy_W(53, 143) <= 1; flappy_W(53, 144) <= 1; flappy_W(53, 145) <= 1; flappy_W(53, 146) <= 1; flappy_W(53, 147) <= 1; flappy_W(53, 148) <= 1; flappy_W(53, 149) <= 1; flappy_W(53, 150) <= 0; flappy_W(53, 151) <= 0; flappy_W(53, 152) <= 0; flappy_W(53, 153) <= 0; flappy_W(53, 154) <= 0; flappy_W(53, 155) <= 0; flappy_W(53, 156) <= 0; flappy_W(53, 157) <= 0; flappy_W(53, 158) <= 0; flappy_W(53, 159) <= 0; flappy_W(53, 160) <= 0; flappy_W(53, 161) <= 0; flappy_W(53, 162) <= 0; flappy_W(53, 163) <= 0; flappy_W(53, 164) <= 0; flappy_W(53, 165) <= 0; flappy_W(53, 166) <= 0; flappy_W(53, 167) <= 0; flappy_W(53, 168) <= 1; flappy_W(53, 169) <= 1; flappy_W(53, 170) <= 1; flappy_W(53, 171) <= 1; flappy_W(53, 172) <= 1; flappy_W(53, 173) <= 1; flappy_W(53, 174) <= 1; flappy_W(53, 175) <= 1; flappy_W(53, 176) <= 1; flappy_W(53, 177) <= 1; flappy_W(53, 178) <= 1; flappy_W(53, 179) <= 1; flappy_W(53, 180) <= 0; flappy_W(53, 181) <= 0; flappy_W(53, 182) <= 0; flappy_W(53, 183) <= 0; flappy_W(53, 184) <= 0; flappy_W(53, 185) <= 0; flappy_W(53, 186) <= 0; flappy_W(53, 187) <= 0; flappy_W(53, 188) <= 0; flappy_W(53, 189) <= 0; flappy_W(53, 190) <= 0; flappy_W(53, 191) <= 0; flappy_W(53, 192) <= 0; flappy_W(53, 193) <= 0; flappy_W(53, 194) <= 0; flappy_W(53, 195) <= 0; flappy_W(53, 196) <= 0; flappy_W(53, 197) <= 0; flappy_W(53, 198) <= 0; flappy_W(53, 199) <= 0; flappy_W(53, 200) <= 0; flappy_W(53, 201) <= 0; flappy_W(53, 202) <= 0; flappy_W(53, 203) <= 0; flappy_W(53, 204) <= 0; flappy_W(53, 205) <= 0; flappy_W(53, 206) <= 0; flappy_W(53, 207) <= 0; flappy_W(53, 208) <= 0; flappy_W(53, 209) <= 0; flappy_W(53, 210) <= 0; flappy_W(53, 211) <= 0; flappy_W(53, 212) <= 0; flappy_W(53, 213) <= 0; flappy_W(53, 214) <= 0; flappy_W(53, 215) <= 0; flappy_W(53, 216) <= 0; flappy_W(53, 217) <= 0; flappy_W(53, 218) <= 0; flappy_W(53, 219) <= 0; flappy_W(53, 220) <= 0; flappy_W(53, 221) <= 0; flappy_W(53, 222) <= 1; flappy_W(53, 223) <= 1; flappy_W(53, 224) <= 1; flappy_W(53, 225) <= 1; flappy_W(53, 226) <= 1; flappy_W(53, 227) <= 1; flappy_W(53, 228) <= 1; flappy_W(53, 229) <= 1; flappy_W(53, 230) <= 1; flappy_W(53, 231) <= 1; flappy_W(53, 232) <= 1; flappy_W(53, 233) <= 1; flappy_W(53, 234) <= 0; flappy_W(53, 235) <= 0; flappy_W(53, 236) <= 0; flappy_W(53, 237) <= 0; flappy_W(53, 238) <= 0; flappy_W(53, 239) <= 0; flappy_W(53, 240) <= 0; flappy_W(53, 241) <= 0; flappy_W(53, 242) <= 0; flappy_W(53, 243) <= 0; flappy_W(53, 244) <= 0; flappy_W(53, 245) <= 0; flappy_W(53, 246) <= 0; flappy_W(53, 247) <= 0; flappy_W(53, 248) <= 0; flappy_W(53, 249) <= 0; flappy_W(53, 250) <= 0; flappy_W(53, 251) <= 0; flappy_W(53, 252) <= 0; flappy_W(53, 253) <= 0; flappy_W(53, 254) <= 0; flappy_W(53, 255) <= 0; flappy_W(53, 256) <= 0; flappy_W(53, 257) <= 0; flappy_W(53, 258) <= 0; flappy_W(53, 259) <= 0; flappy_W(53, 260) <= 0; flappy_W(53, 261) <= 0; flappy_W(53, 262) <= 0; flappy_W(53, 263) <= 0; flappy_W(53, 264) <= 0; flappy_W(53, 265) <= 0; flappy_W(53, 266) <= 0; flappy_W(53, 267) <= 0; flappy_W(53, 268) <= 0; flappy_W(53, 269) <= 0; flappy_W(53, 270) <= 0; flappy_W(53, 271) <= 0; flappy_W(53, 272) <= 0; flappy_W(53, 273) <= 0; flappy_W(53, 274) <= 0; flappy_W(53, 275) <= 0; flappy_W(53, 276) <= 0; flappy_W(53, 277) <= 0; flappy_W(53, 278) <= 0; flappy_W(53, 279) <= 0; flappy_W(53, 280) <= 0; flappy_W(53, 281) <= 0; flappy_W(53, 282) <= 0; flappy_W(53, 283) <= 0; flappy_W(53, 284) <= 0; flappy_W(53, 285) <= 0; flappy_W(53, 286) <= 0; flappy_W(53, 287) <= 0; flappy_W(53, 288) <= 1; flappy_W(53, 289) <= 1; flappy_W(53, 290) <= 1; flappy_W(53, 291) <= 1; flappy_W(53, 292) <= 1; flappy_W(53, 293) <= 1; flappy_W(53, 294) <= 1; flappy_W(53, 295) <= 1; flappy_W(53, 296) <= 1; flappy_W(53, 297) <= 1; flappy_W(53, 298) <= 1; flappy_W(53, 299) <= 1; flappy_W(53, 300) <= 0; flappy_W(53, 301) <= 0; flappy_W(53, 302) <= 0; flappy_W(53, 303) <= 0; flappy_W(53, 304) <= 0; flappy_W(53, 305) <= 0; flappy_W(53, 306) <= 0; flappy_W(53, 307) <= 0; flappy_W(53, 308) <= 0; flappy_W(53, 309) <= 0; flappy_W(53, 310) <= 0; flappy_W(53, 311) <= 0; flappy_W(53, 312) <= 0; flappy_W(53, 313) <= 0; flappy_W(53, 314) <= 0; flappy_W(53, 315) <= 0; flappy_W(53, 316) <= 0; flappy_W(53, 317) <= 0; flappy_W(53, 318) <= 0; flappy_W(53, 319) <= 0; flappy_W(53, 320) <= 0; flappy_W(53, 321) <= 0; flappy_W(53, 322) <= 0; flappy_W(53, 323) <= 0; flappy_W(53, 324) <= 0; flappy_W(53, 325) <= 0; flappy_W(53, 326) <= 0; flappy_W(53, 327) <= 0; flappy_W(53, 328) <= 0; flappy_W(53, 329) <= 0; flappy_W(53, 330) <= 0; flappy_W(53, 331) <= 0; flappy_W(53, 332) <= 0; flappy_W(53, 333) <= 0; flappy_W(53, 334) <= 0; flappy_W(53, 335) <= 0; flappy_W(53, 336) <= 0; flappy_W(53, 337) <= 0; flappy_W(53, 338) <= 0; flappy_W(53, 339) <= 0; flappy_W(53, 340) <= 0; flappy_W(53, 341) <= 0; flappy_W(53, 342) <= 0; flappy_W(53, 343) <= 0; flappy_W(53, 344) <= 0; flappy_W(53, 345) <= 0; flappy_W(53, 346) <= 0; flappy_W(53, 347) <= 0; flappy_W(53, 348) <= 0; flappy_W(53, 349) <= 0; flappy_W(53, 350) <= 0; flappy_W(53, 351) <= 0; flappy_W(53, 352) <= 0; flappy_W(53, 353) <= 0; flappy_W(53, 354) <= 0; flappy_W(53, 355) <= 0; flappy_W(53, 356) <= 0; flappy_W(53, 357) <= 0; flappy_W(53, 358) <= 0; flappy_W(53, 359) <= 0; flappy_W(53, 360) <= 0; flappy_W(53, 361) <= 0; flappy_W(53, 362) <= 0; flappy_W(53, 363) <= 0; flappy_W(53, 364) <= 0; flappy_W(53, 365) <= 0; flappy_W(53, 366) <= 0; flappy_W(53, 367) <= 0; flappy_W(53, 368) <= 0; flappy_W(53, 369) <= 0; flappy_W(53, 370) <= 0; flappy_W(53, 371) <= 0; flappy_W(53, 372) <= 0; flappy_W(53, 373) <= 0; flappy_W(53, 374) <= 0; flappy_W(53, 375) <= 0; flappy_W(53, 376) <= 0; flappy_W(53, 377) <= 0; flappy_W(53, 378) <= 0; flappy_W(53, 379) <= 0; flappy_W(53, 380) <= 0; flappy_W(53, 381) <= 0; flappy_W(53, 382) <= 0; flappy_W(53, 383) <= 0; flappy_W(53, 384) <= 0; flappy_W(53, 385) <= 0; flappy_W(53, 386) <= 0; flappy_W(53, 387) <= 0; flappy_W(53, 388) <= 0; flappy_W(53, 389) <= 0; flappy_W(53, 390) <= 0; flappy_W(53, 391) <= 0; flappy_W(53, 392) <= 0; flappy_W(53, 393) <= 0; flappy_W(53, 394) <= 0; flappy_W(53, 395) <= 0; flappy_W(53, 396) <= 0; flappy_W(53, 397) <= 0; flappy_W(53, 398) <= 0; flappy_W(53, 399) <= 0; flappy_W(53, 400) <= 0; flappy_W(53, 401) <= 0; flappy_W(53, 402) <= 1; flappy_W(53, 403) <= 1; flappy_W(53, 404) <= 1; flappy_W(53, 405) <= 1; flappy_W(53, 406) <= 1; flappy_W(53, 407) <= 1; flappy_W(53, 408) <= 1; flappy_W(53, 409) <= 1; flappy_W(53, 410) <= 1; flappy_W(53, 411) <= 1; flappy_W(53, 412) <= 1; flappy_W(53, 413) <= 1; flappy_W(53, 414) <= 0; flappy_W(53, 415) <= 0; flappy_W(53, 416) <= 0; flappy_W(53, 417) <= 0; flappy_W(53, 418) <= 0; flappy_W(53, 419) <= 0; flappy_W(53, 420) <= 0; flappy_W(53, 421) <= 0; flappy_W(53, 422) <= 0; flappy_W(53, 423) <= 0; flappy_W(53, 424) <= 0; flappy_W(53, 425) <= 0; flappy_W(53, 426) <= 1; flappy_W(53, 427) <= 1; flappy_W(53, 428) <= 1; flappy_W(53, 429) <= 1; flappy_W(53, 430) <= 1; flappy_W(53, 431) <= 1; flappy_W(53, 432) <= 1; flappy_W(53, 433) <= 1; flappy_W(53, 434) <= 1; flappy_W(53, 435) <= 1; flappy_W(53, 436) <= 1; flappy_W(53, 437) <= 1; flappy_W(53, 438) <= 0; flappy_W(53, 439) <= 0; flappy_W(53, 440) <= 0; flappy_W(53, 441) <= 0; flappy_W(53, 442) <= 0; flappy_W(53, 443) <= 0; flappy_W(53, 444) <= 0; flappy_W(53, 445) <= 0; flappy_W(53, 446) <= 0; flappy_W(53, 447) <= 0; flappy_W(53, 448) <= 0; flappy_W(53, 449) <= 0; flappy_W(53, 450) <= 0; flappy_W(53, 451) <= 0; flappy_W(53, 452) <= 0; flappy_W(53, 453) <= 0; flappy_W(53, 454) <= 0; flappy_W(53, 455) <= 0; flappy_W(53, 456) <= 0; flappy_W(53, 457) <= 0; flappy_W(53, 458) <= 0; flappy_W(53, 459) <= 0; flappy_W(53, 460) <= 0; flappy_W(53, 461) <= 0; flappy_W(53, 462) <= 0; flappy_W(53, 463) <= 0; flappy_W(53, 464) <= 0; flappy_W(53, 465) <= 0; flappy_W(53, 466) <= 0; flappy_W(53, 467) <= 0; flappy_W(53, 468) <= 1; flappy_W(53, 469) <= 1; flappy_W(53, 470) <= 1; flappy_W(53, 471) <= 1; flappy_W(53, 472) <= 1; flappy_W(53, 473) <= 1; flappy_W(53, 474) <= 1; flappy_W(53, 475) <= 1; flappy_W(53, 476) <= 1; flappy_W(53, 477) <= 1; flappy_W(53, 478) <= 1; flappy_W(53, 479) <= 1; flappy_W(53, 480) <= 0; flappy_W(53, 481) <= 0; flappy_W(53, 482) <= 0; flappy_W(53, 483) <= 0; flappy_W(53, 484) <= 0; flappy_W(53, 485) <= 0; flappy_W(53, 486) <= 0; flappy_W(53, 487) <= 0; flappy_W(53, 488) <= 0; flappy_W(53, 489) <= 0; flappy_W(53, 490) <= 0; flappy_W(53, 491) <= 0; flappy_W(53, 492) <= 0; flappy_W(53, 493) <= 0; flappy_W(53, 494) <= 0; flappy_W(53, 495) <= 0; flappy_W(53, 496) <= 0; flappy_W(53, 497) <= 0; flappy_W(53, 498) <= 0; flappy_W(53, 499) <= 0; flappy_W(53, 500) <= 0; flappy_W(53, 501) <= 0; flappy_W(53, 502) <= 0; flappy_W(53, 503) <= 0; flappy_W(53, 504) <= 0; flappy_W(53, 505) <= 0; flappy_W(53, 506) <= 0; flappy_W(53, 507) <= 0; flappy_W(53, 508) <= 0; flappy_W(53, 509) <= 0; flappy_W(53, 510) <= 1; flappy_W(53, 511) <= 1; flappy_W(53, 512) <= 1; flappy_W(53, 513) <= 1; flappy_W(53, 514) <= 1; flappy_W(53, 515) <= 1; flappy_W(53, 516) <= 1; flappy_W(53, 517) <= 1; flappy_W(53, 518) <= 1; flappy_W(53, 519) <= 1; flappy_W(53, 520) <= 1; flappy_W(53, 521) <= 1; flappy_W(53, 522) <= 0; flappy_W(53, 523) <= 0; flappy_W(53, 524) <= 0; flappy_W(53, 525) <= 0; flappy_W(53, 526) <= 0; flappy_W(53, 527) <= 0; flappy_W(53, 528) <= 0; flappy_W(53, 529) <= 0; flappy_W(53, 530) <= 0; flappy_W(53, 531) <= 0; flappy_W(53, 532) <= 0; flappy_W(53, 533) <= 0; flappy_W(53, 534) <= 1; flappy_W(53, 535) <= 1; flappy_W(53, 536) <= 1; flappy_W(53, 537) <= 1; flappy_W(53, 538) <= 1; flappy_W(53, 539) <= 1; flappy_W(53, 540) <= 1; flappy_W(53, 541) <= 1; flappy_W(53, 542) <= 1; flappy_W(53, 543) <= 1; flappy_W(53, 544) <= 1; flappy_W(53, 545) <= 1; flappy_W(53, 546) <= 0; flappy_W(53, 547) <= 0; flappy_W(53, 548) <= 0; flappy_W(53, 549) <= 0; flappy_W(53, 550) <= 0; flappy_W(53, 551) <= 0; flappy_W(53, 552) <= 0; flappy_W(53, 553) <= 0; flappy_W(53, 554) <= 0; flappy_W(53, 555) <= 0; flappy_W(53, 556) <= 0; flappy_W(53, 557) <= 0; flappy_W(53, 558) <= 0; flappy_W(53, 559) <= 0; flappy_W(53, 560) <= 0; flappy_W(53, 561) <= 0; flappy_W(53, 562) <= 0; flappy_W(53, 563) <= 0; flappy_W(53, 564) <= 1; flappy_W(53, 565) <= 1; flappy_W(53, 566) <= 1; flappy_W(53, 567) <= 1; flappy_W(53, 568) <= 1; flappy_W(53, 569) <= 1; flappy_W(53, 570) <= 1; flappy_W(53, 571) <= 1; flappy_W(53, 572) <= 1; flappy_W(53, 573) <= 1; flappy_W(53, 574) <= 1; flappy_W(53, 575) <= 1; flappy_W(53, 576) <= 0; flappy_W(53, 577) <= 0; flappy_W(53, 578) <= 0; flappy_W(53, 579) <= 0; flappy_W(53, 580) <= 0; flappy_W(53, 581) <= 0; flappy_W(53, 582) <= 1; flappy_W(53, 583) <= 1; flappy_W(53, 584) <= 1; flappy_W(53, 585) <= 1; flappy_W(53, 586) <= 1; flappy_W(53, 587) <= 1; flappy_W(53, 588) <= 1; flappy_W(53, 589) <= 1; flappy_W(53, 590) <= 1; flappy_W(53, 591) <= 1; flappy_W(53, 592) <= 1; flappy_W(53, 593) <= 1; 
flappy_W(54, 0) <= 1; flappy_W(54, 1) <= 1; flappy_W(54, 2) <= 1; flappy_W(54, 3) <= 1; flappy_W(54, 4) <= 1; flappy_W(54, 5) <= 1; flappy_W(54, 6) <= 1; flappy_W(54, 7) <= 1; flappy_W(54, 8) <= 1; flappy_W(54, 9) <= 1; flappy_W(54, 10) <= 1; flappy_W(54, 11) <= 1; flappy_W(54, 12) <= 1; flappy_W(54, 13) <= 1; flappy_W(54, 14) <= 1; flappy_W(54, 15) <= 1; flappy_W(54, 16) <= 1; flappy_W(54, 17) <= 1; flappy_W(54, 18) <= 1; flappy_W(54, 19) <= 1; flappy_W(54, 20) <= 1; flappy_W(54, 21) <= 1; flappy_W(54, 22) <= 1; flappy_W(54, 23) <= 1; flappy_W(54, 24) <= 0; flappy_W(54, 25) <= 0; flappy_W(54, 26) <= 0; flappy_W(54, 27) <= 0; flappy_W(54, 28) <= 0; flappy_W(54, 29) <= 0; flappy_W(54, 30) <= 0; flappy_W(54, 31) <= 0; flappy_W(54, 32) <= 0; flappy_W(54, 33) <= 0; flappy_W(54, 34) <= 0; flappy_W(54, 35) <= 0; flappy_W(54, 36) <= 0; flappy_W(54, 37) <= 0; flappy_W(54, 38) <= 0; flappy_W(54, 39) <= 0; flappy_W(54, 40) <= 0; flappy_W(54, 41) <= 0; flappy_W(54, 42) <= 0; flappy_W(54, 43) <= 0; flappy_W(54, 44) <= 0; flappy_W(54, 45) <= 0; flappy_W(54, 46) <= 0; flappy_W(54, 47) <= 0; flappy_W(54, 48) <= 0; flappy_W(54, 49) <= 0; flappy_W(54, 50) <= 0; flappy_W(54, 51) <= 0; flappy_W(54, 52) <= 0; flappy_W(54, 53) <= 0; flappy_W(54, 54) <= 1; flappy_W(54, 55) <= 1; flappy_W(54, 56) <= 1; flappy_W(54, 57) <= 1; flappy_W(54, 58) <= 1; flappy_W(54, 59) <= 1; flappy_W(54, 60) <= 1; flappy_W(54, 61) <= 1; flappy_W(54, 62) <= 1; flappy_W(54, 63) <= 1; flappy_W(54, 64) <= 1; flappy_W(54, 65) <= 1; flappy_W(54, 66) <= 1; flappy_W(54, 67) <= 1; flappy_W(54, 68) <= 1; flappy_W(54, 69) <= 1; flappy_W(54, 70) <= 1; flappy_W(54, 71) <= 1; flappy_W(54, 72) <= 1; flappy_W(54, 73) <= 1; flappy_W(54, 74) <= 1; flappy_W(54, 75) <= 1; flappy_W(54, 76) <= 1; flappy_W(54, 77) <= 1; flappy_W(54, 78) <= 1; flappy_W(54, 79) <= 1; flappy_W(54, 80) <= 1; flappy_W(54, 81) <= 1; flappy_W(54, 82) <= 1; flappy_W(54, 83) <= 1; flappy_W(54, 84) <= 1; flappy_W(54, 85) <= 1; flappy_W(54, 86) <= 1; flappy_W(54, 87) <= 1; flappy_W(54, 88) <= 1; flappy_W(54, 89) <= 1; flappy_W(54, 90) <= 1; flappy_W(54, 91) <= 1; flappy_W(54, 92) <= 1; flappy_W(54, 93) <= 1; flappy_W(54, 94) <= 1; flappy_W(54, 95) <= 1; flappy_W(54, 96) <= 0; flappy_W(54, 97) <= 0; flappy_W(54, 98) <= 0; flappy_W(54, 99) <= 0; flappy_W(54, 100) <= 0; flappy_W(54, 101) <= 0; flappy_W(54, 102) <= 0; flappy_W(54, 103) <= 0; flappy_W(54, 104) <= 0; flappy_W(54, 105) <= 0; flappy_W(54, 106) <= 0; flappy_W(54, 107) <= 0; flappy_W(54, 108) <= 1; flappy_W(54, 109) <= 1; flappy_W(54, 110) <= 1; flappy_W(54, 111) <= 1; flappy_W(54, 112) <= 1; flappy_W(54, 113) <= 1; flappy_W(54, 114) <= 1; flappy_W(54, 115) <= 1; flappy_W(54, 116) <= 1; flappy_W(54, 117) <= 1; flappy_W(54, 118) <= 1; flappy_W(54, 119) <= 1; flappy_W(54, 120) <= 0; flappy_W(54, 121) <= 0; flappy_W(54, 122) <= 0; flappy_W(54, 123) <= 0; flappy_W(54, 124) <= 0; flappy_W(54, 125) <= 0; flappy_W(54, 126) <= 0; flappy_W(54, 127) <= 0; flappy_W(54, 128) <= 0; flappy_W(54, 129) <= 0; flappy_W(54, 130) <= 0; flappy_W(54, 131) <= 0; flappy_W(54, 132) <= 0; flappy_W(54, 133) <= 0; flappy_W(54, 134) <= 0; flappy_W(54, 135) <= 0; flappy_W(54, 136) <= 0; flappy_W(54, 137) <= 0; flappy_W(54, 138) <= 1; flappy_W(54, 139) <= 1; flappy_W(54, 140) <= 1; flappy_W(54, 141) <= 1; flappy_W(54, 142) <= 1; flappy_W(54, 143) <= 1; flappy_W(54, 144) <= 1; flappy_W(54, 145) <= 1; flappy_W(54, 146) <= 1; flappy_W(54, 147) <= 1; flappy_W(54, 148) <= 1; flappy_W(54, 149) <= 1; flappy_W(54, 150) <= 0; flappy_W(54, 151) <= 0; flappy_W(54, 152) <= 0; flappy_W(54, 153) <= 0; flappy_W(54, 154) <= 0; flappy_W(54, 155) <= 0; flappy_W(54, 156) <= 0; flappy_W(54, 157) <= 0; flappy_W(54, 158) <= 0; flappy_W(54, 159) <= 0; flappy_W(54, 160) <= 0; flappy_W(54, 161) <= 0; flappy_W(54, 162) <= 1; flappy_W(54, 163) <= 1; flappy_W(54, 164) <= 1; flappy_W(54, 165) <= 1; flappy_W(54, 166) <= 1; flappy_W(54, 167) <= 1; flappy_W(54, 168) <= 1; flappy_W(54, 169) <= 1; flappy_W(54, 170) <= 1; flappy_W(54, 171) <= 1; flappy_W(54, 172) <= 1; flappy_W(54, 173) <= 1; flappy_W(54, 174) <= 1; flappy_W(54, 175) <= 1; flappy_W(54, 176) <= 1; flappy_W(54, 177) <= 1; flappy_W(54, 178) <= 1; flappy_W(54, 179) <= 1; flappy_W(54, 180) <= 1; flappy_W(54, 181) <= 1; flappy_W(54, 182) <= 1; flappy_W(54, 183) <= 1; flappy_W(54, 184) <= 1; flappy_W(54, 185) <= 1; flappy_W(54, 186) <= 0; flappy_W(54, 187) <= 0; flappy_W(54, 188) <= 0; flappy_W(54, 189) <= 0; flappy_W(54, 190) <= 0; flappy_W(54, 191) <= 0; flappy_W(54, 192) <= 0; flappy_W(54, 193) <= 0; flappy_W(54, 194) <= 0; flappy_W(54, 195) <= 0; flappy_W(54, 196) <= 0; flappy_W(54, 197) <= 0; flappy_W(54, 198) <= 0; flappy_W(54, 199) <= 0; flappy_W(54, 200) <= 0; flappy_W(54, 201) <= 0; flappy_W(54, 202) <= 0; flappy_W(54, 203) <= 0; flappy_W(54, 204) <= 0; flappy_W(54, 205) <= 0; flappy_W(54, 206) <= 0; flappy_W(54, 207) <= 0; flappy_W(54, 208) <= 0; flappy_W(54, 209) <= 0; flappy_W(54, 210) <= 0; flappy_W(54, 211) <= 0; flappy_W(54, 212) <= 0; flappy_W(54, 213) <= 0; flappy_W(54, 214) <= 0; flappy_W(54, 215) <= 0; flappy_W(54, 216) <= 1; flappy_W(54, 217) <= 1; flappy_W(54, 218) <= 1; flappy_W(54, 219) <= 1; flappy_W(54, 220) <= 1; flappy_W(54, 221) <= 1; flappy_W(54, 222) <= 1; flappy_W(54, 223) <= 1; flappy_W(54, 224) <= 1; flappy_W(54, 225) <= 1; flappy_W(54, 226) <= 1; flappy_W(54, 227) <= 1; flappy_W(54, 228) <= 1; flappy_W(54, 229) <= 1; flappy_W(54, 230) <= 1; flappy_W(54, 231) <= 1; flappy_W(54, 232) <= 1; flappy_W(54, 233) <= 1; flappy_W(54, 234) <= 1; flappy_W(54, 235) <= 1; flappy_W(54, 236) <= 1; flappy_W(54, 237) <= 1; flappy_W(54, 238) <= 1; flappy_W(54, 239) <= 1; flappy_W(54, 240) <= 0; flappy_W(54, 241) <= 0; flappy_W(54, 242) <= 0; flappy_W(54, 243) <= 0; flappy_W(54, 244) <= 0; flappy_W(54, 245) <= 0; flappy_W(54, 246) <= 0; flappy_W(54, 247) <= 0; flappy_W(54, 248) <= 0; flappy_W(54, 249) <= 0; flappy_W(54, 250) <= 0; flappy_W(54, 251) <= 0; flappy_W(54, 252) <= 0; flappy_W(54, 253) <= 0; flappy_W(54, 254) <= 0; flappy_W(54, 255) <= 0; flappy_W(54, 256) <= 0; flappy_W(54, 257) <= 0; flappy_W(54, 258) <= 0; flappy_W(54, 259) <= 0; flappy_W(54, 260) <= 0; flappy_W(54, 261) <= 0; flappy_W(54, 262) <= 0; flappy_W(54, 263) <= 0; flappy_W(54, 264) <= 0; flappy_W(54, 265) <= 0; flappy_W(54, 266) <= 0; flappy_W(54, 267) <= 0; flappy_W(54, 268) <= 0; flappy_W(54, 269) <= 0; flappy_W(54, 270) <= 0; flappy_W(54, 271) <= 0; flappy_W(54, 272) <= 0; flappy_W(54, 273) <= 0; flappy_W(54, 274) <= 0; flappy_W(54, 275) <= 0; flappy_W(54, 276) <= 0; flappy_W(54, 277) <= 0; flappy_W(54, 278) <= 0; flappy_W(54, 279) <= 0; flappy_W(54, 280) <= 0; flappy_W(54, 281) <= 0; flappy_W(54, 282) <= 1; flappy_W(54, 283) <= 1; flappy_W(54, 284) <= 1; flappy_W(54, 285) <= 1; flappy_W(54, 286) <= 1; flappy_W(54, 287) <= 1; flappy_W(54, 288) <= 1; flappy_W(54, 289) <= 1; flappy_W(54, 290) <= 1; flappy_W(54, 291) <= 1; flappy_W(54, 292) <= 1; flappy_W(54, 293) <= 1; flappy_W(54, 294) <= 1; flappy_W(54, 295) <= 1; flappy_W(54, 296) <= 1; flappy_W(54, 297) <= 1; flappy_W(54, 298) <= 1; flappy_W(54, 299) <= 1; flappy_W(54, 300) <= 1; flappy_W(54, 301) <= 1; flappy_W(54, 302) <= 1; flappy_W(54, 303) <= 1; flappy_W(54, 304) <= 1; flappy_W(54, 305) <= 1; flappy_W(54, 306) <= 0; flappy_W(54, 307) <= 0; flappy_W(54, 308) <= 0; flappy_W(54, 309) <= 0; flappy_W(54, 310) <= 0; flappy_W(54, 311) <= 0; flappy_W(54, 312) <= 0; flappy_W(54, 313) <= 0; flappy_W(54, 314) <= 0; flappy_W(54, 315) <= 0; flappy_W(54, 316) <= 0; flappy_W(54, 317) <= 0; flappy_W(54, 318) <= 0; flappy_W(54, 319) <= 0; flappy_W(54, 320) <= 0; flappy_W(54, 321) <= 0; flappy_W(54, 322) <= 0; flappy_W(54, 323) <= 0; flappy_W(54, 324) <= 0; flappy_W(54, 325) <= 0; flappy_W(54, 326) <= 0; flappy_W(54, 327) <= 0; flappy_W(54, 328) <= 0; flappy_W(54, 329) <= 0; flappy_W(54, 330) <= 0; flappy_W(54, 331) <= 0; flappy_W(54, 332) <= 0; flappy_W(54, 333) <= 0; flappy_W(54, 334) <= 0; flappy_W(54, 335) <= 0; flappy_W(54, 336) <= 0; flappy_W(54, 337) <= 0; flappy_W(54, 338) <= 0; flappy_W(54, 339) <= 0; flappy_W(54, 340) <= 0; flappy_W(54, 341) <= 0; flappy_W(54, 342) <= 0; flappy_W(54, 343) <= 0; flappy_W(54, 344) <= 0; flappy_W(54, 345) <= 0; flappy_W(54, 346) <= 0; flappy_W(54, 347) <= 0; flappy_W(54, 348) <= 0; flappy_W(54, 349) <= 0; flappy_W(54, 350) <= 0; flappy_W(54, 351) <= 0; flappy_W(54, 352) <= 0; flappy_W(54, 353) <= 0; flappy_W(54, 354) <= 0; flappy_W(54, 355) <= 0; flappy_W(54, 356) <= 0; flappy_W(54, 357) <= 0; flappy_W(54, 358) <= 0; flappy_W(54, 359) <= 0; flappy_W(54, 360) <= 0; flappy_W(54, 361) <= 0; flappy_W(54, 362) <= 0; flappy_W(54, 363) <= 0; flappy_W(54, 364) <= 0; flappy_W(54, 365) <= 0; flappy_W(54, 366) <= 0; flappy_W(54, 367) <= 0; flappy_W(54, 368) <= 0; flappy_W(54, 369) <= 0; flappy_W(54, 370) <= 0; flappy_W(54, 371) <= 0; flappy_W(54, 372) <= 0; flappy_W(54, 373) <= 0; flappy_W(54, 374) <= 0; flappy_W(54, 375) <= 0; flappy_W(54, 376) <= 0; flappy_W(54, 377) <= 0; flappy_W(54, 378) <= 0; flappy_W(54, 379) <= 0; flappy_W(54, 380) <= 0; flappy_W(54, 381) <= 0; flappy_W(54, 382) <= 0; flappy_W(54, 383) <= 0; flappy_W(54, 384) <= 0; flappy_W(54, 385) <= 0; flappy_W(54, 386) <= 0; flappy_W(54, 387) <= 0; flappy_W(54, 388) <= 0; flappy_W(54, 389) <= 0; flappy_W(54, 390) <= 0; flappy_W(54, 391) <= 0; flappy_W(54, 392) <= 0; flappy_W(54, 393) <= 0; flappy_W(54, 394) <= 0; flappy_W(54, 395) <= 0; flappy_W(54, 396) <= 1; flappy_W(54, 397) <= 1; flappy_W(54, 398) <= 1; flappy_W(54, 399) <= 1; flappy_W(54, 400) <= 1; flappy_W(54, 401) <= 1; flappy_W(54, 402) <= 1; flappy_W(54, 403) <= 1; flappy_W(54, 404) <= 1; flappy_W(54, 405) <= 1; flappy_W(54, 406) <= 1; flappy_W(54, 407) <= 1; flappy_W(54, 408) <= 1; flappy_W(54, 409) <= 1; flappy_W(54, 410) <= 1; flappy_W(54, 411) <= 1; flappy_W(54, 412) <= 1; flappy_W(54, 413) <= 1; flappy_W(54, 414) <= 1; flappy_W(54, 415) <= 1; flappy_W(54, 416) <= 1; flappy_W(54, 417) <= 1; flappy_W(54, 418) <= 1; flappy_W(54, 419) <= 1; flappy_W(54, 420) <= 1; flappy_W(54, 421) <= 1; flappy_W(54, 422) <= 1; flappy_W(54, 423) <= 1; flappy_W(54, 424) <= 1; flappy_W(54, 425) <= 1; flappy_W(54, 426) <= 1; flappy_W(54, 427) <= 1; flappy_W(54, 428) <= 1; flappy_W(54, 429) <= 1; flappy_W(54, 430) <= 1; flappy_W(54, 431) <= 1; flappy_W(54, 432) <= 0; flappy_W(54, 433) <= 0; flappy_W(54, 434) <= 0; flappy_W(54, 435) <= 0; flappy_W(54, 436) <= 0; flappy_W(54, 437) <= 0; flappy_W(54, 438) <= 0; flappy_W(54, 439) <= 0; flappy_W(54, 440) <= 0; flappy_W(54, 441) <= 0; flappy_W(54, 442) <= 0; flappy_W(54, 443) <= 0; flappy_W(54, 444) <= 0; flappy_W(54, 445) <= 0; flappy_W(54, 446) <= 0; flappy_W(54, 447) <= 0; flappy_W(54, 448) <= 0; flappy_W(54, 449) <= 0; flappy_W(54, 450) <= 0; flappy_W(54, 451) <= 0; flappy_W(54, 452) <= 0; flappy_W(54, 453) <= 0; flappy_W(54, 454) <= 0; flappy_W(54, 455) <= 0; flappy_W(54, 456) <= 0; flappy_W(54, 457) <= 0; flappy_W(54, 458) <= 0; flappy_W(54, 459) <= 0; flappy_W(54, 460) <= 0; flappy_W(54, 461) <= 0; flappy_W(54, 462) <= 1; flappy_W(54, 463) <= 1; flappy_W(54, 464) <= 1; flappy_W(54, 465) <= 1; flappy_W(54, 466) <= 1; flappy_W(54, 467) <= 1; flappy_W(54, 468) <= 1; flappy_W(54, 469) <= 1; flappy_W(54, 470) <= 1; flappy_W(54, 471) <= 1; flappy_W(54, 472) <= 1; flappy_W(54, 473) <= 1; flappy_W(54, 474) <= 1; flappy_W(54, 475) <= 1; flappy_W(54, 476) <= 1; flappy_W(54, 477) <= 1; flappy_W(54, 478) <= 1; flappy_W(54, 479) <= 1; flappy_W(54, 480) <= 1; flappy_W(54, 481) <= 1; flappy_W(54, 482) <= 1; flappy_W(54, 483) <= 1; flappy_W(54, 484) <= 1; flappy_W(54, 485) <= 1; flappy_W(54, 486) <= 0; flappy_W(54, 487) <= 0; flappy_W(54, 488) <= 0; flappy_W(54, 489) <= 0; flappy_W(54, 490) <= 0; flappy_W(54, 491) <= 0; flappy_W(54, 492) <= 0; flappy_W(54, 493) <= 0; flappy_W(54, 494) <= 0; flappy_W(54, 495) <= 0; flappy_W(54, 496) <= 0; flappy_W(54, 497) <= 0; flappy_W(54, 498) <= 0; flappy_W(54, 499) <= 0; flappy_W(54, 500) <= 0; flappy_W(54, 501) <= 0; flappy_W(54, 502) <= 0; flappy_W(54, 503) <= 0; flappy_W(54, 504) <= 1; flappy_W(54, 505) <= 1; flappy_W(54, 506) <= 1; flappy_W(54, 507) <= 1; flappy_W(54, 508) <= 1; flappy_W(54, 509) <= 1; flappy_W(54, 510) <= 1; flappy_W(54, 511) <= 1; flappy_W(54, 512) <= 1; flappy_W(54, 513) <= 1; flappy_W(54, 514) <= 1; flappy_W(54, 515) <= 1; flappy_W(54, 516) <= 1; flappy_W(54, 517) <= 1; flappy_W(54, 518) <= 1; flappy_W(54, 519) <= 1; flappy_W(54, 520) <= 1; flappy_W(54, 521) <= 1; flappy_W(54, 522) <= 0; flappy_W(54, 523) <= 0; flappy_W(54, 524) <= 0; flappy_W(54, 525) <= 0; flappy_W(54, 526) <= 0; flappy_W(54, 527) <= 0; flappy_W(54, 528) <= 0; flappy_W(54, 529) <= 0; flappy_W(54, 530) <= 0; flappy_W(54, 531) <= 0; flappy_W(54, 532) <= 0; flappy_W(54, 533) <= 0; flappy_W(54, 534) <= 1; flappy_W(54, 535) <= 1; flappy_W(54, 536) <= 1; flappy_W(54, 537) <= 1; flappy_W(54, 538) <= 1; flappy_W(54, 539) <= 1; flappy_W(54, 540) <= 1; flappy_W(54, 541) <= 1; flappy_W(54, 542) <= 1; flappy_W(54, 543) <= 1; flappy_W(54, 544) <= 1; flappy_W(54, 545) <= 1; flappy_W(54, 546) <= 0; flappy_W(54, 547) <= 0; flappy_W(54, 548) <= 0; flappy_W(54, 549) <= 0; flappy_W(54, 550) <= 0; flappy_W(54, 551) <= 0; flappy_W(54, 552) <= 0; flappy_W(54, 553) <= 0; flappy_W(54, 554) <= 0; flappy_W(54, 555) <= 0; flappy_W(54, 556) <= 0; flappy_W(54, 557) <= 0; flappy_W(54, 558) <= 1; flappy_W(54, 559) <= 1; flappy_W(54, 560) <= 1; flappy_W(54, 561) <= 1; flappy_W(54, 562) <= 1; flappy_W(54, 563) <= 1; flappy_W(54, 564) <= 1; flappy_W(54, 565) <= 1; flappy_W(54, 566) <= 1; flappy_W(54, 567) <= 1; flappy_W(54, 568) <= 1; flappy_W(54, 569) <= 1; flappy_W(54, 570) <= 1; flappy_W(54, 571) <= 1; flappy_W(54, 572) <= 1; flappy_W(54, 573) <= 1; flappy_W(54, 574) <= 1; flappy_W(54, 575) <= 1; flappy_W(54, 576) <= 1; flappy_W(54, 577) <= 1; flappy_W(54, 578) <= 1; flappy_W(54, 579) <= 1; flappy_W(54, 580) <= 1; flappy_W(54, 581) <= 1; flappy_W(54, 582) <= 1; flappy_W(54, 583) <= 1; flappy_W(54, 584) <= 1; flappy_W(54, 585) <= 1; flappy_W(54, 586) <= 1; flappy_W(54, 587) <= 1; flappy_W(54, 588) <= 0; flappy_W(54, 589) <= 0; flappy_W(54, 590) <= 0; flappy_W(54, 591) <= 0; flappy_W(54, 592) <= 0; flappy_W(54, 593) <= 0; 
flappy_W(55, 0) <= 1; flappy_W(55, 1) <= 1; flappy_W(55, 2) <= 1; flappy_W(55, 3) <= 1; flappy_W(55, 4) <= 1; flappy_W(55, 5) <= 1; flappy_W(55, 6) <= 1; flappy_W(55, 7) <= 1; flappy_W(55, 8) <= 1; flappy_W(55, 9) <= 1; flappy_W(55, 10) <= 1; flappy_W(55, 11) <= 1; flappy_W(55, 12) <= 1; flappy_W(55, 13) <= 1; flappy_W(55, 14) <= 1; flappy_W(55, 15) <= 1; flappy_W(55, 16) <= 1; flappy_W(55, 17) <= 1; flappy_W(55, 18) <= 1; flappy_W(55, 19) <= 1; flappy_W(55, 20) <= 1; flappy_W(55, 21) <= 1; flappy_W(55, 22) <= 1; flappy_W(55, 23) <= 1; flappy_W(55, 24) <= 0; flappy_W(55, 25) <= 0; flappy_W(55, 26) <= 0; flappy_W(55, 27) <= 0; flappy_W(55, 28) <= 0; flappy_W(55, 29) <= 0; flappy_W(55, 30) <= 0; flappy_W(55, 31) <= 0; flappy_W(55, 32) <= 0; flappy_W(55, 33) <= 0; flappy_W(55, 34) <= 0; flappy_W(55, 35) <= 0; flappy_W(55, 36) <= 0; flappy_W(55, 37) <= 0; flappy_W(55, 38) <= 0; flappy_W(55, 39) <= 0; flappy_W(55, 40) <= 0; flappy_W(55, 41) <= 0; flappy_W(55, 42) <= 0; flappy_W(55, 43) <= 0; flappy_W(55, 44) <= 0; flappy_W(55, 45) <= 0; flappy_W(55, 46) <= 0; flappy_W(55, 47) <= 0; flappy_W(55, 48) <= 0; flappy_W(55, 49) <= 0; flappy_W(55, 50) <= 0; flappy_W(55, 51) <= 0; flappy_W(55, 52) <= 0; flappy_W(55, 53) <= 0; flappy_W(55, 54) <= 1; flappy_W(55, 55) <= 1; flappy_W(55, 56) <= 1; flappy_W(55, 57) <= 1; flappy_W(55, 58) <= 1; flappy_W(55, 59) <= 1; flappy_W(55, 60) <= 1; flappy_W(55, 61) <= 1; flappy_W(55, 62) <= 1; flappy_W(55, 63) <= 1; flappy_W(55, 64) <= 1; flappy_W(55, 65) <= 1; flappy_W(55, 66) <= 1; flappy_W(55, 67) <= 1; flappy_W(55, 68) <= 1; flappy_W(55, 69) <= 1; flappy_W(55, 70) <= 1; flappy_W(55, 71) <= 1; flappy_W(55, 72) <= 1; flappy_W(55, 73) <= 1; flappy_W(55, 74) <= 1; flappy_W(55, 75) <= 1; flappy_W(55, 76) <= 1; flappy_W(55, 77) <= 1; flappy_W(55, 78) <= 1; flappy_W(55, 79) <= 1; flappy_W(55, 80) <= 1; flappy_W(55, 81) <= 1; flappy_W(55, 82) <= 1; flappy_W(55, 83) <= 1; flappy_W(55, 84) <= 1; flappy_W(55, 85) <= 1; flappy_W(55, 86) <= 1; flappy_W(55, 87) <= 1; flappy_W(55, 88) <= 1; flappy_W(55, 89) <= 1; flappy_W(55, 90) <= 1; flappy_W(55, 91) <= 1; flappy_W(55, 92) <= 1; flappy_W(55, 93) <= 1; flappy_W(55, 94) <= 1; flappy_W(55, 95) <= 1; flappy_W(55, 96) <= 0; flappy_W(55, 97) <= 0; flappy_W(55, 98) <= 0; flappy_W(55, 99) <= 0; flappy_W(55, 100) <= 0; flappy_W(55, 101) <= 0; flappy_W(55, 102) <= 0; flappy_W(55, 103) <= 0; flappy_W(55, 104) <= 0; flappy_W(55, 105) <= 0; flappy_W(55, 106) <= 0; flappy_W(55, 107) <= 0; flappy_W(55, 108) <= 1; flappy_W(55, 109) <= 1; flappy_W(55, 110) <= 1; flappy_W(55, 111) <= 1; flappy_W(55, 112) <= 1; flappy_W(55, 113) <= 1; flappy_W(55, 114) <= 1; flappy_W(55, 115) <= 1; flappy_W(55, 116) <= 1; flappy_W(55, 117) <= 1; flappy_W(55, 118) <= 1; flappy_W(55, 119) <= 1; flappy_W(55, 120) <= 0; flappy_W(55, 121) <= 0; flappy_W(55, 122) <= 0; flappy_W(55, 123) <= 0; flappy_W(55, 124) <= 0; flappy_W(55, 125) <= 0; flappy_W(55, 126) <= 0; flappy_W(55, 127) <= 0; flappy_W(55, 128) <= 0; flappy_W(55, 129) <= 0; flappy_W(55, 130) <= 0; flappy_W(55, 131) <= 0; flappy_W(55, 132) <= 0; flappy_W(55, 133) <= 0; flappy_W(55, 134) <= 0; flappy_W(55, 135) <= 0; flappy_W(55, 136) <= 0; flappy_W(55, 137) <= 0; flappy_W(55, 138) <= 1; flappy_W(55, 139) <= 1; flappy_W(55, 140) <= 1; flappy_W(55, 141) <= 1; flappy_W(55, 142) <= 1; flappy_W(55, 143) <= 1; flappy_W(55, 144) <= 1; flappy_W(55, 145) <= 1; flappy_W(55, 146) <= 1; flappy_W(55, 147) <= 1; flappy_W(55, 148) <= 1; flappy_W(55, 149) <= 1; flappy_W(55, 150) <= 0; flappy_W(55, 151) <= 0; flappy_W(55, 152) <= 0; flappy_W(55, 153) <= 0; flappy_W(55, 154) <= 0; flappy_W(55, 155) <= 0; flappy_W(55, 156) <= 0; flappy_W(55, 157) <= 0; flappy_W(55, 158) <= 0; flappy_W(55, 159) <= 0; flappy_W(55, 160) <= 0; flappy_W(55, 161) <= 0; flappy_W(55, 162) <= 1; flappy_W(55, 163) <= 1; flappy_W(55, 164) <= 1; flappy_W(55, 165) <= 1; flappy_W(55, 166) <= 1; flappy_W(55, 167) <= 1; flappy_W(55, 168) <= 1; flappy_W(55, 169) <= 1; flappy_W(55, 170) <= 1; flappy_W(55, 171) <= 1; flappy_W(55, 172) <= 1; flappy_W(55, 173) <= 1; flappy_W(55, 174) <= 1; flappy_W(55, 175) <= 1; flappy_W(55, 176) <= 1; flappy_W(55, 177) <= 1; flappy_W(55, 178) <= 1; flappy_W(55, 179) <= 1; flappy_W(55, 180) <= 1; flappy_W(55, 181) <= 1; flappy_W(55, 182) <= 1; flappy_W(55, 183) <= 1; flappy_W(55, 184) <= 1; flappy_W(55, 185) <= 1; flappy_W(55, 186) <= 0; flappy_W(55, 187) <= 0; flappy_W(55, 188) <= 0; flappy_W(55, 189) <= 0; flappy_W(55, 190) <= 0; flappy_W(55, 191) <= 0; flappy_W(55, 192) <= 0; flappy_W(55, 193) <= 0; flappy_W(55, 194) <= 0; flappy_W(55, 195) <= 0; flappy_W(55, 196) <= 0; flappy_W(55, 197) <= 0; flappy_W(55, 198) <= 0; flappy_W(55, 199) <= 0; flappy_W(55, 200) <= 0; flappy_W(55, 201) <= 0; flappy_W(55, 202) <= 0; flappy_W(55, 203) <= 0; flappy_W(55, 204) <= 0; flappy_W(55, 205) <= 0; flappy_W(55, 206) <= 0; flappy_W(55, 207) <= 0; flappy_W(55, 208) <= 0; flappy_W(55, 209) <= 0; flappy_W(55, 210) <= 0; flappy_W(55, 211) <= 0; flappy_W(55, 212) <= 0; flappy_W(55, 213) <= 0; flappy_W(55, 214) <= 0; flappy_W(55, 215) <= 0; flappy_W(55, 216) <= 1; flappy_W(55, 217) <= 1; flappy_W(55, 218) <= 1; flappy_W(55, 219) <= 1; flappy_W(55, 220) <= 1; flappy_W(55, 221) <= 1; flappy_W(55, 222) <= 1; flappy_W(55, 223) <= 1; flappy_W(55, 224) <= 1; flappy_W(55, 225) <= 1; flappy_W(55, 226) <= 1; flappy_W(55, 227) <= 1; flappy_W(55, 228) <= 1; flappy_W(55, 229) <= 1; flappy_W(55, 230) <= 1; flappy_W(55, 231) <= 1; flappy_W(55, 232) <= 1; flappy_W(55, 233) <= 1; flappy_W(55, 234) <= 1; flappy_W(55, 235) <= 1; flappy_W(55, 236) <= 1; flappy_W(55, 237) <= 1; flappy_W(55, 238) <= 1; flappy_W(55, 239) <= 1; flappy_W(55, 240) <= 0; flappy_W(55, 241) <= 0; flappy_W(55, 242) <= 0; flappy_W(55, 243) <= 0; flappy_W(55, 244) <= 0; flappy_W(55, 245) <= 0; flappy_W(55, 246) <= 0; flappy_W(55, 247) <= 0; flappy_W(55, 248) <= 0; flappy_W(55, 249) <= 0; flappy_W(55, 250) <= 0; flappy_W(55, 251) <= 0; flappy_W(55, 252) <= 0; flappy_W(55, 253) <= 0; flappy_W(55, 254) <= 0; flappy_W(55, 255) <= 0; flappy_W(55, 256) <= 0; flappy_W(55, 257) <= 0; flappy_W(55, 258) <= 0; flappy_W(55, 259) <= 0; flappy_W(55, 260) <= 0; flappy_W(55, 261) <= 0; flappy_W(55, 262) <= 0; flappy_W(55, 263) <= 0; flappy_W(55, 264) <= 0; flappy_W(55, 265) <= 0; flappy_W(55, 266) <= 0; flappy_W(55, 267) <= 0; flappy_W(55, 268) <= 0; flappy_W(55, 269) <= 0; flappy_W(55, 270) <= 0; flappy_W(55, 271) <= 0; flappy_W(55, 272) <= 0; flappy_W(55, 273) <= 0; flappy_W(55, 274) <= 0; flappy_W(55, 275) <= 0; flappy_W(55, 276) <= 0; flappy_W(55, 277) <= 0; flappy_W(55, 278) <= 0; flappy_W(55, 279) <= 0; flappy_W(55, 280) <= 0; flappy_W(55, 281) <= 0; flappy_W(55, 282) <= 1; flappy_W(55, 283) <= 1; flappy_W(55, 284) <= 1; flappy_W(55, 285) <= 1; flappy_W(55, 286) <= 1; flappy_W(55, 287) <= 1; flappy_W(55, 288) <= 1; flappy_W(55, 289) <= 1; flappy_W(55, 290) <= 1; flappy_W(55, 291) <= 1; flappy_W(55, 292) <= 1; flappy_W(55, 293) <= 1; flappy_W(55, 294) <= 1; flappy_W(55, 295) <= 1; flappy_W(55, 296) <= 1; flappy_W(55, 297) <= 1; flappy_W(55, 298) <= 1; flappy_W(55, 299) <= 1; flappy_W(55, 300) <= 1; flappy_W(55, 301) <= 1; flappy_W(55, 302) <= 1; flappy_W(55, 303) <= 1; flappy_W(55, 304) <= 1; flappy_W(55, 305) <= 1; flappy_W(55, 306) <= 0; flappy_W(55, 307) <= 0; flappy_W(55, 308) <= 0; flappy_W(55, 309) <= 0; flappy_W(55, 310) <= 0; flappy_W(55, 311) <= 0; flappy_W(55, 312) <= 0; flappy_W(55, 313) <= 0; flappy_W(55, 314) <= 0; flappy_W(55, 315) <= 0; flappy_W(55, 316) <= 0; flappy_W(55, 317) <= 0; flappy_W(55, 318) <= 0; flappy_W(55, 319) <= 0; flappy_W(55, 320) <= 0; flappy_W(55, 321) <= 0; flappy_W(55, 322) <= 0; flappy_W(55, 323) <= 0; flappy_W(55, 324) <= 0; flappy_W(55, 325) <= 0; flappy_W(55, 326) <= 0; flappy_W(55, 327) <= 0; flappy_W(55, 328) <= 0; flappy_W(55, 329) <= 0; flappy_W(55, 330) <= 0; flappy_W(55, 331) <= 0; flappy_W(55, 332) <= 0; flappy_W(55, 333) <= 0; flappy_W(55, 334) <= 0; flappy_W(55, 335) <= 0; flappy_W(55, 336) <= 0; flappy_W(55, 337) <= 0; flappy_W(55, 338) <= 0; flappy_W(55, 339) <= 0; flappy_W(55, 340) <= 0; flappy_W(55, 341) <= 0; flappy_W(55, 342) <= 0; flappy_W(55, 343) <= 0; flappy_W(55, 344) <= 0; flappy_W(55, 345) <= 0; flappy_W(55, 346) <= 0; flappy_W(55, 347) <= 0; flappy_W(55, 348) <= 0; flappy_W(55, 349) <= 0; flappy_W(55, 350) <= 0; flappy_W(55, 351) <= 0; flappy_W(55, 352) <= 0; flappy_W(55, 353) <= 0; flappy_W(55, 354) <= 0; flappy_W(55, 355) <= 0; flappy_W(55, 356) <= 0; flappy_W(55, 357) <= 0; flappy_W(55, 358) <= 0; flappy_W(55, 359) <= 0; flappy_W(55, 360) <= 0; flappy_W(55, 361) <= 0; flappy_W(55, 362) <= 0; flappy_W(55, 363) <= 0; flappy_W(55, 364) <= 0; flappy_W(55, 365) <= 0; flappy_W(55, 366) <= 0; flappy_W(55, 367) <= 0; flappy_W(55, 368) <= 0; flappy_W(55, 369) <= 0; flappy_W(55, 370) <= 0; flappy_W(55, 371) <= 0; flappy_W(55, 372) <= 0; flappy_W(55, 373) <= 0; flappy_W(55, 374) <= 0; flappy_W(55, 375) <= 0; flappy_W(55, 376) <= 0; flappy_W(55, 377) <= 0; flappy_W(55, 378) <= 0; flappy_W(55, 379) <= 0; flappy_W(55, 380) <= 0; flappy_W(55, 381) <= 0; flappy_W(55, 382) <= 0; flappy_W(55, 383) <= 0; flappy_W(55, 384) <= 0; flappy_W(55, 385) <= 0; flappy_W(55, 386) <= 0; flappy_W(55, 387) <= 0; flappy_W(55, 388) <= 0; flappy_W(55, 389) <= 0; flappy_W(55, 390) <= 0; flappy_W(55, 391) <= 0; flappy_W(55, 392) <= 0; flappy_W(55, 393) <= 0; flappy_W(55, 394) <= 0; flappy_W(55, 395) <= 0; flappy_W(55, 396) <= 1; flappy_W(55, 397) <= 1; flappy_W(55, 398) <= 1; flappy_W(55, 399) <= 1; flappy_W(55, 400) <= 1; flappy_W(55, 401) <= 1; flappy_W(55, 402) <= 1; flappy_W(55, 403) <= 1; flappy_W(55, 404) <= 1; flappy_W(55, 405) <= 1; flappy_W(55, 406) <= 1; flappy_W(55, 407) <= 1; flappy_W(55, 408) <= 1; flappy_W(55, 409) <= 1; flappy_W(55, 410) <= 1; flappy_W(55, 411) <= 1; flappy_W(55, 412) <= 1; flappy_W(55, 413) <= 1; flappy_W(55, 414) <= 1; flappy_W(55, 415) <= 1; flappy_W(55, 416) <= 1; flappy_W(55, 417) <= 1; flappy_W(55, 418) <= 1; flappy_W(55, 419) <= 1; flappy_W(55, 420) <= 1; flappy_W(55, 421) <= 1; flappy_W(55, 422) <= 1; flappy_W(55, 423) <= 1; flappy_W(55, 424) <= 1; flappy_W(55, 425) <= 1; flappy_W(55, 426) <= 1; flappy_W(55, 427) <= 1; flappy_W(55, 428) <= 1; flappy_W(55, 429) <= 1; flappy_W(55, 430) <= 1; flappy_W(55, 431) <= 1; flappy_W(55, 432) <= 0; flappy_W(55, 433) <= 0; flappy_W(55, 434) <= 0; flappy_W(55, 435) <= 0; flappy_W(55, 436) <= 0; flappy_W(55, 437) <= 0; flappy_W(55, 438) <= 0; flappy_W(55, 439) <= 0; flappy_W(55, 440) <= 0; flappy_W(55, 441) <= 0; flappy_W(55, 442) <= 0; flappy_W(55, 443) <= 0; flappy_W(55, 444) <= 0; flappy_W(55, 445) <= 0; flappy_W(55, 446) <= 0; flappy_W(55, 447) <= 0; flappy_W(55, 448) <= 0; flappy_W(55, 449) <= 0; flappy_W(55, 450) <= 0; flappy_W(55, 451) <= 0; flappy_W(55, 452) <= 0; flappy_W(55, 453) <= 0; flappy_W(55, 454) <= 0; flappy_W(55, 455) <= 0; flappy_W(55, 456) <= 0; flappy_W(55, 457) <= 0; flappy_W(55, 458) <= 0; flappy_W(55, 459) <= 0; flappy_W(55, 460) <= 0; flappy_W(55, 461) <= 0; flappy_W(55, 462) <= 1; flappy_W(55, 463) <= 1; flappy_W(55, 464) <= 1; flappy_W(55, 465) <= 1; flappy_W(55, 466) <= 1; flappy_W(55, 467) <= 1; flappy_W(55, 468) <= 1; flappy_W(55, 469) <= 1; flappy_W(55, 470) <= 1; flappy_W(55, 471) <= 1; flappy_W(55, 472) <= 1; flappy_W(55, 473) <= 1; flappy_W(55, 474) <= 1; flappy_W(55, 475) <= 1; flappy_W(55, 476) <= 1; flappy_W(55, 477) <= 1; flappy_W(55, 478) <= 1; flappy_W(55, 479) <= 1; flappy_W(55, 480) <= 1; flappy_W(55, 481) <= 1; flappy_W(55, 482) <= 1; flappy_W(55, 483) <= 1; flappy_W(55, 484) <= 1; flappy_W(55, 485) <= 1; flappy_W(55, 486) <= 0; flappy_W(55, 487) <= 0; flappy_W(55, 488) <= 0; flappy_W(55, 489) <= 0; flappy_W(55, 490) <= 0; flappy_W(55, 491) <= 0; flappy_W(55, 492) <= 0; flappy_W(55, 493) <= 0; flappy_W(55, 494) <= 0; flappy_W(55, 495) <= 0; flappy_W(55, 496) <= 0; flappy_W(55, 497) <= 0; flappy_W(55, 498) <= 0; flappy_W(55, 499) <= 0; flappy_W(55, 500) <= 0; flappy_W(55, 501) <= 0; flappy_W(55, 502) <= 0; flappy_W(55, 503) <= 0; flappy_W(55, 504) <= 1; flappy_W(55, 505) <= 1; flappy_W(55, 506) <= 1; flappy_W(55, 507) <= 1; flappy_W(55, 508) <= 1; flappy_W(55, 509) <= 1; flappy_W(55, 510) <= 1; flappy_W(55, 511) <= 1; flappy_W(55, 512) <= 1; flappy_W(55, 513) <= 1; flappy_W(55, 514) <= 1; flappy_W(55, 515) <= 1; flappy_W(55, 516) <= 1; flappy_W(55, 517) <= 1; flappy_W(55, 518) <= 1; flappy_W(55, 519) <= 1; flappy_W(55, 520) <= 1; flappy_W(55, 521) <= 1; flappy_W(55, 522) <= 0; flappy_W(55, 523) <= 0; flappy_W(55, 524) <= 0; flappy_W(55, 525) <= 0; flappy_W(55, 526) <= 0; flappy_W(55, 527) <= 0; flappy_W(55, 528) <= 0; flappy_W(55, 529) <= 0; flappy_W(55, 530) <= 0; flappy_W(55, 531) <= 0; flappy_W(55, 532) <= 0; flappy_W(55, 533) <= 0; flappy_W(55, 534) <= 1; flappy_W(55, 535) <= 1; flappy_W(55, 536) <= 1; flappy_W(55, 537) <= 1; flappy_W(55, 538) <= 1; flappy_W(55, 539) <= 1; flappy_W(55, 540) <= 1; flappy_W(55, 541) <= 1; flappy_W(55, 542) <= 1; flappy_W(55, 543) <= 1; flappy_W(55, 544) <= 1; flappy_W(55, 545) <= 1; flappy_W(55, 546) <= 0; flappy_W(55, 547) <= 0; flappy_W(55, 548) <= 0; flappy_W(55, 549) <= 0; flappy_W(55, 550) <= 0; flappy_W(55, 551) <= 0; flappy_W(55, 552) <= 0; flappy_W(55, 553) <= 0; flappy_W(55, 554) <= 0; flappy_W(55, 555) <= 0; flappy_W(55, 556) <= 0; flappy_W(55, 557) <= 0; flappy_W(55, 558) <= 1; flappy_W(55, 559) <= 1; flappy_W(55, 560) <= 1; flappy_W(55, 561) <= 1; flappy_W(55, 562) <= 1; flappy_W(55, 563) <= 1; flappy_W(55, 564) <= 1; flappy_W(55, 565) <= 1; flappy_W(55, 566) <= 1; flappy_W(55, 567) <= 1; flappy_W(55, 568) <= 1; flappy_W(55, 569) <= 1; flappy_W(55, 570) <= 1; flappy_W(55, 571) <= 1; flappy_W(55, 572) <= 1; flappy_W(55, 573) <= 1; flappy_W(55, 574) <= 1; flappy_W(55, 575) <= 1; flappy_W(55, 576) <= 1; flappy_W(55, 577) <= 1; flappy_W(55, 578) <= 1; flappy_W(55, 579) <= 1; flappy_W(55, 580) <= 1; flappy_W(55, 581) <= 1; flappy_W(55, 582) <= 1; flappy_W(55, 583) <= 1; flappy_W(55, 584) <= 1; flappy_W(55, 585) <= 1; flappy_W(55, 586) <= 1; flappy_W(55, 587) <= 1; flappy_W(55, 588) <= 0; flappy_W(55, 589) <= 0; flappy_W(55, 590) <= 0; flappy_W(55, 591) <= 0; flappy_W(55, 592) <= 0; flappy_W(55, 593) <= 0; 
flappy_W(56, 0) <= 1; flappy_W(56, 1) <= 1; flappy_W(56, 2) <= 1; flappy_W(56, 3) <= 1; flappy_W(56, 4) <= 1; flappy_W(56, 5) <= 1; flappy_W(56, 6) <= 1; flappy_W(56, 7) <= 1; flappy_W(56, 8) <= 1; flappy_W(56, 9) <= 1; flappy_W(56, 10) <= 1; flappy_W(56, 11) <= 1; flappy_W(56, 12) <= 1; flappy_W(56, 13) <= 1; flappy_W(56, 14) <= 1; flappy_W(56, 15) <= 1; flappy_W(56, 16) <= 1; flappy_W(56, 17) <= 1; flappy_W(56, 18) <= 1; flappy_W(56, 19) <= 1; flappy_W(56, 20) <= 1; flappy_W(56, 21) <= 1; flappy_W(56, 22) <= 1; flappy_W(56, 23) <= 1; flappy_W(56, 24) <= 0; flappy_W(56, 25) <= 0; flappy_W(56, 26) <= 0; flappy_W(56, 27) <= 0; flappy_W(56, 28) <= 0; flappy_W(56, 29) <= 0; flappy_W(56, 30) <= 0; flappy_W(56, 31) <= 0; flappy_W(56, 32) <= 0; flappy_W(56, 33) <= 0; flappy_W(56, 34) <= 0; flappy_W(56, 35) <= 0; flappy_W(56, 36) <= 0; flappy_W(56, 37) <= 0; flappy_W(56, 38) <= 0; flappy_W(56, 39) <= 0; flappy_W(56, 40) <= 0; flappy_W(56, 41) <= 0; flappy_W(56, 42) <= 0; flappy_W(56, 43) <= 0; flappy_W(56, 44) <= 0; flappy_W(56, 45) <= 0; flappy_W(56, 46) <= 0; flappy_W(56, 47) <= 0; flappy_W(56, 48) <= 0; flappy_W(56, 49) <= 0; flappy_W(56, 50) <= 0; flappy_W(56, 51) <= 0; flappy_W(56, 52) <= 0; flappy_W(56, 53) <= 0; flappy_W(56, 54) <= 1; flappy_W(56, 55) <= 1; flappy_W(56, 56) <= 1; flappy_W(56, 57) <= 1; flappy_W(56, 58) <= 1; flappy_W(56, 59) <= 1; flappy_W(56, 60) <= 1; flappy_W(56, 61) <= 1; flappy_W(56, 62) <= 1; flappy_W(56, 63) <= 1; flappy_W(56, 64) <= 1; flappy_W(56, 65) <= 1; flappy_W(56, 66) <= 1; flappy_W(56, 67) <= 1; flappy_W(56, 68) <= 1; flappy_W(56, 69) <= 1; flappy_W(56, 70) <= 1; flappy_W(56, 71) <= 1; flappy_W(56, 72) <= 1; flappy_W(56, 73) <= 1; flappy_W(56, 74) <= 1; flappy_W(56, 75) <= 1; flappy_W(56, 76) <= 1; flappy_W(56, 77) <= 1; flappy_W(56, 78) <= 1; flappy_W(56, 79) <= 1; flappy_W(56, 80) <= 1; flappy_W(56, 81) <= 1; flappy_W(56, 82) <= 1; flappy_W(56, 83) <= 1; flappy_W(56, 84) <= 1; flappy_W(56, 85) <= 1; flappy_W(56, 86) <= 1; flappy_W(56, 87) <= 1; flappy_W(56, 88) <= 1; flappy_W(56, 89) <= 1; flappy_W(56, 90) <= 1; flappy_W(56, 91) <= 1; flappy_W(56, 92) <= 1; flappy_W(56, 93) <= 1; flappy_W(56, 94) <= 1; flappy_W(56, 95) <= 1; flappy_W(56, 96) <= 0; flappy_W(56, 97) <= 0; flappy_W(56, 98) <= 0; flappy_W(56, 99) <= 0; flappy_W(56, 100) <= 0; flappy_W(56, 101) <= 0; flappy_W(56, 102) <= 0; flappy_W(56, 103) <= 0; flappy_W(56, 104) <= 0; flappy_W(56, 105) <= 0; flappy_W(56, 106) <= 0; flappy_W(56, 107) <= 0; flappy_W(56, 108) <= 1; flappy_W(56, 109) <= 1; flappy_W(56, 110) <= 1; flappy_W(56, 111) <= 1; flappy_W(56, 112) <= 1; flappy_W(56, 113) <= 1; flappy_W(56, 114) <= 1; flappy_W(56, 115) <= 1; flappy_W(56, 116) <= 1; flappy_W(56, 117) <= 1; flappy_W(56, 118) <= 1; flappy_W(56, 119) <= 1; flappy_W(56, 120) <= 0; flappy_W(56, 121) <= 0; flappy_W(56, 122) <= 0; flappy_W(56, 123) <= 0; flappy_W(56, 124) <= 0; flappy_W(56, 125) <= 0; flappy_W(56, 126) <= 0; flappy_W(56, 127) <= 0; flappy_W(56, 128) <= 0; flappy_W(56, 129) <= 0; flappy_W(56, 130) <= 0; flappy_W(56, 131) <= 0; flappy_W(56, 132) <= 0; flappy_W(56, 133) <= 0; flappy_W(56, 134) <= 0; flappy_W(56, 135) <= 0; flappy_W(56, 136) <= 0; flappy_W(56, 137) <= 0; flappy_W(56, 138) <= 1; flappy_W(56, 139) <= 1; flappy_W(56, 140) <= 1; flappy_W(56, 141) <= 1; flappy_W(56, 142) <= 1; flappy_W(56, 143) <= 1; flappy_W(56, 144) <= 1; flappy_W(56, 145) <= 1; flappy_W(56, 146) <= 1; flappy_W(56, 147) <= 1; flappy_W(56, 148) <= 1; flappy_W(56, 149) <= 1; flappy_W(56, 150) <= 0; flappy_W(56, 151) <= 0; flappy_W(56, 152) <= 0; flappy_W(56, 153) <= 0; flappy_W(56, 154) <= 0; flappy_W(56, 155) <= 0; flappy_W(56, 156) <= 0; flappy_W(56, 157) <= 0; flappy_W(56, 158) <= 0; flappy_W(56, 159) <= 0; flappy_W(56, 160) <= 0; flappy_W(56, 161) <= 0; flappy_W(56, 162) <= 1; flappy_W(56, 163) <= 1; flappy_W(56, 164) <= 1; flappy_W(56, 165) <= 1; flappy_W(56, 166) <= 1; flappy_W(56, 167) <= 1; flappy_W(56, 168) <= 1; flappy_W(56, 169) <= 1; flappy_W(56, 170) <= 1; flappy_W(56, 171) <= 1; flappy_W(56, 172) <= 1; flappy_W(56, 173) <= 1; flappy_W(56, 174) <= 1; flappy_W(56, 175) <= 1; flappy_W(56, 176) <= 1; flappy_W(56, 177) <= 1; flappy_W(56, 178) <= 1; flappy_W(56, 179) <= 1; flappy_W(56, 180) <= 1; flappy_W(56, 181) <= 1; flappy_W(56, 182) <= 1; flappy_W(56, 183) <= 1; flappy_W(56, 184) <= 1; flappy_W(56, 185) <= 1; flappy_W(56, 186) <= 0; flappy_W(56, 187) <= 0; flappy_W(56, 188) <= 0; flappy_W(56, 189) <= 0; flappy_W(56, 190) <= 0; flappy_W(56, 191) <= 0; flappy_W(56, 192) <= 0; flappy_W(56, 193) <= 0; flappy_W(56, 194) <= 0; flappy_W(56, 195) <= 0; flappy_W(56, 196) <= 0; flappy_W(56, 197) <= 0; flappy_W(56, 198) <= 0; flappy_W(56, 199) <= 0; flappy_W(56, 200) <= 0; flappy_W(56, 201) <= 0; flappy_W(56, 202) <= 0; flappy_W(56, 203) <= 0; flappy_W(56, 204) <= 0; flappy_W(56, 205) <= 0; flappy_W(56, 206) <= 0; flappy_W(56, 207) <= 0; flappy_W(56, 208) <= 0; flappy_W(56, 209) <= 0; flappy_W(56, 210) <= 0; flappy_W(56, 211) <= 0; flappy_W(56, 212) <= 0; flappy_W(56, 213) <= 0; flappy_W(56, 214) <= 0; flappy_W(56, 215) <= 0; flappy_W(56, 216) <= 1; flappy_W(56, 217) <= 1; flappy_W(56, 218) <= 1; flappy_W(56, 219) <= 1; flappy_W(56, 220) <= 1; flappy_W(56, 221) <= 1; flappy_W(56, 222) <= 1; flappy_W(56, 223) <= 1; flappy_W(56, 224) <= 1; flappy_W(56, 225) <= 1; flappy_W(56, 226) <= 1; flappy_W(56, 227) <= 1; flappy_W(56, 228) <= 1; flappy_W(56, 229) <= 1; flappy_W(56, 230) <= 1; flappy_W(56, 231) <= 1; flappy_W(56, 232) <= 1; flappy_W(56, 233) <= 1; flappy_W(56, 234) <= 1; flappy_W(56, 235) <= 1; flappy_W(56, 236) <= 1; flappy_W(56, 237) <= 1; flappy_W(56, 238) <= 1; flappy_W(56, 239) <= 1; flappy_W(56, 240) <= 0; flappy_W(56, 241) <= 0; flappy_W(56, 242) <= 0; flappy_W(56, 243) <= 0; flappy_W(56, 244) <= 0; flappy_W(56, 245) <= 0; flappy_W(56, 246) <= 0; flappy_W(56, 247) <= 0; flappy_W(56, 248) <= 0; flappy_W(56, 249) <= 0; flappy_W(56, 250) <= 0; flappy_W(56, 251) <= 0; flappy_W(56, 252) <= 0; flappy_W(56, 253) <= 0; flappy_W(56, 254) <= 0; flappy_W(56, 255) <= 0; flappy_W(56, 256) <= 0; flappy_W(56, 257) <= 0; flappy_W(56, 258) <= 0; flappy_W(56, 259) <= 0; flappy_W(56, 260) <= 0; flappy_W(56, 261) <= 0; flappy_W(56, 262) <= 0; flappy_W(56, 263) <= 0; flappy_W(56, 264) <= 0; flappy_W(56, 265) <= 0; flappy_W(56, 266) <= 0; flappy_W(56, 267) <= 0; flappy_W(56, 268) <= 0; flappy_W(56, 269) <= 0; flappy_W(56, 270) <= 0; flappy_W(56, 271) <= 0; flappy_W(56, 272) <= 0; flappy_W(56, 273) <= 0; flappy_W(56, 274) <= 0; flappy_W(56, 275) <= 0; flappy_W(56, 276) <= 0; flappy_W(56, 277) <= 0; flappy_W(56, 278) <= 0; flappy_W(56, 279) <= 0; flappy_W(56, 280) <= 0; flappy_W(56, 281) <= 0; flappy_W(56, 282) <= 1; flappy_W(56, 283) <= 1; flappy_W(56, 284) <= 1; flappy_W(56, 285) <= 1; flappy_W(56, 286) <= 1; flappy_W(56, 287) <= 1; flappy_W(56, 288) <= 1; flappy_W(56, 289) <= 1; flappy_W(56, 290) <= 1; flappy_W(56, 291) <= 1; flappy_W(56, 292) <= 1; flappy_W(56, 293) <= 1; flappy_W(56, 294) <= 1; flappy_W(56, 295) <= 1; flappy_W(56, 296) <= 1; flappy_W(56, 297) <= 1; flappy_W(56, 298) <= 1; flappy_W(56, 299) <= 1; flappy_W(56, 300) <= 1; flappy_W(56, 301) <= 1; flappy_W(56, 302) <= 1; flappy_W(56, 303) <= 1; flappy_W(56, 304) <= 1; flappy_W(56, 305) <= 1; flappy_W(56, 306) <= 0; flappy_W(56, 307) <= 0; flappy_W(56, 308) <= 0; flappy_W(56, 309) <= 0; flappy_W(56, 310) <= 0; flappy_W(56, 311) <= 0; flappy_W(56, 312) <= 0; flappy_W(56, 313) <= 0; flappy_W(56, 314) <= 0; flappy_W(56, 315) <= 0; flappy_W(56, 316) <= 0; flappy_W(56, 317) <= 0; flappy_W(56, 318) <= 0; flappy_W(56, 319) <= 0; flappy_W(56, 320) <= 0; flappy_W(56, 321) <= 0; flappy_W(56, 322) <= 0; flappy_W(56, 323) <= 0; flappy_W(56, 324) <= 0; flappy_W(56, 325) <= 0; flappy_W(56, 326) <= 0; flappy_W(56, 327) <= 0; flappy_W(56, 328) <= 0; flappy_W(56, 329) <= 0; flappy_W(56, 330) <= 0; flappy_W(56, 331) <= 0; flappy_W(56, 332) <= 0; flappy_W(56, 333) <= 0; flappy_W(56, 334) <= 0; flappy_W(56, 335) <= 0; flappy_W(56, 336) <= 0; flappy_W(56, 337) <= 0; flappy_W(56, 338) <= 0; flappy_W(56, 339) <= 0; flappy_W(56, 340) <= 0; flappy_W(56, 341) <= 0; flappy_W(56, 342) <= 0; flappy_W(56, 343) <= 0; flappy_W(56, 344) <= 0; flappy_W(56, 345) <= 0; flappy_W(56, 346) <= 0; flappy_W(56, 347) <= 0; flappy_W(56, 348) <= 0; flappy_W(56, 349) <= 0; flappy_W(56, 350) <= 0; flappy_W(56, 351) <= 0; flappy_W(56, 352) <= 0; flappy_W(56, 353) <= 0; flappy_W(56, 354) <= 0; flappy_W(56, 355) <= 0; flappy_W(56, 356) <= 0; flappy_W(56, 357) <= 0; flappy_W(56, 358) <= 0; flappy_W(56, 359) <= 0; flappy_W(56, 360) <= 0; flappy_W(56, 361) <= 0; flappy_W(56, 362) <= 0; flappy_W(56, 363) <= 0; flappy_W(56, 364) <= 0; flappy_W(56, 365) <= 0; flappy_W(56, 366) <= 0; flappy_W(56, 367) <= 0; flappy_W(56, 368) <= 0; flappy_W(56, 369) <= 0; flappy_W(56, 370) <= 0; flappy_W(56, 371) <= 0; flappy_W(56, 372) <= 0; flappy_W(56, 373) <= 0; flappy_W(56, 374) <= 0; flappy_W(56, 375) <= 0; flappy_W(56, 376) <= 0; flappy_W(56, 377) <= 0; flappy_W(56, 378) <= 0; flappy_W(56, 379) <= 0; flappy_W(56, 380) <= 0; flappy_W(56, 381) <= 0; flappy_W(56, 382) <= 0; flappy_W(56, 383) <= 0; flappy_W(56, 384) <= 0; flappy_W(56, 385) <= 0; flappy_W(56, 386) <= 0; flappy_W(56, 387) <= 0; flappy_W(56, 388) <= 0; flappy_W(56, 389) <= 0; flappy_W(56, 390) <= 0; flappy_W(56, 391) <= 0; flappy_W(56, 392) <= 0; flappy_W(56, 393) <= 0; flappy_W(56, 394) <= 0; flappy_W(56, 395) <= 0; flappy_W(56, 396) <= 1; flappy_W(56, 397) <= 1; flappy_W(56, 398) <= 1; flappy_W(56, 399) <= 1; flappy_W(56, 400) <= 1; flappy_W(56, 401) <= 1; flappy_W(56, 402) <= 1; flappy_W(56, 403) <= 1; flappy_W(56, 404) <= 1; flappy_W(56, 405) <= 1; flappy_W(56, 406) <= 1; flappy_W(56, 407) <= 1; flappy_W(56, 408) <= 1; flappy_W(56, 409) <= 1; flappy_W(56, 410) <= 1; flappy_W(56, 411) <= 1; flappy_W(56, 412) <= 1; flappy_W(56, 413) <= 1; flappy_W(56, 414) <= 1; flappy_W(56, 415) <= 1; flappy_W(56, 416) <= 1; flappy_W(56, 417) <= 1; flappy_W(56, 418) <= 1; flappy_W(56, 419) <= 1; flappy_W(56, 420) <= 1; flappy_W(56, 421) <= 1; flappy_W(56, 422) <= 1; flappy_W(56, 423) <= 1; flappy_W(56, 424) <= 1; flappy_W(56, 425) <= 1; flappy_W(56, 426) <= 1; flappy_W(56, 427) <= 1; flappy_W(56, 428) <= 1; flappy_W(56, 429) <= 1; flappy_W(56, 430) <= 1; flappy_W(56, 431) <= 1; flappy_W(56, 432) <= 0; flappy_W(56, 433) <= 0; flappy_W(56, 434) <= 0; flappy_W(56, 435) <= 0; flappy_W(56, 436) <= 0; flappy_W(56, 437) <= 0; flappy_W(56, 438) <= 0; flappy_W(56, 439) <= 0; flappy_W(56, 440) <= 0; flappy_W(56, 441) <= 0; flappy_W(56, 442) <= 0; flappy_W(56, 443) <= 0; flappy_W(56, 444) <= 0; flappy_W(56, 445) <= 0; flappy_W(56, 446) <= 0; flappy_W(56, 447) <= 0; flappy_W(56, 448) <= 0; flappy_W(56, 449) <= 0; flappy_W(56, 450) <= 0; flappy_W(56, 451) <= 0; flappy_W(56, 452) <= 0; flappy_W(56, 453) <= 0; flappy_W(56, 454) <= 0; flappy_W(56, 455) <= 0; flappy_W(56, 456) <= 0; flappy_W(56, 457) <= 0; flappy_W(56, 458) <= 0; flappy_W(56, 459) <= 0; flappy_W(56, 460) <= 0; flappy_W(56, 461) <= 0; flappy_W(56, 462) <= 1; flappy_W(56, 463) <= 1; flappy_W(56, 464) <= 1; flappy_W(56, 465) <= 1; flappy_W(56, 466) <= 1; flappy_W(56, 467) <= 1; flappy_W(56, 468) <= 1; flappy_W(56, 469) <= 1; flappy_W(56, 470) <= 1; flappy_W(56, 471) <= 1; flappy_W(56, 472) <= 1; flappy_W(56, 473) <= 1; flappy_W(56, 474) <= 1; flappy_W(56, 475) <= 1; flappy_W(56, 476) <= 1; flappy_W(56, 477) <= 1; flappy_W(56, 478) <= 1; flappy_W(56, 479) <= 1; flappy_W(56, 480) <= 1; flappy_W(56, 481) <= 1; flappy_W(56, 482) <= 1; flappy_W(56, 483) <= 1; flappy_W(56, 484) <= 1; flappy_W(56, 485) <= 1; flappy_W(56, 486) <= 0; flappy_W(56, 487) <= 0; flappy_W(56, 488) <= 0; flappy_W(56, 489) <= 0; flappy_W(56, 490) <= 0; flappy_W(56, 491) <= 0; flappy_W(56, 492) <= 0; flappy_W(56, 493) <= 0; flappy_W(56, 494) <= 0; flappy_W(56, 495) <= 0; flappy_W(56, 496) <= 0; flappy_W(56, 497) <= 0; flappy_W(56, 498) <= 0; flappy_W(56, 499) <= 0; flappy_W(56, 500) <= 0; flappy_W(56, 501) <= 0; flappy_W(56, 502) <= 0; flappy_W(56, 503) <= 0; flappy_W(56, 504) <= 1; flappy_W(56, 505) <= 1; flappy_W(56, 506) <= 1; flappy_W(56, 507) <= 1; flappy_W(56, 508) <= 1; flappy_W(56, 509) <= 1; flappy_W(56, 510) <= 1; flappy_W(56, 511) <= 1; flappy_W(56, 512) <= 1; flappy_W(56, 513) <= 1; flappy_W(56, 514) <= 1; flappy_W(56, 515) <= 1; flappy_W(56, 516) <= 1; flappy_W(56, 517) <= 1; flappy_W(56, 518) <= 1; flappy_W(56, 519) <= 1; flappy_W(56, 520) <= 1; flappy_W(56, 521) <= 1; flappy_W(56, 522) <= 0; flappy_W(56, 523) <= 0; flappy_W(56, 524) <= 0; flappy_W(56, 525) <= 0; flappy_W(56, 526) <= 0; flappy_W(56, 527) <= 0; flappy_W(56, 528) <= 0; flappy_W(56, 529) <= 0; flappy_W(56, 530) <= 0; flappy_W(56, 531) <= 0; flappy_W(56, 532) <= 0; flappy_W(56, 533) <= 0; flappy_W(56, 534) <= 1; flappy_W(56, 535) <= 1; flappy_W(56, 536) <= 1; flappy_W(56, 537) <= 1; flappy_W(56, 538) <= 1; flappy_W(56, 539) <= 1; flappy_W(56, 540) <= 1; flappy_W(56, 541) <= 1; flappy_W(56, 542) <= 1; flappy_W(56, 543) <= 1; flappy_W(56, 544) <= 1; flappy_W(56, 545) <= 1; flappy_W(56, 546) <= 0; flappy_W(56, 547) <= 0; flappy_W(56, 548) <= 0; flappy_W(56, 549) <= 0; flappy_W(56, 550) <= 0; flappy_W(56, 551) <= 0; flappy_W(56, 552) <= 0; flappy_W(56, 553) <= 0; flappy_W(56, 554) <= 0; flappy_W(56, 555) <= 0; flappy_W(56, 556) <= 0; flappy_W(56, 557) <= 0; flappy_W(56, 558) <= 1; flappy_W(56, 559) <= 1; flappy_W(56, 560) <= 1; flappy_W(56, 561) <= 1; flappy_W(56, 562) <= 1; flappy_W(56, 563) <= 1; flappy_W(56, 564) <= 1; flappy_W(56, 565) <= 1; flappy_W(56, 566) <= 1; flappy_W(56, 567) <= 1; flappy_W(56, 568) <= 1; flappy_W(56, 569) <= 1; flappy_W(56, 570) <= 1; flappy_W(56, 571) <= 1; flappy_W(56, 572) <= 1; flappy_W(56, 573) <= 1; flappy_W(56, 574) <= 1; flappy_W(56, 575) <= 1; flappy_W(56, 576) <= 1; flappy_W(56, 577) <= 1; flappy_W(56, 578) <= 1; flappy_W(56, 579) <= 1; flappy_W(56, 580) <= 1; flappy_W(56, 581) <= 1; flappy_W(56, 582) <= 1; flappy_W(56, 583) <= 1; flappy_W(56, 584) <= 1; flappy_W(56, 585) <= 1; flappy_W(56, 586) <= 1; flappy_W(56, 587) <= 1; flappy_W(56, 588) <= 0; flappy_W(56, 589) <= 0; flappy_W(56, 590) <= 0; flappy_W(56, 591) <= 0; flappy_W(56, 592) <= 0; flappy_W(56, 593) <= 0; 
flappy_W(57, 0) <= 1; flappy_W(57, 1) <= 1; flappy_W(57, 2) <= 1; flappy_W(57, 3) <= 1; flappy_W(57, 4) <= 1; flappy_W(57, 5) <= 1; flappy_W(57, 6) <= 1; flappy_W(57, 7) <= 1; flappy_W(57, 8) <= 1; flappy_W(57, 9) <= 1; flappy_W(57, 10) <= 1; flappy_W(57, 11) <= 1; flappy_W(57, 12) <= 1; flappy_W(57, 13) <= 1; flappy_W(57, 14) <= 1; flappy_W(57, 15) <= 1; flappy_W(57, 16) <= 1; flappy_W(57, 17) <= 1; flappy_W(57, 18) <= 1; flappy_W(57, 19) <= 1; flappy_W(57, 20) <= 1; flappy_W(57, 21) <= 1; flappy_W(57, 22) <= 1; flappy_W(57, 23) <= 1; flappy_W(57, 24) <= 0; flappy_W(57, 25) <= 0; flappy_W(57, 26) <= 0; flappy_W(57, 27) <= 0; flappy_W(57, 28) <= 0; flappy_W(57, 29) <= 0; flappy_W(57, 30) <= 0; flappy_W(57, 31) <= 0; flappy_W(57, 32) <= 0; flappy_W(57, 33) <= 0; flappy_W(57, 34) <= 0; flappy_W(57, 35) <= 0; flappy_W(57, 36) <= 0; flappy_W(57, 37) <= 0; flappy_W(57, 38) <= 0; flappy_W(57, 39) <= 0; flappy_W(57, 40) <= 0; flappy_W(57, 41) <= 0; flappy_W(57, 42) <= 0; flappy_W(57, 43) <= 0; flappy_W(57, 44) <= 0; flappy_W(57, 45) <= 0; flappy_W(57, 46) <= 0; flappy_W(57, 47) <= 0; flappy_W(57, 48) <= 0; flappy_W(57, 49) <= 0; flappy_W(57, 50) <= 0; flappy_W(57, 51) <= 0; flappy_W(57, 52) <= 0; flappy_W(57, 53) <= 0; flappy_W(57, 54) <= 1; flappy_W(57, 55) <= 1; flappy_W(57, 56) <= 1; flappy_W(57, 57) <= 1; flappy_W(57, 58) <= 1; flappy_W(57, 59) <= 1; flappy_W(57, 60) <= 1; flappy_W(57, 61) <= 1; flappy_W(57, 62) <= 1; flappy_W(57, 63) <= 1; flappy_W(57, 64) <= 1; flappy_W(57, 65) <= 1; flappy_W(57, 66) <= 1; flappy_W(57, 67) <= 1; flappy_W(57, 68) <= 1; flappy_W(57, 69) <= 1; flappy_W(57, 70) <= 1; flappy_W(57, 71) <= 1; flappy_W(57, 72) <= 1; flappy_W(57, 73) <= 1; flappy_W(57, 74) <= 1; flappy_W(57, 75) <= 1; flappy_W(57, 76) <= 1; flappy_W(57, 77) <= 1; flappy_W(57, 78) <= 1; flappy_W(57, 79) <= 1; flappy_W(57, 80) <= 1; flappy_W(57, 81) <= 1; flappy_W(57, 82) <= 1; flappy_W(57, 83) <= 1; flappy_W(57, 84) <= 1; flappy_W(57, 85) <= 1; flappy_W(57, 86) <= 1; flappy_W(57, 87) <= 1; flappy_W(57, 88) <= 1; flappy_W(57, 89) <= 1; flappy_W(57, 90) <= 1; flappy_W(57, 91) <= 1; flappy_W(57, 92) <= 1; flappy_W(57, 93) <= 1; flappy_W(57, 94) <= 1; flappy_W(57, 95) <= 1; flappy_W(57, 96) <= 0; flappy_W(57, 97) <= 0; flappy_W(57, 98) <= 0; flappy_W(57, 99) <= 0; flappy_W(57, 100) <= 0; flappy_W(57, 101) <= 0; flappy_W(57, 102) <= 0; flappy_W(57, 103) <= 0; flappy_W(57, 104) <= 0; flappy_W(57, 105) <= 0; flappy_W(57, 106) <= 0; flappy_W(57, 107) <= 0; flappy_W(57, 108) <= 1; flappy_W(57, 109) <= 1; flappy_W(57, 110) <= 1; flappy_W(57, 111) <= 1; flappy_W(57, 112) <= 1; flappy_W(57, 113) <= 1; flappy_W(57, 114) <= 1; flappy_W(57, 115) <= 1; flappy_W(57, 116) <= 1; flappy_W(57, 117) <= 1; flappy_W(57, 118) <= 1; flappy_W(57, 119) <= 1; flappy_W(57, 120) <= 0; flappy_W(57, 121) <= 0; flappy_W(57, 122) <= 0; flappy_W(57, 123) <= 0; flappy_W(57, 124) <= 0; flappy_W(57, 125) <= 0; flappy_W(57, 126) <= 0; flappy_W(57, 127) <= 0; flappy_W(57, 128) <= 0; flappy_W(57, 129) <= 0; flappy_W(57, 130) <= 0; flappy_W(57, 131) <= 0; flappy_W(57, 132) <= 0; flappy_W(57, 133) <= 0; flappy_W(57, 134) <= 0; flappy_W(57, 135) <= 0; flappy_W(57, 136) <= 0; flappy_W(57, 137) <= 0; flappy_W(57, 138) <= 1; flappy_W(57, 139) <= 1; flappy_W(57, 140) <= 1; flappy_W(57, 141) <= 1; flappy_W(57, 142) <= 1; flappy_W(57, 143) <= 1; flappy_W(57, 144) <= 1; flappy_W(57, 145) <= 1; flappy_W(57, 146) <= 1; flappy_W(57, 147) <= 1; flappy_W(57, 148) <= 1; flappy_W(57, 149) <= 1; flappy_W(57, 150) <= 0; flappy_W(57, 151) <= 0; flappy_W(57, 152) <= 0; flappy_W(57, 153) <= 0; flappy_W(57, 154) <= 0; flappy_W(57, 155) <= 0; flappy_W(57, 156) <= 0; flappy_W(57, 157) <= 0; flappy_W(57, 158) <= 0; flappy_W(57, 159) <= 0; flappy_W(57, 160) <= 0; flappy_W(57, 161) <= 0; flappy_W(57, 162) <= 1; flappy_W(57, 163) <= 1; flappy_W(57, 164) <= 1; flappy_W(57, 165) <= 1; flappy_W(57, 166) <= 1; flappy_W(57, 167) <= 1; flappy_W(57, 168) <= 1; flappy_W(57, 169) <= 1; flappy_W(57, 170) <= 1; flappy_W(57, 171) <= 1; flappy_W(57, 172) <= 1; flappy_W(57, 173) <= 1; flappy_W(57, 174) <= 1; flappy_W(57, 175) <= 1; flappy_W(57, 176) <= 1; flappy_W(57, 177) <= 1; flappy_W(57, 178) <= 1; flappy_W(57, 179) <= 1; flappy_W(57, 180) <= 1; flappy_W(57, 181) <= 1; flappy_W(57, 182) <= 1; flappy_W(57, 183) <= 1; flappy_W(57, 184) <= 1; flappy_W(57, 185) <= 1; flappy_W(57, 186) <= 0; flappy_W(57, 187) <= 0; flappy_W(57, 188) <= 0; flappy_W(57, 189) <= 0; flappy_W(57, 190) <= 0; flappy_W(57, 191) <= 0; flappy_W(57, 192) <= 0; flappy_W(57, 193) <= 0; flappy_W(57, 194) <= 0; flappy_W(57, 195) <= 0; flappy_W(57, 196) <= 0; flappy_W(57, 197) <= 0; flappy_W(57, 198) <= 0; flappy_W(57, 199) <= 0; flappy_W(57, 200) <= 0; flappy_W(57, 201) <= 0; flappy_W(57, 202) <= 0; flappy_W(57, 203) <= 0; flappy_W(57, 204) <= 0; flappy_W(57, 205) <= 0; flappy_W(57, 206) <= 0; flappy_W(57, 207) <= 0; flappy_W(57, 208) <= 0; flappy_W(57, 209) <= 0; flappy_W(57, 210) <= 0; flappy_W(57, 211) <= 0; flappy_W(57, 212) <= 0; flappy_W(57, 213) <= 0; flappy_W(57, 214) <= 0; flappy_W(57, 215) <= 0; flappy_W(57, 216) <= 1; flappy_W(57, 217) <= 1; flappy_W(57, 218) <= 1; flappy_W(57, 219) <= 1; flappy_W(57, 220) <= 1; flappy_W(57, 221) <= 1; flappy_W(57, 222) <= 1; flappy_W(57, 223) <= 1; flappy_W(57, 224) <= 1; flappy_W(57, 225) <= 1; flappy_W(57, 226) <= 1; flappy_W(57, 227) <= 1; flappy_W(57, 228) <= 1; flappy_W(57, 229) <= 1; flappy_W(57, 230) <= 1; flappy_W(57, 231) <= 1; flappy_W(57, 232) <= 1; flappy_W(57, 233) <= 1; flappy_W(57, 234) <= 1; flappy_W(57, 235) <= 1; flappy_W(57, 236) <= 1; flappy_W(57, 237) <= 1; flappy_W(57, 238) <= 1; flappy_W(57, 239) <= 1; flappy_W(57, 240) <= 0; flappy_W(57, 241) <= 0; flappy_W(57, 242) <= 0; flappy_W(57, 243) <= 0; flappy_W(57, 244) <= 0; flappy_W(57, 245) <= 0; flappy_W(57, 246) <= 0; flappy_W(57, 247) <= 0; flappy_W(57, 248) <= 0; flappy_W(57, 249) <= 0; flappy_W(57, 250) <= 0; flappy_W(57, 251) <= 0; flappy_W(57, 252) <= 0; flappy_W(57, 253) <= 0; flappy_W(57, 254) <= 0; flappy_W(57, 255) <= 0; flappy_W(57, 256) <= 0; flappy_W(57, 257) <= 0; flappy_W(57, 258) <= 0; flappy_W(57, 259) <= 0; flappy_W(57, 260) <= 0; flappy_W(57, 261) <= 0; flappy_W(57, 262) <= 0; flappy_W(57, 263) <= 0; flappy_W(57, 264) <= 0; flappy_W(57, 265) <= 0; flappy_W(57, 266) <= 0; flappy_W(57, 267) <= 0; flappy_W(57, 268) <= 0; flappy_W(57, 269) <= 0; flappy_W(57, 270) <= 0; flappy_W(57, 271) <= 0; flappy_W(57, 272) <= 0; flappy_W(57, 273) <= 0; flappy_W(57, 274) <= 0; flappy_W(57, 275) <= 0; flappy_W(57, 276) <= 0; flappy_W(57, 277) <= 0; flappy_W(57, 278) <= 0; flappy_W(57, 279) <= 0; flappy_W(57, 280) <= 0; flappy_W(57, 281) <= 0; flappy_W(57, 282) <= 1; flappy_W(57, 283) <= 1; flappy_W(57, 284) <= 1; flappy_W(57, 285) <= 1; flappy_W(57, 286) <= 1; flappy_W(57, 287) <= 1; flappy_W(57, 288) <= 1; flappy_W(57, 289) <= 1; flappy_W(57, 290) <= 1; flappy_W(57, 291) <= 1; flappy_W(57, 292) <= 1; flappy_W(57, 293) <= 1; flappy_W(57, 294) <= 1; flappy_W(57, 295) <= 1; flappy_W(57, 296) <= 1; flappy_W(57, 297) <= 1; flappy_W(57, 298) <= 1; flappy_W(57, 299) <= 1; flappy_W(57, 300) <= 1; flappy_W(57, 301) <= 1; flappy_W(57, 302) <= 1; flappy_W(57, 303) <= 1; flappy_W(57, 304) <= 1; flappy_W(57, 305) <= 1; flappy_W(57, 306) <= 0; flappy_W(57, 307) <= 0; flappy_W(57, 308) <= 0; flappy_W(57, 309) <= 0; flappy_W(57, 310) <= 0; flappy_W(57, 311) <= 0; flappy_W(57, 312) <= 0; flappy_W(57, 313) <= 0; flappy_W(57, 314) <= 0; flappy_W(57, 315) <= 0; flappy_W(57, 316) <= 0; flappy_W(57, 317) <= 0; flappy_W(57, 318) <= 0; flappy_W(57, 319) <= 0; flappy_W(57, 320) <= 0; flappy_W(57, 321) <= 0; flappy_W(57, 322) <= 0; flappy_W(57, 323) <= 0; flappy_W(57, 324) <= 0; flappy_W(57, 325) <= 0; flappy_W(57, 326) <= 0; flappy_W(57, 327) <= 0; flappy_W(57, 328) <= 0; flappy_W(57, 329) <= 0; flappy_W(57, 330) <= 0; flappy_W(57, 331) <= 0; flappy_W(57, 332) <= 0; flappy_W(57, 333) <= 0; flappy_W(57, 334) <= 0; flappy_W(57, 335) <= 0; flappy_W(57, 336) <= 0; flappy_W(57, 337) <= 0; flappy_W(57, 338) <= 0; flappy_W(57, 339) <= 0; flappy_W(57, 340) <= 0; flappy_W(57, 341) <= 0; flappy_W(57, 342) <= 0; flappy_W(57, 343) <= 0; flappy_W(57, 344) <= 0; flappy_W(57, 345) <= 0; flappy_W(57, 346) <= 0; flappy_W(57, 347) <= 0; flappy_W(57, 348) <= 0; flappy_W(57, 349) <= 0; flappy_W(57, 350) <= 0; flappy_W(57, 351) <= 0; flappy_W(57, 352) <= 0; flappy_W(57, 353) <= 0; flappy_W(57, 354) <= 0; flappy_W(57, 355) <= 0; flappy_W(57, 356) <= 0; flappy_W(57, 357) <= 0; flappy_W(57, 358) <= 0; flappy_W(57, 359) <= 0; flappy_W(57, 360) <= 0; flappy_W(57, 361) <= 0; flappy_W(57, 362) <= 0; flappy_W(57, 363) <= 0; flappy_W(57, 364) <= 0; flappy_W(57, 365) <= 0; flappy_W(57, 366) <= 0; flappy_W(57, 367) <= 0; flappy_W(57, 368) <= 0; flappy_W(57, 369) <= 0; flappy_W(57, 370) <= 0; flappy_W(57, 371) <= 0; flappy_W(57, 372) <= 0; flappy_W(57, 373) <= 0; flappy_W(57, 374) <= 0; flappy_W(57, 375) <= 0; flappy_W(57, 376) <= 0; flappy_W(57, 377) <= 0; flappy_W(57, 378) <= 0; flappy_W(57, 379) <= 0; flappy_W(57, 380) <= 0; flappy_W(57, 381) <= 0; flappy_W(57, 382) <= 0; flappy_W(57, 383) <= 0; flappy_W(57, 384) <= 0; flappy_W(57, 385) <= 0; flappy_W(57, 386) <= 0; flappy_W(57, 387) <= 0; flappy_W(57, 388) <= 0; flappy_W(57, 389) <= 0; flappy_W(57, 390) <= 0; flappy_W(57, 391) <= 0; flappy_W(57, 392) <= 0; flappy_W(57, 393) <= 0; flappy_W(57, 394) <= 0; flappy_W(57, 395) <= 0; flappy_W(57, 396) <= 1; flappy_W(57, 397) <= 1; flappy_W(57, 398) <= 1; flappy_W(57, 399) <= 1; flappy_W(57, 400) <= 1; flappy_W(57, 401) <= 1; flappy_W(57, 402) <= 1; flappy_W(57, 403) <= 1; flappy_W(57, 404) <= 1; flappy_W(57, 405) <= 1; flappy_W(57, 406) <= 1; flappy_W(57, 407) <= 1; flappy_W(57, 408) <= 1; flappy_W(57, 409) <= 1; flappy_W(57, 410) <= 1; flappy_W(57, 411) <= 1; flappy_W(57, 412) <= 1; flappy_W(57, 413) <= 1; flappy_W(57, 414) <= 1; flappy_W(57, 415) <= 1; flappy_W(57, 416) <= 1; flappy_W(57, 417) <= 1; flappy_W(57, 418) <= 1; flappy_W(57, 419) <= 1; flappy_W(57, 420) <= 1; flappy_W(57, 421) <= 1; flappy_W(57, 422) <= 1; flappy_W(57, 423) <= 1; flappy_W(57, 424) <= 1; flappy_W(57, 425) <= 1; flappy_W(57, 426) <= 1; flappy_W(57, 427) <= 1; flappy_W(57, 428) <= 1; flappy_W(57, 429) <= 1; flappy_W(57, 430) <= 1; flappy_W(57, 431) <= 1; flappy_W(57, 432) <= 0; flappy_W(57, 433) <= 0; flappy_W(57, 434) <= 0; flappy_W(57, 435) <= 0; flappy_W(57, 436) <= 0; flappy_W(57, 437) <= 0; flappy_W(57, 438) <= 0; flappy_W(57, 439) <= 0; flappy_W(57, 440) <= 0; flappy_W(57, 441) <= 0; flappy_W(57, 442) <= 0; flappy_W(57, 443) <= 0; flappy_W(57, 444) <= 0; flappy_W(57, 445) <= 0; flappy_W(57, 446) <= 0; flappy_W(57, 447) <= 0; flappy_W(57, 448) <= 0; flappy_W(57, 449) <= 0; flappy_W(57, 450) <= 0; flappy_W(57, 451) <= 0; flappy_W(57, 452) <= 0; flappy_W(57, 453) <= 0; flappy_W(57, 454) <= 0; flappy_W(57, 455) <= 0; flappy_W(57, 456) <= 0; flappy_W(57, 457) <= 0; flappy_W(57, 458) <= 0; flappy_W(57, 459) <= 0; flappy_W(57, 460) <= 0; flappy_W(57, 461) <= 0; flappy_W(57, 462) <= 1; flappy_W(57, 463) <= 1; flappy_W(57, 464) <= 1; flappy_W(57, 465) <= 1; flappy_W(57, 466) <= 1; flappy_W(57, 467) <= 1; flappy_W(57, 468) <= 1; flappy_W(57, 469) <= 1; flappy_W(57, 470) <= 1; flappy_W(57, 471) <= 1; flappy_W(57, 472) <= 1; flappy_W(57, 473) <= 1; flappy_W(57, 474) <= 1; flappy_W(57, 475) <= 1; flappy_W(57, 476) <= 1; flappy_W(57, 477) <= 1; flappy_W(57, 478) <= 1; flappy_W(57, 479) <= 1; flappy_W(57, 480) <= 1; flappy_W(57, 481) <= 1; flappy_W(57, 482) <= 1; flappy_W(57, 483) <= 1; flappy_W(57, 484) <= 1; flappy_W(57, 485) <= 1; flappy_W(57, 486) <= 0; flappy_W(57, 487) <= 0; flappy_W(57, 488) <= 0; flappy_W(57, 489) <= 0; flappy_W(57, 490) <= 0; flappy_W(57, 491) <= 0; flappy_W(57, 492) <= 0; flappy_W(57, 493) <= 0; flappy_W(57, 494) <= 0; flappy_W(57, 495) <= 0; flappy_W(57, 496) <= 0; flappy_W(57, 497) <= 0; flappy_W(57, 498) <= 0; flappy_W(57, 499) <= 0; flappy_W(57, 500) <= 0; flappy_W(57, 501) <= 0; flappy_W(57, 502) <= 0; flappy_W(57, 503) <= 0; flappy_W(57, 504) <= 1; flappy_W(57, 505) <= 1; flappy_W(57, 506) <= 1; flappy_W(57, 507) <= 1; flappy_W(57, 508) <= 1; flappy_W(57, 509) <= 1; flappy_W(57, 510) <= 1; flappy_W(57, 511) <= 1; flappy_W(57, 512) <= 1; flappy_W(57, 513) <= 1; flappy_W(57, 514) <= 1; flappy_W(57, 515) <= 1; flappy_W(57, 516) <= 1; flappy_W(57, 517) <= 1; flappy_W(57, 518) <= 1; flappy_W(57, 519) <= 1; flappy_W(57, 520) <= 1; flappy_W(57, 521) <= 1; flappy_W(57, 522) <= 0; flappy_W(57, 523) <= 0; flappy_W(57, 524) <= 0; flappy_W(57, 525) <= 0; flappy_W(57, 526) <= 0; flappy_W(57, 527) <= 0; flappy_W(57, 528) <= 0; flappy_W(57, 529) <= 0; flappy_W(57, 530) <= 0; flappy_W(57, 531) <= 0; flappy_W(57, 532) <= 0; flappy_W(57, 533) <= 0; flappy_W(57, 534) <= 1; flappy_W(57, 535) <= 1; flappy_W(57, 536) <= 1; flappy_W(57, 537) <= 1; flappy_W(57, 538) <= 1; flappy_W(57, 539) <= 1; flappy_W(57, 540) <= 1; flappy_W(57, 541) <= 1; flappy_W(57, 542) <= 1; flappy_W(57, 543) <= 1; flappy_W(57, 544) <= 1; flappy_W(57, 545) <= 1; flappy_W(57, 546) <= 0; flappy_W(57, 547) <= 0; flappy_W(57, 548) <= 0; flappy_W(57, 549) <= 0; flappy_W(57, 550) <= 0; flappy_W(57, 551) <= 0; flappy_W(57, 552) <= 0; flappy_W(57, 553) <= 0; flappy_W(57, 554) <= 0; flappy_W(57, 555) <= 0; flappy_W(57, 556) <= 0; flappy_W(57, 557) <= 0; flappy_W(57, 558) <= 1; flappy_W(57, 559) <= 1; flappy_W(57, 560) <= 1; flappy_W(57, 561) <= 1; flappy_W(57, 562) <= 1; flappy_W(57, 563) <= 1; flappy_W(57, 564) <= 1; flappy_W(57, 565) <= 1; flappy_W(57, 566) <= 1; flappy_W(57, 567) <= 1; flappy_W(57, 568) <= 1; flappy_W(57, 569) <= 1; flappy_W(57, 570) <= 1; flappy_W(57, 571) <= 1; flappy_W(57, 572) <= 1; flappy_W(57, 573) <= 1; flappy_W(57, 574) <= 1; flappy_W(57, 575) <= 1; flappy_W(57, 576) <= 1; flappy_W(57, 577) <= 1; flappy_W(57, 578) <= 1; flappy_W(57, 579) <= 1; flappy_W(57, 580) <= 1; flappy_W(57, 581) <= 1; flappy_W(57, 582) <= 1; flappy_W(57, 583) <= 1; flappy_W(57, 584) <= 1; flappy_W(57, 585) <= 1; flappy_W(57, 586) <= 1; flappy_W(57, 587) <= 1; flappy_W(57, 588) <= 0; flappy_W(57, 589) <= 0; flappy_W(57, 590) <= 0; flappy_W(57, 591) <= 0; flappy_W(57, 592) <= 0; flappy_W(57, 593) <= 0; 
flappy_W(58, 0) <= 1; flappy_W(58, 1) <= 1; flappy_W(58, 2) <= 1; flappy_W(58, 3) <= 1; flappy_W(58, 4) <= 1; flappy_W(58, 5) <= 1; flappy_W(58, 6) <= 1; flappy_W(58, 7) <= 1; flappy_W(58, 8) <= 1; flappy_W(58, 9) <= 1; flappy_W(58, 10) <= 1; flappy_W(58, 11) <= 1; flappy_W(58, 12) <= 1; flappy_W(58, 13) <= 1; flappy_W(58, 14) <= 1; flappy_W(58, 15) <= 1; flappy_W(58, 16) <= 1; flappy_W(58, 17) <= 1; flappy_W(58, 18) <= 1; flappy_W(58, 19) <= 1; flappy_W(58, 20) <= 1; flappy_W(58, 21) <= 1; flappy_W(58, 22) <= 1; flappy_W(58, 23) <= 1; flappy_W(58, 24) <= 0; flappy_W(58, 25) <= 0; flappy_W(58, 26) <= 0; flappy_W(58, 27) <= 0; flappy_W(58, 28) <= 0; flappy_W(58, 29) <= 0; flappy_W(58, 30) <= 0; flappy_W(58, 31) <= 0; flappy_W(58, 32) <= 0; flappy_W(58, 33) <= 0; flappy_W(58, 34) <= 0; flappy_W(58, 35) <= 0; flappy_W(58, 36) <= 0; flappy_W(58, 37) <= 0; flappy_W(58, 38) <= 0; flappy_W(58, 39) <= 0; flappy_W(58, 40) <= 0; flappy_W(58, 41) <= 0; flappy_W(58, 42) <= 0; flappy_W(58, 43) <= 0; flappy_W(58, 44) <= 0; flappy_W(58, 45) <= 0; flappy_W(58, 46) <= 0; flappy_W(58, 47) <= 0; flappy_W(58, 48) <= 0; flappy_W(58, 49) <= 0; flappy_W(58, 50) <= 0; flappy_W(58, 51) <= 0; flappy_W(58, 52) <= 0; flappy_W(58, 53) <= 0; flappy_W(58, 54) <= 1; flappy_W(58, 55) <= 1; flappy_W(58, 56) <= 1; flappy_W(58, 57) <= 1; flappy_W(58, 58) <= 1; flappy_W(58, 59) <= 1; flappy_W(58, 60) <= 1; flappy_W(58, 61) <= 1; flappy_W(58, 62) <= 1; flappy_W(58, 63) <= 1; flappy_W(58, 64) <= 1; flappy_W(58, 65) <= 1; flappy_W(58, 66) <= 1; flappy_W(58, 67) <= 1; flappy_W(58, 68) <= 1; flappy_W(58, 69) <= 1; flappy_W(58, 70) <= 1; flappy_W(58, 71) <= 1; flappy_W(58, 72) <= 1; flappy_W(58, 73) <= 1; flappy_W(58, 74) <= 1; flappy_W(58, 75) <= 1; flappy_W(58, 76) <= 1; flappy_W(58, 77) <= 1; flappy_W(58, 78) <= 1; flappy_W(58, 79) <= 1; flappy_W(58, 80) <= 1; flappy_W(58, 81) <= 1; flappy_W(58, 82) <= 1; flappy_W(58, 83) <= 1; flappy_W(58, 84) <= 1; flappy_W(58, 85) <= 1; flappy_W(58, 86) <= 1; flappy_W(58, 87) <= 1; flappy_W(58, 88) <= 1; flappy_W(58, 89) <= 1; flappy_W(58, 90) <= 1; flappy_W(58, 91) <= 1; flappy_W(58, 92) <= 1; flappy_W(58, 93) <= 1; flappy_W(58, 94) <= 1; flappy_W(58, 95) <= 1; flappy_W(58, 96) <= 0; flappy_W(58, 97) <= 0; flappy_W(58, 98) <= 0; flappy_W(58, 99) <= 0; flappy_W(58, 100) <= 0; flappy_W(58, 101) <= 0; flappy_W(58, 102) <= 0; flappy_W(58, 103) <= 0; flappy_W(58, 104) <= 0; flappy_W(58, 105) <= 0; flappy_W(58, 106) <= 0; flappy_W(58, 107) <= 0; flappy_W(58, 108) <= 1; flappy_W(58, 109) <= 1; flappy_W(58, 110) <= 1; flappy_W(58, 111) <= 1; flappy_W(58, 112) <= 1; flappy_W(58, 113) <= 1; flappy_W(58, 114) <= 1; flappy_W(58, 115) <= 1; flappy_W(58, 116) <= 1; flappy_W(58, 117) <= 1; flappy_W(58, 118) <= 1; flappy_W(58, 119) <= 1; flappy_W(58, 120) <= 0; flappy_W(58, 121) <= 0; flappy_W(58, 122) <= 0; flappy_W(58, 123) <= 0; flappy_W(58, 124) <= 0; flappy_W(58, 125) <= 0; flappy_W(58, 126) <= 0; flappy_W(58, 127) <= 0; flappy_W(58, 128) <= 0; flappy_W(58, 129) <= 0; flappy_W(58, 130) <= 0; flappy_W(58, 131) <= 0; flappy_W(58, 132) <= 0; flappy_W(58, 133) <= 0; flappy_W(58, 134) <= 0; flappy_W(58, 135) <= 0; flappy_W(58, 136) <= 0; flappy_W(58, 137) <= 0; flappy_W(58, 138) <= 1; flappy_W(58, 139) <= 1; flappy_W(58, 140) <= 1; flappy_W(58, 141) <= 1; flappy_W(58, 142) <= 1; flappy_W(58, 143) <= 1; flappy_W(58, 144) <= 1; flappy_W(58, 145) <= 1; flappy_W(58, 146) <= 1; flappy_W(58, 147) <= 1; flappy_W(58, 148) <= 1; flappy_W(58, 149) <= 1; flappy_W(58, 150) <= 0; flappy_W(58, 151) <= 0; flappy_W(58, 152) <= 0; flappy_W(58, 153) <= 0; flappy_W(58, 154) <= 0; flappy_W(58, 155) <= 0; flappy_W(58, 156) <= 0; flappy_W(58, 157) <= 0; flappy_W(58, 158) <= 0; flappy_W(58, 159) <= 0; flappy_W(58, 160) <= 0; flappy_W(58, 161) <= 0; flappy_W(58, 162) <= 1; flappy_W(58, 163) <= 1; flappy_W(58, 164) <= 1; flappy_W(58, 165) <= 1; flappy_W(58, 166) <= 1; flappy_W(58, 167) <= 1; flappy_W(58, 168) <= 1; flappy_W(58, 169) <= 1; flappy_W(58, 170) <= 1; flappy_W(58, 171) <= 1; flappy_W(58, 172) <= 1; flappy_W(58, 173) <= 1; flappy_W(58, 174) <= 1; flappy_W(58, 175) <= 1; flappy_W(58, 176) <= 1; flappy_W(58, 177) <= 1; flappy_W(58, 178) <= 1; flappy_W(58, 179) <= 1; flappy_W(58, 180) <= 1; flappy_W(58, 181) <= 1; flappy_W(58, 182) <= 1; flappy_W(58, 183) <= 1; flappy_W(58, 184) <= 1; flappy_W(58, 185) <= 1; flappy_W(58, 186) <= 0; flappy_W(58, 187) <= 0; flappy_W(58, 188) <= 0; flappy_W(58, 189) <= 0; flappy_W(58, 190) <= 0; flappy_W(58, 191) <= 0; flappy_W(58, 192) <= 0; flappy_W(58, 193) <= 0; flappy_W(58, 194) <= 0; flappy_W(58, 195) <= 0; flappy_W(58, 196) <= 0; flappy_W(58, 197) <= 0; flappy_W(58, 198) <= 0; flappy_W(58, 199) <= 0; flappy_W(58, 200) <= 0; flappy_W(58, 201) <= 0; flappy_W(58, 202) <= 0; flappy_W(58, 203) <= 0; flappy_W(58, 204) <= 0; flappy_W(58, 205) <= 0; flappy_W(58, 206) <= 0; flappy_W(58, 207) <= 0; flappy_W(58, 208) <= 0; flappy_W(58, 209) <= 0; flappy_W(58, 210) <= 0; flappy_W(58, 211) <= 0; flappy_W(58, 212) <= 0; flappy_W(58, 213) <= 0; flappy_W(58, 214) <= 0; flappy_W(58, 215) <= 0; flappy_W(58, 216) <= 1; flappy_W(58, 217) <= 1; flappy_W(58, 218) <= 1; flappy_W(58, 219) <= 1; flappy_W(58, 220) <= 1; flappy_W(58, 221) <= 1; flappy_W(58, 222) <= 1; flappy_W(58, 223) <= 1; flappy_W(58, 224) <= 1; flappy_W(58, 225) <= 1; flappy_W(58, 226) <= 1; flappy_W(58, 227) <= 1; flappy_W(58, 228) <= 1; flappy_W(58, 229) <= 1; flappy_W(58, 230) <= 1; flappy_W(58, 231) <= 1; flappy_W(58, 232) <= 1; flappy_W(58, 233) <= 1; flappy_W(58, 234) <= 1; flappy_W(58, 235) <= 1; flappy_W(58, 236) <= 1; flappy_W(58, 237) <= 1; flappy_W(58, 238) <= 1; flappy_W(58, 239) <= 1; flappy_W(58, 240) <= 0; flappy_W(58, 241) <= 0; flappy_W(58, 242) <= 0; flappy_W(58, 243) <= 0; flappy_W(58, 244) <= 0; flappy_W(58, 245) <= 0; flappy_W(58, 246) <= 0; flappy_W(58, 247) <= 0; flappy_W(58, 248) <= 0; flappy_W(58, 249) <= 0; flappy_W(58, 250) <= 0; flappy_W(58, 251) <= 0; flappy_W(58, 252) <= 0; flappy_W(58, 253) <= 0; flappy_W(58, 254) <= 0; flappy_W(58, 255) <= 0; flappy_W(58, 256) <= 0; flappy_W(58, 257) <= 0; flappy_W(58, 258) <= 0; flappy_W(58, 259) <= 0; flappy_W(58, 260) <= 0; flappy_W(58, 261) <= 0; flappy_W(58, 262) <= 0; flappy_W(58, 263) <= 0; flappy_W(58, 264) <= 0; flappy_W(58, 265) <= 0; flappy_W(58, 266) <= 0; flappy_W(58, 267) <= 0; flappy_W(58, 268) <= 0; flappy_W(58, 269) <= 0; flappy_W(58, 270) <= 0; flappy_W(58, 271) <= 0; flappy_W(58, 272) <= 0; flappy_W(58, 273) <= 0; flappy_W(58, 274) <= 0; flappy_W(58, 275) <= 0; flappy_W(58, 276) <= 0; flappy_W(58, 277) <= 0; flappy_W(58, 278) <= 0; flappy_W(58, 279) <= 0; flappy_W(58, 280) <= 0; flappy_W(58, 281) <= 0; flappy_W(58, 282) <= 1; flappy_W(58, 283) <= 1; flappy_W(58, 284) <= 1; flappy_W(58, 285) <= 1; flappy_W(58, 286) <= 1; flappy_W(58, 287) <= 1; flappy_W(58, 288) <= 1; flappy_W(58, 289) <= 1; flappy_W(58, 290) <= 1; flappy_W(58, 291) <= 1; flappy_W(58, 292) <= 1; flappy_W(58, 293) <= 1; flappy_W(58, 294) <= 1; flappy_W(58, 295) <= 1; flappy_W(58, 296) <= 1; flappy_W(58, 297) <= 1; flappy_W(58, 298) <= 1; flappy_W(58, 299) <= 1; flappy_W(58, 300) <= 1; flappy_W(58, 301) <= 1; flappy_W(58, 302) <= 1; flappy_W(58, 303) <= 1; flappy_W(58, 304) <= 1; flappy_W(58, 305) <= 1; flappy_W(58, 306) <= 0; flappy_W(58, 307) <= 0; flappy_W(58, 308) <= 0; flappy_W(58, 309) <= 0; flappy_W(58, 310) <= 0; flappy_W(58, 311) <= 0; flappy_W(58, 312) <= 0; flappy_W(58, 313) <= 0; flappy_W(58, 314) <= 0; flappy_W(58, 315) <= 0; flappy_W(58, 316) <= 0; flappy_W(58, 317) <= 0; flappy_W(58, 318) <= 0; flappy_W(58, 319) <= 0; flappy_W(58, 320) <= 0; flappy_W(58, 321) <= 0; flappy_W(58, 322) <= 0; flappy_W(58, 323) <= 0; flappy_W(58, 324) <= 0; flappy_W(58, 325) <= 0; flappy_W(58, 326) <= 0; flappy_W(58, 327) <= 0; flappy_W(58, 328) <= 0; flappy_W(58, 329) <= 0; flappy_W(58, 330) <= 0; flappy_W(58, 331) <= 0; flappy_W(58, 332) <= 0; flappy_W(58, 333) <= 0; flappy_W(58, 334) <= 0; flappy_W(58, 335) <= 0; flappy_W(58, 336) <= 0; flappy_W(58, 337) <= 0; flappy_W(58, 338) <= 0; flappy_W(58, 339) <= 0; flappy_W(58, 340) <= 0; flappy_W(58, 341) <= 0; flappy_W(58, 342) <= 0; flappy_W(58, 343) <= 0; flappy_W(58, 344) <= 0; flappy_W(58, 345) <= 0; flappy_W(58, 346) <= 0; flappy_W(58, 347) <= 0; flappy_W(58, 348) <= 0; flappy_W(58, 349) <= 0; flappy_W(58, 350) <= 0; flappy_W(58, 351) <= 0; flappy_W(58, 352) <= 0; flappy_W(58, 353) <= 0; flappy_W(58, 354) <= 0; flappy_W(58, 355) <= 0; flappy_W(58, 356) <= 0; flappy_W(58, 357) <= 0; flappy_W(58, 358) <= 0; flappy_W(58, 359) <= 0; flappy_W(58, 360) <= 0; flappy_W(58, 361) <= 0; flappy_W(58, 362) <= 0; flappy_W(58, 363) <= 0; flappy_W(58, 364) <= 0; flappy_W(58, 365) <= 0; flappy_W(58, 366) <= 0; flappy_W(58, 367) <= 0; flappy_W(58, 368) <= 0; flappy_W(58, 369) <= 0; flappy_W(58, 370) <= 0; flappy_W(58, 371) <= 0; flappy_W(58, 372) <= 0; flappy_W(58, 373) <= 0; flappy_W(58, 374) <= 0; flappy_W(58, 375) <= 0; flappy_W(58, 376) <= 0; flappy_W(58, 377) <= 0; flappy_W(58, 378) <= 0; flappy_W(58, 379) <= 0; flappy_W(58, 380) <= 0; flappy_W(58, 381) <= 0; flappy_W(58, 382) <= 0; flappy_W(58, 383) <= 0; flappy_W(58, 384) <= 0; flappy_W(58, 385) <= 0; flappy_W(58, 386) <= 0; flappy_W(58, 387) <= 0; flappy_W(58, 388) <= 0; flappy_W(58, 389) <= 0; flappy_W(58, 390) <= 0; flappy_W(58, 391) <= 0; flappy_W(58, 392) <= 0; flappy_W(58, 393) <= 0; flappy_W(58, 394) <= 0; flappy_W(58, 395) <= 0; flappy_W(58, 396) <= 1; flappy_W(58, 397) <= 1; flappy_W(58, 398) <= 1; flappy_W(58, 399) <= 1; flappy_W(58, 400) <= 1; flappy_W(58, 401) <= 1; flappy_W(58, 402) <= 1; flappy_W(58, 403) <= 1; flappy_W(58, 404) <= 1; flappy_W(58, 405) <= 1; flappy_W(58, 406) <= 1; flappy_W(58, 407) <= 1; flappy_W(58, 408) <= 1; flappy_W(58, 409) <= 1; flappy_W(58, 410) <= 1; flappy_W(58, 411) <= 1; flappy_W(58, 412) <= 1; flappy_W(58, 413) <= 1; flappy_W(58, 414) <= 1; flappy_W(58, 415) <= 1; flappy_W(58, 416) <= 1; flappy_W(58, 417) <= 1; flappy_W(58, 418) <= 1; flappy_W(58, 419) <= 1; flappy_W(58, 420) <= 1; flappy_W(58, 421) <= 1; flappy_W(58, 422) <= 1; flappy_W(58, 423) <= 1; flappy_W(58, 424) <= 1; flappy_W(58, 425) <= 1; flappy_W(58, 426) <= 1; flappy_W(58, 427) <= 1; flappy_W(58, 428) <= 1; flappy_W(58, 429) <= 1; flappy_W(58, 430) <= 1; flappy_W(58, 431) <= 1; flappy_W(58, 432) <= 0; flappy_W(58, 433) <= 0; flappy_W(58, 434) <= 0; flappy_W(58, 435) <= 0; flappy_W(58, 436) <= 0; flappy_W(58, 437) <= 0; flappy_W(58, 438) <= 0; flappy_W(58, 439) <= 0; flappy_W(58, 440) <= 0; flappy_W(58, 441) <= 0; flappy_W(58, 442) <= 0; flappy_W(58, 443) <= 0; flappy_W(58, 444) <= 0; flappy_W(58, 445) <= 0; flappy_W(58, 446) <= 0; flappy_W(58, 447) <= 0; flappy_W(58, 448) <= 0; flappy_W(58, 449) <= 0; flappy_W(58, 450) <= 0; flappy_W(58, 451) <= 0; flappy_W(58, 452) <= 0; flappy_W(58, 453) <= 0; flappy_W(58, 454) <= 0; flappy_W(58, 455) <= 0; flappy_W(58, 456) <= 0; flappy_W(58, 457) <= 0; flappy_W(58, 458) <= 0; flappy_W(58, 459) <= 0; flappy_W(58, 460) <= 0; flappy_W(58, 461) <= 0; flappy_W(58, 462) <= 1; flappy_W(58, 463) <= 1; flappy_W(58, 464) <= 1; flappy_W(58, 465) <= 1; flappy_W(58, 466) <= 1; flappy_W(58, 467) <= 1; flappy_W(58, 468) <= 1; flappy_W(58, 469) <= 1; flappy_W(58, 470) <= 1; flappy_W(58, 471) <= 1; flappy_W(58, 472) <= 1; flappy_W(58, 473) <= 1; flappy_W(58, 474) <= 1; flappy_W(58, 475) <= 1; flappy_W(58, 476) <= 1; flappy_W(58, 477) <= 1; flappy_W(58, 478) <= 1; flappy_W(58, 479) <= 1; flappy_W(58, 480) <= 1; flappy_W(58, 481) <= 1; flappy_W(58, 482) <= 1; flappy_W(58, 483) <= 1; flappy_W(58, 484) <= 1; flappy_W(58, 485) <= 1; flappy_W(58, 486) <= 0; flappy_W(58, 487) <= 0; flappy_W(58, 488) <= 0; flappy_W(58, 489) <= 0; flappy_W(58, 490) <= 0; flappy_W(58, 491) <= 0; flappy_W(58, 492) <= 0; flappy_W(58, 493) <= 0; flappy_W(58, 494) <= 0; flappy_W(58, 495) <= 0; flappy_W(58, 496) <= 0; flappy_W(58, 497) <= 0; flappy_W(58, 498) <= 0; flappy_W(58, 499) <= 0; flappy_W(58, 500) <= 0; flappy_W(58, 501) <= 0; flappy_W(58, 502) <= 0; flappy_W(58, 503) <= 0; flappy_W(58, 504) <= 1; flappy_W(58, 505) <= 1; flappy_W(58, 506) <= 1; flappy_W(58, 507) <= 1; flappy_W(58, 508) <= 1; flappy_W(58, 509) <= 1; flappy_W(58, 510) <= 1; flappy_W(58, 511) <= 1; flappy_W(58, 512) <= 1; flappy_W(58, 513) <= 1; flappy_W(58, 514) <= 1; flappy_W(58, 515) <= 1; flappy_W(58, 516) <= 1; flappy_W(58, 517) <= 1; flappy_W(58, 518) <= 1; flappy_W(58, 519) <= 1; flappy_W(58, 520) <= 1; flappy_W(58, 521) <= 1; flappy_W(58, 522) <= 0; flappy_W(58, 523) <= 0; flappy_W(58, 524) <= 0; flappy_W(58, 525) <= 0; flappy_W(58, 526) <= 0; flappy_W(58, 527) <= 0; flappy_W(58, 528) <= 0; flappy_W(58, 529) <= 0; flappy_W(58, 530) <= 0; flappy_W(58, 531) <= 0; flappy_W(58, 532) <= 0; flappy_W(58, 533) <= 0; flappy_W(58, 534) <= 1; flappy_W(58, 535) <= 1; flappy_W(58, 536) <= 1; flappy_W(58, 537) <= 1; flappy_W(58, 538) <= 1; flappy_W(58, 539) <= 1; flappy_W(58, 540) <= 1; flappy_W(58, 541) <= 1; flappy_W(58, 542) <= 1; flappy_W(58, 543) <= 1; flappy_W(58, 544) <= 1; flappy_W(58, 545) <= 1; flappy_W(58, 546) <= 0; flappy_W(58, 547) <= 0; flappy_W(58, 548) <= 0; flappy_W(58, 549) <= 0; flappy_W(58, 550) <= 0; flappy_W(58, 551) <= 0; flappy_W(58, 552) <= 0; flappy_W(58, 553) <= 0; flappy_W(58, 554) <= 0; flappy_W(58, 555) <= 0; flappy_W(58, 556) <= 0; flappy_W(58, 557) <= 0; flappy_W(58, 558) <= 1; flappy_W(58, 559) <= 1; flappy_W(58, 560) <= 1; flappy_W(58, 561) <= 1; flappy_W(58, 562) <= 1; flappy_W(58, 563) <= 1; flappy_W(58, 564) <= 1; flappy_W(58, 565) <= 1; flappy_W(58, 566) <= 1; flappy_W(58, 567) <= 1; flappy_W(58, 568) <= 1; flappy_W(58, 569) <= 1; flappy_W(58, 570) <= 1; flappy_W(58, 571) <= 1; flappy_W(58, 572) <= 1; flappy_W(58, 573) <= 1; flappy_W(58, 574) <= 1; flappy_W(58, 575) <= 1; flappy_W(58, 576) <= 1; flappy_W(58, 577) <= 1; flappy_W(58, 578) <= 1; flappy_W(58, 579) <= 1; flappy_W(58, 580) <= 1; flappy_W(58, 581) <= 1; flappy_W(58, 582) <= 1; flappy_W(58, 583) <= 1; flappy_W(58, 584) <= 1; flappy_W(58, 585) <= 1; flappy_W(58, 586) <= 1; flappy_W(58, 587) <= 1; flappy_W(58, 588) <= 0; flappy_W(58, 589) <= 0; flappy_W(58, 590) <= 0; flappy_W(58, 591) <= 0; flappy_W(58, 592) <= 0; flappy_W(58, 593) <= 0; 
flappy_W(59, 0) <= 1; flappy_W(59, 1) <= 1; flappy_W(59, 2) <= 1; flappy_W(59, 3) <= 1; flappy_W(59, 4) <= 1; flappy_W(59, 5) <= 1; flappy_W(59, 6) <= 1; flappy_W(59, 7) <= 1; flappy_W(59, 8) <= 1; flappy_W(59, 9) <= 1; flappy_W(59, 10) <= 1; flappy_W(59, 11) <= 1; flappy_W(59, 12) <= 1; flappy_W(59, 13) <= 1; flappy_W(59, 14) <= 1; flappy_W(59, 15) <= 1; flappy_W(59, 16) <= 1; flappy_W(59, 17) <= 1; flappy_W(59, 18) <= 1; flappy_W(59, 19) <= 1; flappy_W(59, 20) <= 1; flappy_W(59, 21) <= 1; flappy_W(59, 22) <= 1; flappy_W(59, 23) <= 1; flappy_W(59, 24) <= 0; flappy_W(59, 25) <= 0; flappy_W(59, 26) <= 0; flappy_W(59, 27) <= 0; flappy_W(59, 28) <= 0; flappy_W(59, 29) <= 0; flappy_W(59, 30) <= 0; flappy_W(59, 31) <= 0; flappy_W(59, 32) <= 0; flappy_W(59, 33) <= 0; flappy_W(59, 34) <= 0; flappy_W(59, 35) <= 0; flappy_W(59, 36) <= 0; flappy_W(59, 37) <= 0; flappy_W(59, 38) <= 0; flappy_W(59, 39) <= 0; flappy_W(59, 40) <= 0; flappy_W(59, 41) <= 0; flappy_W(59, 42) <= 0; flappy_W(59, 43) <= 0; flappy_W(59, 44) <= 0; flappy_W(59, 45) <= 0; flappy_W(59, 46) <= 0; flappy_W(59, 47) <= 0; flappy_W(59, 48) <= 0; flappy_W(59, 49) <= 0; flappy_W(59, 50) <= 0; flappy_W(59, 51) <= 0; flappy_W(59, 52) <= 0; flappy_W(59, 53) <= 0; flappy_W(59, 54) <= 1; flappy_W(59, 55) <= 1; flappy_W(59, 56) <= 1; flappy_W(59, 57) <= 1; flappy_W(59, 58) <= 1; flappy_W(59, 59) <= 1; flappy_W(59, 60) <= 1; flappy_W(59, 61) <= 1; flappy_W(59, 62) <= 1; flappy_W(59, 63) <= 1; flappy_W(59, 64) <= 1; flappy_W(59, 65) <= 1; flappy_W(59, 66) <= 1; flappy_W(59, 67) <= 1; flappy_W(59, 68) <= 1; flappy_W(59, 69) <= 1; flappy_W(59, 70) <= 1; flappy_W(59, 71) <= 1; flappy_W(59, 72) <= 1; flappy_W(59, 73) <= 1; flappy_W(59, 74) <= 1; flappy_W(59, 75) <= 1; flappy_W(59, 76) <= 1; flappy_W(59, 77) <= 1; flappy_W(59, 78) <= 1; flappy_W(59, 79) <= 1; flappy_W(59, 80) <= 1; flappy_W(59, 81) <= 1; flappy_W(59, 82) <= 1; flappy_W(59, 83) <= 1; flappy_W(59, 84) <= 1; flappy_W(59, 85) <= 1; flappy_W(59, 86) <= 1; flappy_W(59, 87) <= 1; flappy_W(59, 88) <= 1; flappy_W(59, 89) <= 1; flappy_W(59, 90) <= 1; flappy_W(59, 91) <= 1; flappy_W(59, 92) <= 1; flappy_W(59, 93) <= 1; flappy_W(59, 94) <= 1; flappy_W(59, 95) <= 1; flappy_W(59, 96) <= 0; flappy_W(59, 97) <= 0; flappy_W(59, 98) <= 0; flappy_W(59, 99) <= 0; flappy_W(59, 100) <= 0; flappy_W(59, 101) <= 0; flappy_W(59, 102) <= 0; flappy_W(59, 103) <= 0; flappy_W(59, 104) <= 0; flappy_W(59, 105) <= 0; flappy_W(59, 106) <= 0; flappy_W(59, 107) <= 0; flappy_W(59, 108) <= 1; flappy_W(59, 109) <= 1; flappy_W(59, 110) <= 1; flappy_W(59, 111) <= 1; flappy_W(59, 112) <= 1; flappy_W(59, 113) <= 1; flappy_W(59, 114) <= 1; flappy_W(59, 115) <= 1; flappy_W(59, 116) <= 1; flappy_W(59, 117) <= 1; flappy_W(59, 118) <= 1; flappy_W(59, 119) <= 1; flappy_W(59, 120) <= 0; flappy_W(59, 121) <= 0; flappy_W(59, 122) <= 0; flappy_W(59, 123) <= 0; flappy_W(59, 124) <= 0; flappy_W(59, 125) <= 0; flappy_W(59, 126) <= 0; flappy_W(59, 127) <= 0; flappy_W(59, 128) <= 0; flappy_W(59, 129) <= 0; flappy_W(59, 130) <= 0; flappy_W(59, 131) <= 0; flappy_W(59, 132) <= 0; flappy_W(59, 133) <= 0; flappy_W(59, 134) <= 0; flappy_W(59, 135) <= 0; flappy_W(59, 136) <= 0; flappy_W(59, 137) <= 0; flappy_W(59, 138) <= 1; flappy_W(59, 139) <= 1; flappy_W(59, 140) <= 1; flappy_W(59, 141) <= 1; flappy_W(59, 142) <= 1; flappy_W(59, 143) <= 1; flappy_W(59, 144) <= 1; flappy_W(59, 145) <= 1; flappy_W(59, 146) <= 1; flappy_W(59, 147) <= 1; flappy_W(59, 148) <= 1; flappy_W(59, 149) <= 1; flappy_W(59, 150) <= 0; flappy_W(59, 151) <= 0; flappy_W(59, 152) <= 0; flappy_W(59, 153) <= 0; flappy_W(59, 154) <= 0; flappy_W(59, 155) <= 0; flappy_W(59, 156) <= 0; flappy_W(59, 157) <= 0; flappy_W(59, 158) <= 0; flappy_W(59, 159) <= 0; flappy_W(59, 160) <= 0; flappy_W(59, 161) <= 0; flappy_W(59, 162) <= 1; flappy_W(59, 163) <= 1; flappy_W(59, 164) <= 1; flappy_W(59, 165) <= 1; flappy_W(59, 166) <= 1; flappy_W(59, 167) <= 1; flappy_W(59, 168) <= 1; flappy_W(59, 169) <= 1; flappy_W(59, 170) <= 1; flappy_W(59, 171) <= 1; flappy_W(59, 172) <= 1; flappy_W(59, 173) <= 1; flappy_W(59, 174) <= 1; flappy_W(59, 175) <= 1; flappy_W(59, 176) <= 1; flappy_W(59, 177) <= 1; flappy_W(59, 178) <= 1; flappy_W(59, 179) <= 1; flappy_W(59, 180) <= 1; flappy_W(59, 181) <= 1; flappy_W(59, 182) <= 1; flappy_W(59, 183) <= 1; flappy_W(59, 184) <= 1; flappy_W(59, 185) <= 1; flappy_W(59, 186) <= 0; flappy_W(59, 187) <= 0; flappy_W(59, 188) <= 0; flappy_W(59, 189) <= 0; flappy_W(59, 190) <= 0; flappy_W(59, 191) <= 0; flappy_W(59, 192) <= 0; flappy_W(59, 193) <= 0; flappy_W(59, 194) <= 0; flappy_W(59, 195) <= 0; flappy_W(59, 196) <= 0; flappy_W(59, 197) <= 0; flappy_W(59, 198) <= 0; flappy_W(59, 199) <= 0; flappy_W(59, 200) <= 0; flappy_W(59, 201) <= 0; flappy_W(59, 202) <= 0; flappy_W(59, 203) <= 0; flappy_W(59, 204) <= 0; flappy_W(59, 205) <= 0; flappy_W(59, 206) <= 0; flappy_W(59, 207) <= 0; flappy_W(59, 208) <= 0; flappy_W(59, 209) <= 0; flappy_W(59, 210) <= 0; flappy_W(59, 211) <= 0; flappy_W(59, 212) <= 0; flappy_W(59, 213) <= 0; flappy_W(59, 214) <= 0; flappy_W(59, 215) <= 0; flappy_W(59, 216) <= 1; flappy_W(59, 217) <= 1; flappy_W(59, 218) <= 1; flappy_W(59, 219) <= 1; flappy_W(59, 220) <= 1; flappy_W(59, 221) <= 1; flappy_W(59, 222) <= 1; flappy_W(59, 223) <= 1; flappy_W(59, 224) <= 1; flappy_W(59, 225) <= 1; flappy_W(59, 226) <= 1; flappy_W(59, 227) <= 1; flappy_W(59, 228) <= 1; flappy_W(59, 229) <= 1; flappy_W(59, 230) <= 1; flappy_W(59, 231) <= 1; flappy_W(59, 232) <= 1; flappy_W(59, 233) <= 1; flappy_W(59, 234) <= 1; flappy_W(59, 235) <= 1; flappy_W(59, 236) <= 1; flappy_W(59, 237) <= 1; flappy_W(59, 238) <= 1; flappy_W(59, 239) <= 1; flappy_W(59, 240) <= 0; flappy_W(59, 241) <= 0; flappy_W(59, 242) <= 0; flappy_W(59, 243) <= 0; flappy_W(59, 244) <= 0; flappy_W(59, 245) <= 0; flappy_W(59, 246) <= 0; flappy_W(59, 247) <= 0; flappy_W(59, 248) <= 0; flappy_W(59, 249) <= 0; flappy_W(59, 250) <= 0; flappy_W(59, 251) <= 0; flappy_W(59, 252) <= 0; flappy_W(59, 253) <= 0; flappy_W(59, 254) <= 0; flappy_W(59, 255) <= 0; flappy_W(59, 256) <= 0; flappy_W(59, 257) <= 0; flappy_W(59, 258) <= 0; flappy_W(59, 259) <= 0; flappy_W(59, 260) <= 0; flappy_W(59, 261) <= 0; flappy_W(59, 262) <= 0; flappy_W(59, 263) <= 0; flappy_W(59, 264) <= 0; flappy_W(59, 265) <= 0; flappy_W(59, 266) <= 0; flappy_W(59, 267) <= 0; flappy_W(59, 268) <= 0; flappy_W(59, 269) <= 0; flappy_W(59, 270) <= 0; flappy_W(59, 271) <= 0; flappy_W(59, 272) <= 0; flappy_W(59, 273) <= 0; flappy_W(59, 274) <= 0; flappy_W(59, 275) <= 0; flappy_W(59, 276) <= 0; flappy_W(59, 277) <= 0; flappy_W(59, 278) <= 0; flappy_W(59, 279) <= 0; flappy_W(59, 280) <= 0; flappy_W(59, 281) <= 0; flappy_W(59, 282) <= 1; flappy_W(59, 283) <= 1; flappy_W(59, 284) <= 1; flappy_W(59, 285) <= 1; flappy_W(59, 286) <= 1; flappy_W(59, 287) <= 1; flappy_W(59, 288) <= 1; flappy_W(59, 289) <= 1; flappy_W(59, 290) <= 1; flappy_W(59, 291) <= 1; flappy_W(59, 292) <= 1; flappy_W(59, 293) <= 1; flappy_W(59, 294) <= 1; flappy_W(59, 295) <= 1; flappy_W(59, 296) <= 1; flappy_W(59, 297) <= 1; flappy_W(59, 298) <= 1; flappy_W(59, 299) <= 1; flappy_W(59, 300) <= 1; flappy_W(59, 301) <= 1; flappy_W(59, 302) <= 1; flappy_W(59, 303) <= 1; flappy_W(59, 304) <= 1; flappy_W(59, 305) <= 1; flappy_W(59, 306) <= 0; flappy_W(59, 307) <= 0; flappy_W(59, 308) <= 0; flappy_W(59, 309) <= 0; flappy_W(59, 310) <= 0; flappy_W(59, 311) <= 0; flappy_W(59, 312) <= 0; flappy_W(59, 313) <= 0; flappy_W(59, 314) <= 0; flappy_W(59, 315) <= 0; flappy_W(59, 316) <= 0; flappy_W(59, 317) <= 0; flappy_W(59, 318) <= 0; flappy_W(59, 319) <= 0; flappy_W(59, 320) <= 0; flappy_W(59, 321) <= 0; flappy_W(59, 322) <= 0; flappy_W(59, 323) <= 0; flappy_W(59, 324) <= 0; flappy_W(59, 325) <= 0; flappy_W(59, 326) <= 0; flappy_W(59, 327) <= 0; flappy_W(59, 328) <= 0; flappy_W(59, 329) <= 0; flappy_W(59, 330) <= 0; flappy_W(59, 331) <= 0; flappy_W(59, 332) <= 0; flappy_W(59, 333) <= 0; flappy_W(59, 334) <= 0; flappy_W(59, 335) <= 0; flappy_W(59, 336) <= 0; flappy_W(59, 337) <= 0; flappy_W(59, 338) <= 0; flappy_W(59, 339) <= 0; flappy_W(59, 340) <= 0; flappy_W(59, 341) <= 0; flappy_W(59, 342) <= 0; flappy_W(59, 343) <= 0; flappy_W(59, 344) <= 0; flappy_W(59, 345) <= 0; flappy_W(59, 346) <= 0; flappy_W(59, 347) <= 0; flappy_W(59, 348) <= 0; flappy_W(59, 349) <= 0; flappy_W(59, 350) <= 0; flappy_W(59, 351) <= 0; flappy_W(59, 352) <= 0; flappy_W(59, 353) <= 0; flappy_W(59, 354) <= 0; flappy_W(59, 355) <= 0; flappy_W(59, 356) <= 0; flappy_W(59, 357) <= 0; flappy_W(59, 358) <= 0; flappy_W(59, 359) <= 0; flappy_W(59, 360) <= 0; flappy_W(59, 361) <= 0; flappy_W(59, 362) <= 0; flappy_W(59, 363) <= 0; flappy_W(59, 364) <= 0; flappy_W(59, 365) <= 0; flappy_W(59, 366) <= 0; flappy_W(59, 367) <= 0; flappy_W(59, 368) <= 0; flappy_W(59, 369) <= 0; flappy_W(59, 370) <= 0; flappy_W(59, 371) <= 0; flappy_W(59, 372) <= 0; flappy_W(59, 373) <= 0; flappy_W(59, 374) <= 0; flappy_W(59, 375) <= 0; flappy_W(59, 376) <= 0; flappy_W(59, 377) <= 0; flappy_W(59, 378) <= 0; flappy_W(59, 379) <= 0; flappy_W(59, 380) <= 0; flappy_W(59, 381) <= 0; flappy_W(59, 382) <= 0; flappy_W(59, 383) <= 0; flappy_W(59, 384) <= 0; flappy_W(59, 385) <= 0; flappy_W(59, 386) <= 0; flappy_W(59, 387) <= 0; flappy_W(59, 388) <= 0; flappy_W(59, 389) <= 0; flappy_W(59, 390) <= 0; flappy_W(59, 391) <= 0; flappy_W(59, 392) <= 0; flappy_W(59, 393) <= 0; flappy_W(59, 394) <= 0; flappy_W(59, 395) <= 0; flappy_W(59, 396) <= 1; flappy_W(59, 397) <= 1; flappy_W(59, 398) <= 1; flappy_W(59, 399) <= 1; flappy_W(59, 400) <= 1; flappy_W(59, 401) <= 1; flappy_W(59, 402) <= 1; flappy_W(59, 403) <= 1; flappy_W(59, 404) <= 1; flappy_W(59, 405) <= 1; flappy_W(59, 406) <= 1; flappy_W(59, 407) <= 1; flappy_W(59, 408) <= 1; flappy_W(59, 409) <= 1; flappy_W(59, 410) <= 1; flappy_W(59, 411) <= 1; flappy_W(59, 412) <= 1; flappy_W(59, 413) <= 1; flappy_W(59, 414) <= 1; flappy_W(59, 415) <= 1; flappy_W(59, 416) <= 1; flappy_W(59, 417) <= 1; flappy_W(59, 418) <= 1; flappy_W(59, 419) <= 1; flappy_W(59, 420) <= 1; flappy_W(59, 421) <= 1; flappy_W(59, 422) <= 1; flappy_W(59, 423) <= 1; flappy_W(59, 424) <= 1; flappy_W(59, 425) <= 1; flappy_W(59, 426) <= 1; flappy_W(59, 427) <= 1; flappy_W(59, 428) <= 1; flappy_W(59, 429) <= 1; flappy_W(59, 430) <= 1; flappy_W(59, 431) <= 1; flappy_W(59, 432) <= 0; flappy_W(59, 433) <= 0; flappy_W(59, 434) <= 0; flappy_W(59, 435) <= 0; flappy_W(59, 436) <= 0; flappy_W(59, 437) <= 0; flappy_W(59, 438) <= 0; flappy_W(59, 439) <= 0; flappy_W(59, 440) <= 0; flappy_W(59, 441) <= 0; flappy_W(59, 442) <= 0; flappy_W(59, 443) <= 0; flappy_W(59, 444) <= 0; flappy_W(59, 445) <= 0; flappy_W(59, 446) <= 0; flappy_W(59, 447) <= 0; flappy_W(59, 448) <= 0; flappy_W(59, 449) <= 0; flappy_W(59, 450) <= 0; flappy_W(59, 451) <= 0; flappy_W(59, 452) <= 0; flappy_W(59, 453) <= 0; flappy_W(59, 454) <= 0; flappy_W(59, 455) <= 0; flappy_W(59, 456) <= 0; flappy_W(59, 457) <= 0; flappy_W(59, 458) <= 0; flappy_W(59, 459) <= 0; flappy_W(59, 460) <= 0; flappy_W(59, 461) <= 0; flappy_W(59, 462) <= 1; flappy_W(59, 463) <= 1; flappy_W(59, 464) <= 1; flappy_W(59, 465) <= 1; flappy_W(59, 466) <= 1; flappy_W(59, 467) <= 1; flappy_W(59, 468) <= 1; flappy_W(59, 469) <= 1; flappy_W(59, 470) <= 1; flappy_W(59, 471) <= 1; flappy_W(59, 472) <= 1; flappy_W(59, 473) <= 1; flappy_W(59, 474) <= 1; flappy_W(59, 475) <= 1; flappy_W(59, 476) <= 1; flappy_W(59, 477) <= 1; flappy_W(59, 478) <= 1; flappy_W(59, 479) <= 1; flappy_W(59, 480) <= 1; flappy_W(59, 481) <= 1; flappy_W(59, 482) <= 1; flappy_W(59, 483) <= 1; flappy_W(59, 484) <= 1; flappy_W(59, 485) <= 1; flappy_W(59, 486) <= 0; flappy_W(59, 487) <= 0; flappy_W(59, 488) <= 0; flappy_W(59, 489) <= 0; flappy_W(59, 490) <= 0; flappy_W(59, 491) <= 0; flappy_W(59, 492) <= 0; flappy_W(59, 493) <= 0; flappy_W(59, 494) <= 0; flappy_W(59, 495) <= 0; flappy_W(59, 496) <= 0; flappy_W(59, 497) <= 0; flappy_W(59, 498) <= 0; flappy_W(59, 499) <= 0; flappy_W(59, 500) <= 0; flappy_W(59, 501) <= 0; flappy_W(59, 502) <= 0; flappy_W(59, 503) <= 0; flappy_W(59, 504) <= 1; flappy_W(59, 505) <= 1; flappy_W(59, 506) <= 1; flappy_W(59, 507) <= 1; flappy_W(59, 508) <= 1; flappy_W(59, 509) <= 1; flappy_W(59, 510) <= 1; flappy_W(59, 511) <= 1; flappy_W(59, 512) <= 1; flappy_W(59, 513) <= 1; flappy_W(59, 514) <= 1; flappy_W(59, 515) <= 1; flappy_W(59, 516) <= 1; flappy_W(59, 517) <= 1; flappy_W(59, 518) <= 1; flappy_W(59, 519) <= 1; flappy_W(59, 520) <= 1; flappy_W(59, 521) <= 1; flappy_W(59, 522) <= 0; flappy_W(59, 523) <= 0; flappy_W(59, 524) <= 0; flappy_W(59, 525) <= 0; flappy_W(59, 526) <= 0; flappy_W(59, 527) <= 0; flappy_W(59, 528) <= 0; flappy_W(59, 529) <= 0; flappy_W(59, 530) <= 0; flappy_W(59, 531) <= 0; flappy_W(59, 532) <= 0; flappy_W(59, 533) <= 0; flappy_W(59, 534) <= 1; flappy_W(59, 535) <= 1; flappy_W(59, 536) <= 1; flappy_W(59, 537) <= 1; flappy_W(59, 538) <= 1; flappy_W(59, 539) <= 1; flappy_W(59, 540) <= 1; flappy_W(59, 541) <= 1; flappy_W(59, 542) <= 1; flappy_W(59, 543) <= 1; flappy_W(59, 544) <= 1; flappy_W(59, 545) <= 1; flappy_W(59, 546) <= 0; flappy_W(59, 547) <= 0; flappy_W(59, 548) <= 0; flappy_W(59, 549) <= 0; flappy_W(59, 550) <= 0; flappy_W(59, 551) <= 0; flappy_W(59, 552) <= 0; flappy_W(59, 553) <= 0; flappy_W(59, 554) <= 0; flappy_W(59, 555) <= 0; flappy_W(59, 556) <= 0; flappy_W(59, 557) <= 0; flappy_W(59, 558) <= 1; flappy_W(59, 559) <= 1; flappy_W(59, 560) <= 1; flappy_W(59, 561) <= 1; flappy_W(59, 562) <= 1; flappy_W(59, 563) <= 1; flappy_W(59, 564) <= 1; flappy_W(59, 565) <= 1; flappy_W(59, 566) <= 1; flappy_W(59, 567) <= 1; flappy_W(59, 568) <= 1; flappy_W(59, 569) <= 1; flappy_W(59, 570) <= 1; flappy_W(59, 571) <= 1; flappy_W(59, 572) <= 1; flappy_W(59, 573) <= 1; flappy_W(59, 574) <= 1; flappy_W(59, 575) <= 1; flappy_W(59, 576) <= 1; flappy_W(59, 577) <= 1; flappy_W(59, 578) <= 1; flappy_W(59, 579) <= 1; flappy_W(59, 580) <= 1; flappy_W(59, 581) <= 1; flappy_W(59, 582) <= 1; flappy_W(59, 583) <= 1; flappy_W(59, 584) <= 1; flappy_W(59, 585) <= 1; flappy_W(59, 586) <= 1; flappy_W(59, 587) <= 1; flappy_W(59, 588) <= 0; flappy_W(59, 589) <= 0; flappy_W(59, 590) <= 0; flappy_W(59, 591) <= 0; flappy_W(59, 592) <= 0; flappy_W(59, 593) <= 0; 

end Behavioral;
