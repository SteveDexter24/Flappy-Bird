library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package cloudpkg is
    type cloud_small2D is array(0 to 26, 0 to 38) of integer;
    type cloud_large2D is array(0 to 35, 0 to 51) of integer;
    type cloud_xl2D is array(0 to 53, 0 to 77) of integer;
end package;

use work.cloudpkg.all;

entity clouds is
    Port (cloud_small: out cloud_small2D; cloud_large: out cloud_large2D; cloud_xl: out cloud_xl2D);
end clouds;

architecture Behavioral of clouds is

begin

cloud_large(0, 0) <= 2; cloud_large(0, 1) <= 2; cloud_large(0, 2) <= 2; cloud_large(0, 3) <= 2; cloud_large(0, 4) <= 2; cloud_large(0, 5) <= 2; cloud_large(0, 6) <= 2; cloud_large(0, 7) <= 2; cloud_large(0, 8) <= 2; cloud_large(0, 9) <= 2; cloud_large(0, 10) <= 2; cloud_large(0, 11) <= 2; cloud_large(0, 12) <= 2; cloud_large(0, 13) <= 2; cloud_large(0, 14) <= 2; cloud_large(0, 15) <= 2; cloud_large(0, 16) <= 2; cloud_large(0, 17) <= 2; cloud_large(0, 18) <= 2; cloud_large(0, 19) <= 2; cloud_large(0, 20) <= 1; cloud_large(0, 21) <= 1; cloud_large(0, 22) <= 1; cloud_large(0, 23) <= 1; cloud_large(0, 24) <= 1; cloud_large(0, 25) <= 1; cloud_large(0, 26) <= 1; cloud_large(0, 27) <= 1; cloud_large(0, 28) <= 1; cloud_large(0, 29) <= 1; cloud_large(0, 30) <= 1; cloud_large(0, 31) <= 1; cloud_large(0, 32) <= 2; cloud_large(0, 33) <= 2; cloud_large(0, 34) <= 2; cloud_large(0, 35) <= 2; cloud_large(0, 36) <= 2; cloud_large(0, 37) <= 2; cloud_large(0, 38) <= 2; cloud_large(0, 39) <= 2; cloud_large(0, 40) <= 2; cloud_large(0, 41) <= 2; cloud_large(0, 42) <= 2; cloud_large(0, 43) <= 2; cloud_large(0, 44) <= 2; cloud_large(0, 45) <= 2; cloud_large(0, 46) <= 2; cloud_large(0, 47) <= 2; cloud_large(0, 48) <= 2; cloud_large(0, 49) <= 2; cloud_large(0, 50) <= 2; cloud_large(0, 51) <= 2; 
cloud_large(1, 0) <= 2; cloud_large(1, 1) <= 2; cloud_large(1, 2) <= 2; cloud_large(1, 3) <= 2; cloud_large(1, 4) <= 2; cloud_large(1, 5) <= 2; cloud_large(1, 6) <= 2; cloud_large(1, 7) <= 2; cloud_large(1, 8) <= 2; cloud_large(1, 9) <= 2; cloud_large(1, 10) <= 2; cloud_large(1, 11) <= 2; cloud_large(1, 12) <= 2; cloud_large(1, 13) <= 2; cloud_large(1, 14) <= 2; cloud_large(1, 15) <= 2; cloud_large(1, 16) <= 2; cloud_large(1, 17) <= 2; cloud_large(1, 18) <= 2; cloud_large(1, 19) <= 2; cloud_large(1, 20) <= 1; cloud_large(1, 21) <= 1; cloud_large(1, 22) <= 1; cloud_large(1, 23) <= 1; cloud_large(1, 24) <= 1; cloud_large(1, 25) <= 1; cloud_large(1, 26) <= 1; cloud_large(1, 27) <= 1; cloud_large(1, 28) <= 1; cloud_large(1, 29) <= 1; cloud_large(1, 30) <= 1; cloud_large(1, 31) <= 1; cloud_large(1, 32) <= 2; cloud_large(1, 33) <= 2; cloud_large(1, 34) <= 2; cloud_large(1, 35) <= 2; cloud_large(1, 36) <= 2; cloud_large(1, 37) <= 2; cloud_large(1, 38) <= 2; cloud_large(1, 39) <= 2; cloud_large(1, 40) <= 2; cloud_large(1, 41) <= 2; cloud_large(1, 42) <= 2; cloud_large(1, 43) <= 2; cloud_large(1, 44) <= 2; cloud_large(1, 45) <= 2; cloud_large(1, 46) <= 2; cloud_large(1, 47) <= 2; cloud_large(1, 48) <= 2; cloud_large(1, 49) <= 2; cloud_large(1, 50) <= 2; cloud_large(1, 51) <= 2; 
cloud_large(2, 0) <= 2; cloud_large(2, 1) <= 2; cloud_large(2, 2) <= 2; cloud_large(2, 3) <= 2; cloud_large(2, 4) <= 2; cloud_large(2, 5) <= 2; cloud_large(2, 6) <= 2; cloud_large(2, 7) <= 2; cloud_large(2, 8) <= 2; cloud_large(2, 9) <= 2; cloud_large(2, 10) <= 2; cloud_large(2, 11) <= 2; cloud_large(2, 12) <= 2; cloud_large(2, 13) <= 2; cloud_large(2, 14) <= 2; cloud_large(2, 15) <= 2; cloud_large(2, 16) <= 2; cloud_large(2, 17) <= 2; cloud_large(2, 18) <= 2; cloud_large(2, 19) <= 2; cloud_large(2, 20) <= 1; cloud_large(2, 21) <= 1; cloud_large(2, 22) <= 1; cloud_large(2, 23) <= 1; cloud_large(2, 24) <= 1; cloud_large(2, 25) <= 1; cloud_large(2, 26) <= 1; cloud_large(2, 27) <= 1; cloud_large(2, 28) <= 1; cloud_large(2, 29) <= 1; cloud_large(2, 30) <= 1; cloud_large(2, 31) <= 1; cloud_large(2, 32) <= 2; cloud_large(2, 33) <= 2; cloud_large(2, 34) <= 2; cloud_large(2, 35) <= 2; cloud_large(2, 36) <= 2; cloud_large(2, 37) <= 2; cloud_large(2, 38) <= 2; cloud_large(2, 39) <= 2; cloud_large(2, 40) <= 2; cloud_large(2, 41) <= 2; cloud_large(2, 42) <= 2; cloud_large(2, 43) <= 2; cloud_large(2, 44) <= 2; cloud_large(2, 45) <= 2; cloud_large(2, 46) <= 2; cloud_large(2, 47) <= 2; cloud_large(2, 48) <= 2; cloud_large(2, 49) <= 2; cloud_large(2, 50) <= 2; cloud_large(2, 51) <= 2; 
cloud_large(3, 0) <= 2; cloud_large(3, 1) <= 2; cloud_large(3, 2) <= 2; cloud_large(3, 3) <= 2; cloud_large(3, 4) <= 2; cloud_large(3, 5) <= 2; cloud_large(3, 6) <= 2; cloud_large(3, 7) <= 2; cloud_large(3, 8) <= 2; cloud_large(3, 9) <= 2; cloud_large(3, 10) <= 2; cloud_large(3, 11) <= 2; cloud_large(3, 12) <= 2; cloud_large(3, 13) <= 2; cloud_large(3, 14) <= 2; cloud_large(3, 15) <= 2; cloud_large(3, 16) <= 2; cloud_large(3, 17) <= 2; cloud_large(3, 18) <= 2; cloud_large(3, 19) <= 2; cloud_large(3, 20) <= 1; cloud_large(3, 21) <= 1; cloud_large(3, 22) <= 1; cloud_large(3, 23) <= 1; cloud_large(3, 24) <= 1; cloud_large(3, 25) <= 1; cloud_large(3, 26) <= 1; cloud_large(3, 27) <= 1; cloud_large(3, 28) <= 1; cloud_large(3, 29) <= 1; cloud_large(3, 30) <= 1; cloud_large(3, 31) <= 1; cloud_large(3, 32) <= 2; cloud_large(3, 33) <= 2; cloud_large(3, 34) <= 2; cloud_large(3, 35) <= 2; cloud_large(3, 36) <= 2; cloud_large(3, 37) <= 2; cloud_large(3, 38) <= 2; cloud_large(3, 39) <= 2; cloud_large(3, 40) <= 2; cloud_large(3, 41) <= 2; cloud_large(3, 42) <= 2; cloud_large(3, 43) <= 2; cloud_large(3, 44) <= 2; cloud_large(3, 45) <= 2; cloud_large(3, 46) <= 2; cloud_large(3, 47) <= 2; cloud_large(3, 48) <= 2; cloud_large(3, 49) <= 2; cloud_large(3, 50) <= 2; cloud_large(3, 51) <= 2; 
cloud_large(4, 0) <= 2; cloud_large(4, 1) <= 2; cloud_large(4, 2) <= 2; cloud_large(4, 3) <= 2; cloud_large(4, 4) <= 2; cloud_large(4, 5) <= 2; cloud_large(4, 6) <= 2; cloud_large(4, 7) <= 2; cloud_large(4, 8) <= 2; cloud_large(4, 9) <= 2; cloud_large(4, 10) <= 2; cloud_large(4, 11) <= 2; cloud_large(4, 12) <= 2; cloud_large(4, 13) <= 2; cloud_large(4, 14) <= 2; cloud_large(4, 15) <= 2; cloud_large(4, 16) <= 1; cloud_large(4, 17) <= 1; cloud_large(4, 18) <= 1; cloud_large(4, 19) <= 1; cloud_large(4, 20) <= 0; cloud_large(4, 21) <= 0; cloud_large(4, 22) <= 0; cloud_large(4, 23) <= 0; cloud_large(4, 24) <= 0; cloud_large(4, 25) <= 0; cloud_large(4, 26) <= 0; cloud_large(4, 27) <= 0; cloud_large(4, 28) <= 0; cloud_large(4, 29) <= 0; cloud_large(4, 30) <= 0; cloud_large(4, 31) <= 0; cloud_large(4, 32) <= 1; cloud_large(4, 33) <= 1; cloud_large(4, 34) <= 1; cloud_large(4, 35) <= 1; cloud_large(4, 36) <= 2; cloud_large(4, 37) <= 2; cloud_large(4, 38) <= 2; cloud_large(4, 39) <= 2; cloud_large(4, 40) <= 2; cloud_large(4, 41) <= 2; cloud_large(4, 42) <= 2; cloud_large(4, 43) <= 2; cloud_large(4, 44) <= 2; cloud_large(4, 45) <= 2; cloud_large(4, 46) <= 2; cloud_large(4, 47) <= 2; cloud_large(4, 48) <= 2; cloud_large(4, 49) <= 2; cloud_large(4, 50) <= 2; cloud_large(4, 51) <= 2; 
cloud_large(5, 0) <= 2; cloud_large(5, 1) <= 2; cloud_large(5, 2) <= 2; cloud_large(5, 3) <= 2; cloud_large(5, 4) <= 2; cloud_large(5, 5) <= 2; cloud_large(5, 6) <= 2; cloud_large(5, 7) <= 2; cloud_large(5, 8) <= 2; cloud_large(5, 9) <= 2; cloud_large(5, 10) <= 2; cloud_large(5, 11) <= 2; cloud_large(5, 12) <= 2; cloud_large(5, 13) <= 2; cloud_large(5, 14) <= 2; cloud_large(5, 15) <= 2; cloud_large(5, 16) <= 1; cloud_large(5, 17) <= 1; cloud_large(5, 18) <= 1; cloud_large(5, 19) <= 1; cloud_large(5, 20) <= 0; cloud_large(5, 21) <= 0; cloud_large(5, 22) <= 0; cloud_large(5, 23) <= 0; cloud_large(5, 24) <= 0; cloud_large(5, 25) <= 0; cloud_large(5, 26) <= 0; cloud_large(5, 27) <= 0; cloud_large(5, 28) <= 0; cloud_large(5, 29) <= 0; cloud_large(5, 30) <= 0; cloud_large(5, 31) <= 0; cloud_large(5, 32) <= 1; cloud_large(5, 33) <= 1; cloud_large(5, 34) <= 1; cloud_large(5, 35) <= 1; cloud_large(5, 36) <= 2; cloud_large(5, 37) <= 2; cloud_large(5, 38) <= 2; cloud_large(5, 39) <= 2; cloud_large(5, 40) <= 2; cloud_large(5, 41) <= 2; cloud_large(5, 42) <= 2; cloud_large(5, 43) <= 2; cloud_large(5, 44) <= 2; cloud_large(5, 45) <= 2; cloud_large(5, 46) <= 2; cloud_large(5, 47) <= 2; cloud_large(5, 48) <= 2; cloud_large(5, 49) <= 2; cloud_large(5, 50) <= 2; cloud_large(5, 51) <= 2; 
cloud_large(6, 0) <= 2; cloud_large(6, 1) <= 2; cloud_large(6, 2) <= 2; cloud_large(6, 3) <= 2; cloud_large(6, 4) <= 2; cloud_large(6, 5) <= 2; cloud_large(6, 6) <= 2; cloud_large(6, 7) <= 2; cloud_large(6, 8) <= 2; cloud_large(6, 9) <= 2; cloud_large(6, 10) <= 2; cloud_large(6, 11) <= 2; cloud_large(6, 12) <= 2; cloud_large(6, 13) <= 2; cloud_large(6, 14) <= 2; cloud_large(6, 15) <= 2; cloud_large(6, 16) <= 1; cloud_large(6, 17) <= 1; cloud_large(6, 18) <= 1; cloud_large(6, 19) <= 1; cloud_large(6, 20) <= 0; cloud_large(6, 21) <= 0; cloud_large(6, 22) <= 0; cloud_large(6, 23) <= 0; cloud_large(6, 24) <= 0; cloud_large(6, 25) <= 0; cloud_large(6, 26) <= 0; cloud_large(6, 27) <= 0; cloud_large(6, 28) <= 0; cloud_large(6, 29) <= 0; cloud_large(6, 30) <= 0; cloud_large(6, 31) <= 0; cloud_large(6, 32) <= 1; cloud_large(6, 33) <= 1; cloud_large(6, 34) <= 1; cloud_large(6, 35) <= 1; cloud_large(6, 36) <= 2; cloud_large(6, 37) <= 2; cloud_large(6, 38) <= 2; cloud_large(6, 39) <= 2; cloud_large(6, 40) <= 2; cloud_large(6, 41) <= 2; cloud_large(6, 42) <= 2; cloud_large(6, 43) <= 2; cloud_large(6, 44) <= 2; cloud_large(6, 45) <= 2; cloud_large(6, 46) <= 2; cloud_large(6, 47) <= 2; cloud_large(6, 48) <= 2; cloud_large(6, 49) <= 2; cloud_large(6, 50) <= 2; cloud_large(6, 51) <= 2; 
cloud_large(7, 0) <= 2; cloud_large(7, 1) <= 2; cloud_large(7, 2) <= 2; cloud_large(7, 3) <= 2; cloud_large(7, 4) <= 2; cloud_large(7, 5) <= 2; cloud_large(7, 6) <= 2; cloud_large(7, 7) <= 2; cloud_large(7, 8) <= 2; cloud_large(7, 9) <= 2; cloud_large(7, 10) <= 2; cloud_large(7, 11) <= 2; cloud_large(7, 12) <= 2; cloud_large(7, 13) <= 2; cloud_large(7, 14) <= 2; cloud_large(7, 15) <= 2; cloud_large(7, 16) <= 1; cloud_large(7, 17) <= 1; cloud_large(7, 18) <= 1; cloud_large(7, 19) <= 1; cloud_large(7, 20) <= 0; cloud_large(7, 21) <= 0; cloud_large(7, 22) <= 0; cloud_large(7, 23) <= 0; cloud_large(7, 24) <= 0; cloud_large(7, 25) <= 0; cloud_large(7, 26) <= 0; cloud_large(7, 27) <= 0; cloud_large(7, 28) <= 0; cloud_large(7, 29) <= 0; cloud_large(7, 30) <= 0; cloud_large(7, 31) <= 0; cloud_large(7, 32) <= 1; cloud_large(7, 33) <= 1; cloud_large(7, 34) <= 1; cloud_large(7, 35) <= 1; cloud_large(7, 36) <= 2; cloud_large(7, 37) <= 2; cloud_large(7, 38) <= 2; cloud_large(7, 39) <= 2; cloud_large(7, 40) <= 2; cloud_large(7, 41) <= 2; cloud_large(7, 42) <= 2; cloud_large(7, 43) <= 2; cloud_large(7, 44) <= 2; cloud_large(7, 45) <= 2; cloud_large(7, 46) <= 2; cloud_large(7, 47) <= 2; cloud_large(7, 48) <= 2; cloud_large(7, 49) <= 2; cloud_large(7, 50) <= 2; cloud_large(7, 51) <= 2; 
cloud_large(8, 0) <= 2; cloud_large(8, 1) <= 2; cloud_large(8, 2) <= 2; cloud_large(8, 3) <= 2; cloud_large(8, 4) <= 2; cloud_large(8, 5) <= 2; cloud_large(8, 6) <= 2; cloud_large(8, 7) <= 2; cloud_large(8, 8) <= 1; cloud_large(8, 9) <= 1; cloud_large(8, 10) <= 1; cloud_large(8, 11) <= 1; cloud_large(8, 12) <= 1; cloud_large(8, 13) <= 1; cloud_large(8, 14) <= 1; cloud_large(8, 15) <= 1; cloud_large(8, 16) <= 0; cloud_large(8, 17) <= 0; cloud_large(8, 18) <= 0; cloud_large(8, 19) <= 0; cloud_large(8, 20) <= 0; cloud_large(8, 21) <= 0; cloud_large(8, 22) <= 0; cloud_large(8, 23) <= 0; cloud_large(8, 24) <= 0; cloud_large(8, 25) <= 0; cloud_large(8, 26) <= 0; cloud_large(8, 27) <= 0; cloud_large(8, 28) <= 0; cloud_large(8, 29) <= 0; cloud_large(8, 30) <= 0; cloud_large(8, 31) <= 0; cloud_large(8, 32) <= 0; cloud_large(8, 33) <= 0; cloud_large(8, 34) <= 0; cloud_large(8, 35) <= 0; cloud_large(8, 36) <= 1; cloud_large(8, 37) <= 1; cloud_large(8, 38) <= 1; cloud_large(8, 39) <= 1; cloud_large(8, 40) <= 2; cloud_large(8, 41) <= 2; cloud_large(8, 42) <= 2; cloud_large(8, 43) <= 2; cloud_large(8, 44) <= 2; cloud_large(8, 45) <= 2; cloud_large(8, 46) <= 2; cloud_large(8, 47) <= 2; cloud_large(8, 48) <= 2; cloud_large(8, 49) <= 2; cloud_large(8, 50) <= 2; cloud_large(8, 51) <= 2; 
cloud_large(9, 0) <= 2; cloud_large(9, 1) <= 2; cloud_large(9, 2) <= 2; cloud_large(9, 3) <= 2; cloud_large(9, 4) <= 2; cloud_large(9, 5) <= 2; cloud_large(9, 6) <= 2; cloud_large(9, 7) <= 2; cloud_large(9, 8) <= 1; cloud_large(9, 9) <= 1; cloud_large(9, 10) <= 1; cloud_large(9, 11) <= 1; cloud_large(9, 12) <= 1; cloud_large(9, 13) <= 1; cloud_large(9, 14) <= 1; cloud_large(9, 15) <= 1; cloud_large(9, 16) <= 0; cloud_large(9, 17) <= 0; cloud_large(9, 18) <= 0; cloud_large(9, 19) <= 0; cloud_large(9, 20) <= 0; cloud_large(9, 21) <= 0; cloud_large(9, 22) <= 0; cloud_large(9, 23) <= 0; cloud_large(9, 24) <= 0; cloud_large(9, 25) <= 0; cloud_large(9, 26) <= 0; cloud_large(9, 27) <= 0; cloud_large(9, 28) <= 0; cloud_large(9, 29) <= 0; cloud_large(9, 30) <= 0; cloud_large(9, 31) <= 0; cloud_large(9, 32) <= 0; cloud_large(9, 33) <= 0; cloud_large(9, 34) <= 0; cloud_large(9, 35) <= 0; cloud_large(9, 36) <= 1; cloud_large(9, 37) <= 1; cloud_large(9, 38) <= 1; cloud_large(9, 39) <= 1; cloud_large(9, 40) <= 2; cloud_large(9, 41) <= 2; cloud_large(9, 42) <= 2; cloud_large(9, 43) <= 2; cloud_large(9, 44) <= 2; cloud_large(9, 45) <= 2; cloud_large(9, 46) <= 2; cloud_large(9, 47) <= 2; cloud_large(9, 48) <= 2; cloud_large(9, 49) <= 2; cloud_large(9, 50) <= 2; cloud_large(9, 51) <= 2; 
cloud_large(10, 0) <= 2; cloud_large(10, 1) <= 2; cloud_large(10, 2) <= 2; cloud_large(10, 3) <= 2; cloud_large(10, 4) <= 2; cloud_large(10, 5) <= 2; cloud_large(10, 6) <= 2; cloud_large(10, 7) <= 2; cloud_large(10, 8) <= 1; cloud_large(10, 9) <= 1; cloud_large(10, 10) <= 1; cloud_large(10, 11) <= 1; cloud_large(10, 12) <= 1; cloud_large(10, 13) <= 1; cloud_large(10, 14) <= 1; cloud_large(10, 15) <= 1; cloud_large(10, 16) <= 0; cloud_large(10, 17) <= 0; cloud_large(10, 18) <= 0; cloud_large(10, 19) <= 0; cloud_large(10, 20) <= 0; cloud_large(10, 21) <= 0; cloud_large(10, 22) <= 0; cloud_large(10, 23) <= 0; cloud_large(10, 24) <= 0; cloud_large(10, 25) <= 0; cloud_large(10, 26) <= 0; cloud_large(10, 27) <= 0; cloud_large(10, 28) <= 0; cloud_large(10, 29) <= 0; cloud_large(10, 30) <= 0; cloud_large(10, 31) <= 0; cloud_large(10, 32) <= 0; cloud_large(10, 33) <= 0; cloud_large(10, 34) <= 0; cloud_large(10, 35) <= 0; cloud_large(10, 36) <= 1; cloud_large(10, 37) <= 1; cloud_large(10, 38) <= 1; cloud_large(10, 39) <= 1; cloud_large(10, 40) <= 2; cloud_large(10, 41) <= 2; cloud_large(10, 42) <= 2; cloud_large(10, 43) <= 2; cloud_large(10, 44) <= 2; cloud_large(10, 45) <= 2; cloud_large(10, 46) <= 2; cloud_large(10, 47) <= 2; cloud_large(10, 48) <= 2; cloud_large(10, 49) <= 2; cloud_large(10, 50) <= 2; cloud_large(10, 51) <= 2; 
cloud_large(11, 0) <= 2; cloud_large(11, 1) <= 2; cloud_large(11, 2) <= 2; cloud_large(11, 3) <= 2; cloud_large(11, 4) <= 2; cloud_large(11, 5) <= 2; cloud_large(11, 6) <= 2; cloud_large(11, 7) <= 2; cloud_large(11, 8) <= 1; cloud_large(11, 9) <= 1; cloud_large(11, 10) <= 1; cloud_large(11, 11) <= 1; cloud_large(11, 12) <= 1; cloud_large(11, 13) <= 1; cloud_large(11, 14) <= 1; cloud_large(11, 15) <= 1; cloud_large(11, 16) <= 0; cloud_large(11, 17) <= 0; cloud_large(11, 18) <= 0; cloud_large(11, 19) <= 0; cloud_large(11, 20) <= 0; cloud_large(11, 21) <= 0; cloud_large(11, 22) <= 0; cloud_large(11, 23) <= 0; cloud_large(11, 24) <= 0; cloud_large(11, 25) <= 0; cloud_large(11, 26) <= 0; cloud_large(11, 27) <= 0; cloud_large(11, 28) <= 0; cloud_large(11, 29) <= 0; cloud_large(11, 30) <= 0; cloud_large(11, 31) <= 0; cloud_large(11, 32) <= 0; cloud_large(11, 33) <= 0; cloud_large(11, 34) <= 0; cloud_large(11, 35) <= 0; cloud_large(11, 36) <= 1; cloud_large(11, 37) <= 1; cloud_large(11, 38) <= 1; cloud_large(11, 39) <= 1; cloud_large(11, 40) <= 2; cloud_large(11, 41) <= 2; cloud_large(11, 42) <= 2; cloud_large(11, 43) <= 2; cloud_large(11, 44) <= 2; cloud_large(11, 45) <= 2; cloud_large(11, 46) <= 2; cloud_large(11, 47) <= 2; cloud_large(11, 48) <= 2; cloud_large(11, 49) <= 2; cloud_large(11, 50) <= 2; cloud_large(11, 51) <= 2; 
cloud_large(12, 0) <= 2; cloud_large(12, 1) <= 2; cloud_large(12, 2) <= 2; cloud_large(12, 3) <= 2; cloud_large(12, 4) <= 1; cloud_large(12, 5) <= 1; cloud_large(12, 6) <= 1; cloud_large(12, 7) <= 1; cloud_large(12, 8) <= 0; cloud_large(12, 9) <= 0; cloud_large(12, 10) <= 0; cloud_large(12, 11) <= 0; cloud_large(12, 12) <= 0; cloud_large(12, 13) <= 0; cloud_large(12, 14) <= 0; cloud_large(12, 15) <= 0; cloud_large(12, 16) <= 0; cloud_large(12, 17) <= 0; cloud_large(12, 18) <= 0; cloud_large(12, 19) <= 0; cloud_large(12, 20) <= 0; cloud_large(12, 21) <= 0; cloud_large(12, 22) <= 0; cloud_large(12, 23) <= 0; cloud_large(12, 24) <= 0; cloud_large(12, 25) <= 0; cloud_large(12, 26) <= 0; cloud_large(12, 27) <= 0; cloud_large(12, 28) <= 0; cloud_large(12, 29) <= 0; cloud_large(12, 30) <= 0; cloud_large(12, 31) <= 0; cloud_large(12, 32) <= 0; cloud_large(12, 33) <= 0; cloud_large(12, 34) <= 0; cloud_large(12, 35) <= 0; cloud_large(12, 36) <= 0; cloud_large(12, 37) <= 0; cloud_large(12, 38) <= 0; cloud_large(12, 39) <= 0; cloud_large(12, 40) <= 1; cloud_large(12, 41) <= 1; cloud_large(12, 42) <= 1; cloud_large(12, 43) <= 1; cloud_large(12, 44) <= 1; cloud_large(12, 45) <= 1; cloud_large(12, 46) <= 1; cloud_large(12, 47) <= 1; cloud_large(12, 48) <= 2; cloud_large(12, 49) <= 2; cloud_large(12, 50) <= 2; cloud_large(12, 51) <= 2; 
cloud_large(13, 0) <= 2; cloud_large(13, 1) <= 2; cloud_large(13, 2) <= 2; cloud_large(13, 3) <= 2; cloud_large(13, 4) <= 1; cloud_large(13, 5) <= 1; cloud_large(13, 6) <= 1; cloud_large(13, 7) <= 1; cloud_large(13, 8) <= 0; cloud_large(13, 9) <= 0; cloud_large(13, 10) <= 0; cloud_large(13, 11) <= 0; cloud_large(13, 12) <= 0; cloud_large(13, 13) <= 0; cloud_large(13, 14) <= 0; cloud_large(13, 15) <= 0; cloud_large(13, 16) <= 0; cloud_large(13, 17) <= 0; cloud_large(13, 18) <= 0; cloud_large(13, 19) <= 0; cloud_large(13, 20) <= 0; cloud_large(13, 21) <= 0; cloud_large(13, 22) <= 0; cloud_large(13, 23) <= 0; cloud_large(13, 24) <= 0; cloud_large(13, 25) <= 0; cloud_large(13, 26) <= 0; cloud_large(13, 27) <= 0; cloud_large(13, 28) <= 0; cloud_large(13, 29) <= 0; cloud_large(13, 30) <= 0; cloud_large(13, 31) <= 0; cloud_large(13, 32) <= 0; cloud_large(13, 33) <= 0; cloud_large(13, 34) <= 0; cloud_large(13, 35) <= 0; cloud_large(13, 36) <= 0; cloud_large(13, 37) <= 0; cloud_large(13, 38) <= 0; cloud_large(13, 39) <= 0; cloud_large(13, 40) <= 1; cloud_large(13, 41) <= 1; cloud_large(13, 42) <= 1; cloud_large(13, 43) <= 1; cloud_large(13, 44) <= 1; cloud_large(13, 45) <= 1; cloud_large(13, 46) <= 1; cloud_large(13, 47) <= 1; cloud_large(13, 48) <= 2; cloud_large(13, 49) <= 2; cloud_large(13, 50) <= 2; cloud_large(13, 51) <= 2; 
cloud_large(14, 0) <= 2; cloud_large(14, 1) <= 2; cloud_large(14, 2) <= 2; cloud_large(14, 3) <= 2; cloud_large(14, 4) <= 1; cloud_large(14, 5) <= 1; cloud_large(14, 6) <= 1; cloud_large(14, 7) <= 1; cloud_large(14, 8) <= 0; cloud_large(14, 9) <= 0; cloud_large(14, 10) <= 0; cloud_large(14, 11) <= 0; cloud_large(14, 12) <= 0; cloud_large(14, 13) <= 0; cloud_large(14, 14) <= 0; cloud_large(14, 15) <= 0; cloud_large(14, 16) <= 0; cloud_large(14, 17) <= 0; cloud_large(14, 18) <= 0; cloud_large(14, 19) <= 0; cloud_large(14, 20) <= 0; cloud_large(14, 21) <= 0; cloud_large(14, 22) <= 0; cloud_large(14, 23) <= 0; cloud_large(14, 24) <= 0; cloud_large(14, 25) <= 0; cloud_large(14, 26) <= 0; cloud_large(14, 27) <= 0; cloud_large(14, 28) <= 0; cloud_large(14, 29) <= 0; cloud_large(14, 30) <= 0; cloud_large(14, 31) <= 0; cloud_large(14, 32) <= 0; cloud_large(14, 33) <= 0; cloud_large(14, 34) <= 0; cloud_large(14, 35) <= 0; cloud_large(14, 36) <= 0; cloud_large(14, 37) <= 0; cloud_large(14, 38) <= 0; cloud_large(14, 39) <= 0; cloud_large(14, 40) <= 1; cloud_large(14, 41) <= 1; cloud_large(14, 42) <= 1; cloud_large(14, 43) <= 1; cloud_large(14, 44) <= 1; cloud_large(14, 45) <= 1; cloud_large(14, 46) <= 1; cloud_large(14, 47) <= 1; cloud_large(14, 48) <= 2; cloud_large(14, 49) <= 2; cloud_large(14, 50) <= 2; cloud_large(14, 51) <= 2; 
cloud_large(15, 0) <= 2; cloud_large(15, 1) <= 2; cloud_large(15, 2) <= 2; cloud_large(15, 3) <= 2; cloud_large(15, 4) <= 1; cloud_large(15, 5) <= 1; cloud_large(15, 6) <= 1; cloud_large(15, 7) <= 1; cloud_large(15, 8) <= 0; cloud_large(15, 9) <= 0; cloud_large(15, 10) <= 0; cloud_large(15, 11) <= 0; cloud_large(15, 12) <= 0; cloud_large(15, 13) <= 0; cloud_large(15, 14) <= 0; cloud_large(15, 15) <= 0; cloud_large(15, 16) <= 0; cloud_large(15, 17) <= 0; cloud_large(15, 18) <= 0; cloud_large(15, 19) <= 0; cloud_large(15, 20) <= 0; cloud_large(15, 21) <= 0; cloud_large(15, 22) <= 0; cloud_large(15, 23) <= 0; cloud_large(15, 24) <= 0; cloud_large(15, 25) <= 0; cloud_large(15, 26) <= 0; cloud_large(15, 27) <= 0; cloud_large(15, 28) <= 0; cloud_large(15, 29) <= 0; cloud_large(15, 30) <= 0; cloud_large(15, 31) <= 0; cloud_large(15, 32) <= 0; cloud_large(15, 33) <= 0; cloud_large(15, 34) <= 0; cloud_large(15, 35) <= 0; cloud_large(15, 36) <= 0; cloud_large(15, 37) <= 0; cloud_large(15, 38) <= 0; cloud_large(15, 39) <= 0; cloud_large(15, 40) <= 1; cloud_large(15, 41) <= 1; cloud_large(15, 42) <= 1; cloud_large(15, 43) <= 1; cloud_large(15, 44) <= 1; cloud_large(15, 45) <= 1; cloud_large(15, 46) <= 1; cloud_large(15, 47) <= 1; cloud_large(15, 48) <= 2; cloud_large(15, 49) <= 2; cloud_large(15, 50) <= 2; cloud_large(15, 51) <= 2; 
cloud_large(16, 0) <= 1; cloud_large(16, 1) <= 1; cloud_large(16, 2) <= 1; cloud_large(16, 3) <= 1; cloud_large(16, 4) <= 0; cloud_large(16, 5) <= 0; cloud_large(16, 6) <= 0; cloud_large(16, 7) <= 0; cloud_large(16, 8) <= 0; cloud_large(16, 9) <= 0; cloud_large(16, 10) <= 0; cloud_large(16, 11) <= 0; cloud_large(16, 12) <= 0; cloud_large(16, 13) <= 0; cloud_large(16, 14) <= 0; cloud_large(16, 15) <= 0; cloud_large(16, 16) <= 0; cloud_large(16, 17) <= 0; cloud_large(16, 18) <= 0; cloud_large(16, 19) <= 0; cloud_large(16, 20) <= 0; cloud_large(16, 21) <= 0; cloud_large(16, 22) <= 0; cloud_large(16, 23) <= 0; cloud_large(16, 24) <= 0; cloud_large(16, 25) <= 0; cloud_large(16, 26) <= 0; cloud_large(16, 27) <= 0; cloud_large(16, 28) <= 0; cloud_large(16, 29) <= 0; cloud_large(16, 30) <= 0; cloud_large(16, 31) <= 0; cloud_large(16, 32) <= 0; cloud_large(16, 33) <= 0; cloud_large(16, 34) <= 0; cloud_large(16, 35) <= 0; cloud_large(16, 36) <= 0; cloud_large(16, 37) <= 0; cloud_large(16, 38) <= 0; cloud_large(16, 39) <= 0; cloud_large(16, 40) <= 0; cloud_large(16, 41) <= 0; cloud_large(16, 42) <= 0; cloud_large(16, 43) <= 0; cloud_large(16, 44) <= 0; cloud_large(16, 45) <= 0; cloud_large(16, 46) <= 0; cloud_large(16, 47) <= 0; cloud_large(16, 48) <= 1; cloud_large(16, 49) <= 1; cloud_large(16, 50) <= 1; cloud_large(16, 51) <= 1; 
cloud_large(17, 0) <= 1; cloud_large(17, 1) <= 1; cloud_large(17, 2) <= 1; cloud_large(17, 3) <= 1; cloud_large(17, 4) <= 0; cloud_large(17, 5) <= 0; cloud_large(17, 6) <= 0; cloud_large(17, 7) <= 0; cloud_large(17, 8) <= 0; cloud_large(17, 9) <= 0; cloud_large(17, 10) <= 0; cloud_large(17, 11) <= 0; cloud_large(17, 12) <= 0; cloud_large(17, 13) <= 0; cloud_large(17, 14) <= 0; cloud_large(17, 15) <= 0; cloud_large(17, 16) <= 0; cloud_large(17, 17) <= 0; cloud_large(17, 18) <= 0; cloud_large(17, 19) <= 0; cloud_large(17, 20) <= 0; cloud_large(17, 21) <= 0; cloud_large(17, 22) <= 0; cloud_large(17, 23) <= 0; cloud_large(17, 24) <= 0; cloud_large(17, 25) <= 0; cloud_large(17, 26) <= 0; cloud_large(17, 27) <= 0; cloud_large(17, 28) <= 0; cloud_large(17, 29) <= 0; cloud_large(17, 30) <= 0; cloud_large(17, 31) <= 0; cloud_large(17, 32) <= 0; cloud_large(17, 33) <= 0; cloud_large(17, 34) <= 0; cloud_large(17, 35) <= 0; cloud_large(17, 36) <= 0; cloud_large(17, 37) <= 0; cloud_large(17, 38) <= 0; cloud_large(17, 39) <= 0; cloud_large(17, 40) <= 0; cloud_large(17, 41) <= 0; cloud_large(17, 42) <= 0; cloud_large(17, 43) <= 0; cloud_large(17, 44) <= 0; cloud_large(17, 45) <= 0; cloud_large(17, 46) <= 0; cloud_large(17, 47) <= 0; cloud_large(17, 48) <= 1; cloud_large(17, 49) <= 1; cloud_large(17, 50) <= 1; cloud_large(17, 51) <= 1; 
cloud_large(18, 0) <= 1; cloud_large(18, 1) <= 1; cloud_large(18, 2) <= 1; cloud_large(18, 3) <= 1; cloud_large(18, 4) <= 0; cloud_large(18, 5) <= 0; cloud_large(18, 6) <= 0; cloud_large(18, 7) <= 0; cloud_large(18, 8) <= 0; cloud_large(18, 9) <= 0; cloud_large(18, 10) <= 0; cloud_large(18, 11) <= 0; cloud_large(18, 12) <= 0; cloud_large(18, 13) <= 0; cloud_large(18, 14) <= 0; cloud_large(18, 15) <= 0; cloud_large(18, 16) <= 0; cloud_large(18, 17) <= 0; cloud_large(18, 18) <= 0; cloud_large(18, 19) <= 0; cloud_large(18, 20) <= 0; cloud_large(18, 21) <= 0; cloud_large(18, 22) <= 0; cloud_large(18, 23) <= 0; cloud_large(18, 24) <= 0; cloud_large(18, 25) <= 0; cloud_large(18, 26) <= 0; cloud_large(18, 27) <= 0; cloud_large(18, 28) <= 0; cloud_large(18, 29) <= 0; cloud_large(18, 30) <= 0; cloud_large(18, 31) <= 0; cloud_large(18, 32) <= 0; cloud_large(18, 33) <= 0; cloud_large(18, 34) <= 0; cloud_large(18, 35) <= 0; cloud_large(18, 36) <= 0; cloud_large(18, 37) <= 0; cloud_large(18, 38) <= 0; cloud_large(18, 39) <= 0; cloud_large(18, 40) <= 0; cloud_large(18, 41) <= 0; cloud_large(18, 42) <= 0; cloud_large(18, 43) <= 0; cloud_large(18, 44) <= 0; cloud_large(18, 45) <= 0; cloud_large(18, 46) <= 0; cloud_large(18, 47) <= 0; cloud_large(18, 48) <= 1; cloud_large(18, 49) <= 1; cloud_large(18, 50) <= 1; cloud_large(18, 51) <= 1; 
cloud_large(19, 0) <= 1; cloud_large(19, 1) <= 1; cloud_large(19, 2) <= 1; cloud_large(19, 3) <= 1; cloud_large(19, 4) <= 0; cloud_large(19, 5) <= 0; cloud_large(19, 6) <= 0; cloud_large(19, 7) <= 0; cloud_large(19, 8) <= 0; cloud_large(19, 9) <= 0; cloud_large(19, 10) <= 0; cloud_large(19, 11) <= 0; cloud_large(19, 12) <= 0; cloud_large(19, 13) <= 0; cloud_large(19, 14) <= 0; cloud_large(19, 15) <= 0; cloud_large(19, 16) <= 0; cloud_large(19, 17) <= 0; cloud_large(19, 18) <= 0; cloud_large(19, 19) <= 0; cloud_large(19, 20) <= 0; cloud_large(19, 21) <= 0; cloud_large(19, 22) <= 0; cloud_large(19, 23) <= 0; cloud_large(19, 24) <= 0; cloud_large(19, 25) <= 0; cloud_large(19, 26) <= 0; cloud_large(19, 27) <= 0; cloud_large(19, 28) <= 0; cloud_large(19, 29) <= 0; cloud_large(19, 30) <= 0; cloud_large(19, 31) <= 0; cloud_large(19, 32) <= 0; cloud_large(19, 33) <= 0; cloud_large(19, 34) <= 0; cloud_large(19, 35) <= 0; cloud_large(19, 36) <= 0; cloud_large(19, 37) <= 0; cloud_large(19, 38) <= 0; cloud_large(19, 39) <= 0; cloud_large(19, 40) <= 0; cloud_large(19, 41) <= 0; cloud_large(19, 42) <= 0; cloud_large(19, 43) <= 0; cloud_large(19, 44) <= 0; cloud_large(19, 45) <= 0; cloud_large(19, 46) <= 0; cloud_large(19, 47) <= 0; cloud_large(19, 48) <= 1; cloud_large(19, 49) <= 1; cloud_large(19, 50) <= 1; cloud_large(19, 51) <= 1; 
cloud_large(20, 0) <= 1; cloud_large(20, 1) <= 1; cloud_large(20, 2) <= 1; cloud_large(20, 3) <= 1; cloud_large(20, 4) <= 0; cloud_large(20, 5) <= 0; cloud_large(20, 6) <= 0; cloud_large(20, 7) <= 0; cloud_large(20, 8) <= 0; cloud_large(20, 9) <= 0; cloud_large(20, 10) <= 0; cloud_large(20, 11) <= 0; cloud_large(20, 12) <= 0; cloud_large(20, 13) <= 0; cloud_large(20, 14) <= 0; cloud_large(20, 15) <= 0; cloud_large(20, 16) <= 0; cloud_large(20, 17) <= 0; cloud_large(20, 18) <= 0; cloud_large(20, 19) <= 0; cloud_large(20, 20) <= 0; cloud_large(20, 21) <= 0; cloud_large(20, 22) <= 0; cloud_large(20, 23) <= 0; cloud_large(20, 24) <= 0; cloud_large(20, 25) <= 0; cloud_large(20, 26) <= 0; cloud_large(20, 27) <= 0; cloud_large(20, 28) <= 0; cloud_large(20, 29) <= 0; cloud_large(20, 30) <= 0; cloud_large(20, 31) <= 0; cloud_large(20, 32) <= 0; cloud_large(20, 33) <= 0; cloud_large(20, 34) <= 0; cloud_large(20, 35) <= 0; cloud_large(20, 36) <= 0; cloud_large(20, 37) <= 0; cloud_large(20, 38) <= 0; cloud_large(20, 39) <= 0; cloud_large(20, 40) <= 0; cloud_large(20, 41) <= 0; cloud_large(20, 42) <= 0; cloud_large(20, 43) <= 0; cloud_large(20, 44) <= 0; cloud_large(20, 45) <= 0; cloud_large(20, 46) <= 0; cloud_large(20, 47) <= 0; cloud_large(20, 48) <= 1; cloud_large(20, 49) <= 1; cloud_large(20, 50) <= 1; cloud_large(20, 51) <= 1; 
cloud_large(21, 0) <= 1; cloud_large(21, 1) <= 1; cloud_large(21, 2) <= 1; cloud_large(21, 3) <= 1; cloud_large(21, 4) <= 0; cloud_large(21, 5) <= 0; cloud_large(21, 6) <= 0; cloud_large(21, 7) <= 0; cloud_large(21, 8) <= 0; cloud_large(21, 9) <= 0; cloud_large(21, 10) <= 0; cloud_large(21, 11) <= 0; cloud_large(21, 12) <= 0; cloud_large(21, 13) <= 0; cloud_large(21, 14) <= 0; cloud_large(21, 15) <= 0; cloud_large(21, 16) <= 0; cloud_large(21, 17) <= 0; cloud_large(21, 18) <= 0; cloud_large(21, 19) <= 0; cloud_large(21, 20) <= 0; cloud_large(21, 21) <= 0; cloud_large(21, 22) <= 0; cloud_large(21, 23) <= 0; cloud_large(21, 24) <= 0; cloud_large(21, 25) <= 0; cloud_large(21, 26) <= 0; cloud_large(21, 27) <= 0; cloud_large(21, 28) <= 0; cloud_large(21, 29) <= 0; cloud_large(21, 30) <= 0; cloud_large(21, 31) <= 0; cloud_large(21, 32) <= 0; cloud_large(21, 33) <= 0; cloud_large(21, 34) <= 0; cloud_large(21, 35) <= 0; cloud_large(21, 36) <= 0; cloud_large(21, 37) <= 0; cloud_large(21, 38) <= 0; cloud_large(21, 39) <= 0; cloud_large(21, 40) <= 0; cloud_large(21, 41) <= 0; cloud_large(21, 42) <= 0; cloud_large(21, 43) <= 0; cloud_large(21, 44) <= 0; cloud_large(21, 45) <= 0; cloud_large(21, 46) <= 0; cloud_large(21, 47) <= 0; cloud_large(21, 48) <= 1; cloud_large(21, 49) <= 1; cloud_large(21, 50) <= 1; cloud_large(21, 51) <= 1; 
cloud_large(22, 0) <= 1; cloud_large(22, 1) <= 1; cloud_large(22, 2) <= 1; cloud_large(22, 3) <= 1; cloud_large(22, 4) <= 0; cloud_large(22, 5) <= 0; cloud_large(22, 6) <= 0; cloud_large(22, 7) <= 0; cloud_large(22, 8) <= 0; cloud_large(22, 9) <= 0; cloud_large(22, 10) <= 0; cloud_large(22, 11) <= 0; cloud_large(22, 12) <= 0; cloud_large(22, 13) <= 0; cloud_large(22, 14) <= 0; cloud_large(22, 15) <= 0; cloud_large(22, 16) <= 0; cloud_large(22, 17) <= 0; cloud_large(22, 18) <= 0; cloud_large(22, 19) <= 0; cloud_large(22, 20) <= 0; cloud_large(22, 21) <= 0; cloud_large(22, 22) <= 0; cloud_large(22, 23) <= 0; cloud_large(22, 24) <= 0; cloud_large(22, 25) <= 0; cloud_large(22, 26) <= 0; cloud_large(22, 27) <= 0; cloud_large(22, 28) <= 0; cloud_large(22, 29) <= 0; cloud_large(22, 30) <= 0; cloud_large(22, 31) <= 0; cloud_large(22, 32) <= 0; cloud_large(22, 33) <= 0; cloud_large(22, 34) <= 0; cloud_large(22, 35) <= 0; cloud_large(22, 36) <= 0; cloud_large(22, 37) <= 0; cloud_large(22, 38) <= 0; cloud_large(22, 39) <= 0; cloud_large(22, 40) <= 0; cloud_large(22, 41) <= 0; cloud_large(22, 42) <= 0; cloud_large(22, 43) <= 0; cloud_large(22, 44) <= 0; cloud_large(22, 45) <= 0; cloud_large(22, 46) <= 0; cloud_large(22, 47) <= 0; cloud_large(22, 48) <= 1; cloud_large(22, 49) <= 1; cloud_large(22, 50) <= 1; cloud_large(22, 51) <= 1; 
cloud_large(23, 0) <= 1; cloud_large(23, 1) <= 1; cloud_large(23, 2) <= 1; cloud_large(23, 3) <= 1; cloud_large(23, 4) <= 0; cloud_large(23, 5) <= 0; cloud_large(23, 6) <= 0; cloud_large(23, 7) <= 0; cloud_large(23, 8) <= 0; cloud_large(23, 9) <= 0; cloud_large(23, 10) <= 0; cloud_large(23, 11) <= 0; cloud_large(23, 12) <= 0; cloud_large(23, 13) <= 0; cloud_large(23, 14) <= 0; cloud_large(23, 15) <= 0; cloud_large(23, 16) <= 0; cloud_large(23, 17) <= 0; cloud_large(23, 18) <= 0; cloud_large(23, 19) <= 0; cloud_large(23, 20) <= 0; cloud_large(23, 21) <= 0; cloud_large(23, 22) <= 0; cloud_large(23, 23) <= 0; cloud_large(23, 24) <= 0; cloud_large(23, 25) <= 0; cloud_large(23, 26) <= 0; cloud_large(23, 27) <= 0; cloud_large(23, 28) <= 0; cloud_large(23, 29) <= 0; cloud_large(23, 30) <= 0; cloud_large(23, 31) <= 0; cloud_large(23, 32) <= 0; cloud_large(23, 33) <= 0; cloud_large(23, 34) <= 0; cloud_large(23, 35) <= 0; cloud_large(23, 36) <= 0; cloud_large(23, 37) <= 0; cloud_large(23, 38) <= 0; cloud_large(23, 39) <= 0; cloud_large(23, 40) <= 0; cloud_large(23, 41) <= 0; cloud_large(23, 42) <= 0; cloud_large(23, 43) <= 0; cloud_large(23, 44) <= 0; cloud_large(23, 45) <= 0; cloud_large(23, 46) <= 0; cloud_large(23, 47) <= 0; cloud_large(23, 48) <= 1; cloud_large(23, 49) <= 1; cloud_large(23, 50) <= 1; cloud_large(23, 51) <= 1; 
cloud_large(24, 0) <= 1; cloud_large(24, 1) <= 1; cloud_large(24, 2) <= 1; cloud_large(24, 3) <= 1; cloud_large(24, 4) <= 0; cloud_large(24, 5) <= 0; cloud_large(24, 6) <= 0; cloud_large(24, 7) <= 0; cloud_large(24, 8) <= 0; cloud_large(24, 9) <= 0; cloud_large(24, 10) <= 0; cloud_large(24, 11) <= 0; cloud_large(24, 12) <= 0; cloud_large(24, 13) <= 0; cloud_large(24, 14) <= 0; cloud_large(24, 15) <= 0; cloud_large(24, 16) <= 0; cloud_large(24, 17) <= 0; cloud_large(24, 18) <= 0; cloud_large(24, 19) <= 0; cloud_large(24, 20) <= 0; cloud_large(24, 21) <= 0; cloud_large(24, 22) <= 0; cloud_large(24, 23) <= 0; cloud_large(24, 24) <= 0; cloud_large(24, 25) <= 0; cloud_large(24, 26) <= 0; cloud_large(24, 27) <= 0; cloud_large(24, 28) <= 0; cloud_large(24, 29) <= 0; cloud_large(24, 30) <= 0; cloud_large(24, 31) <= 0; cloud_large(24, 32) <= 0; cloud_large(24, 33) <= 0; cloud_large(24, 34) <= 0; cloud_large(24, 35) <= 0; cloud_large(24, 36) <= 0; cloud_large(24, 37) <= 0; cloud_large(24, 38) <= 0; cloud_large(24, 39) <= 0; cloud_large(24, 40) <= 0; cloud_large(24, 41) <= 0; cloud_large(24, 42) <= 0; cloud_large(24, 43) <= 0; cloud_large(24, 44) <= 0; cloud_large(24, 45) <= 0; cloud_large(24, 46) <= 0; cloud_large(24, 47) <= 0; cloud_large(24, 48) <= 1; cloud_large(24, 49) <= 1; cloud_large(24, 50) <= 1; cloud_large(24, 51) <= 1; 
cloud_large(25, 0) <= 1; cloud_large(25, 1) <= 1; cloud_large(25, 2) <= 1; cloud_large(25, 3) <= 1; cloud_large(25, 4) <= 0; cloud_large(25, 5) <= 0; cloud_large(25, 6) <= 0; cloud_large(25, 7) <= 0; cloud_large(25, 8) <= 0; cloud_large(25, 9) <= 0; cloud_large(25, 10) <= 0; cloud_large(25, 11) <= 0; cloud_large(25, 12) <= 0; cloud_large(25, 13) <= 0; cloud_large(25, 14) <= 0; cloud_large(25, 15) <= 0; cloud_large(25, 16) <= 0; cloud_large(25, 17) <= 0; cloud_large(25, 18) <= 0; cloud_large(25, 19) <= 0; cloud_large(25, 20) <= 0; cloud_large(25, 21) <= 0; cloud_large(25, 22) <= 0; cloud_large(25, 23) <= 0; cloud_large(25, 24) <= 0; cloud_large(25, 25) <= 0; cloud_large(25, 26) <= 0; cloud_large(25, 27) <= 0; cloud_large(25, 28) <= 0; cloud_large(25, 29) <= 0; cloud_large(25, 30) <= 0; cloud_large(25, 31) <= 0; cloud_large(25, 32) <= 0; cloud_large(25, 33) <= 0; cloud_large(25, 34) <= 0; cloud_large(25, 35) <= 0; cloud_large(25, 36) <= 0; cloud_large(25, 37) <= 0; cloud_large(25, 38) <= 0; cloud_large(25, 39) <= 0; cloud_large(25, 40) <= 0; cloud_large(25, 41) <= 0; cloud_large(25, 42) <= 0; cloud_large(25, 43) <= 0; cloud_large(25, 44) <= 0; cloud_large(25, 45) <= 0; cloud_large(25, 46) <= 0; cloud_large(25, 47) <= 0; cloud_large(25, 48) <= 1; cloud_large(25, 49) <= 1; cloud_large(25, 50) <= 1; cloud_large(25, 51) <= 1; 
cloud_large(26, 0) <= 1; cloud_large(26, 1) <= 1; cloud_large(26, 2) <= 1; cloud_large(26, 3) <= 1; cloud_large(26, 4) <= 0; cloud_large(26, 5) <= 0; cloud_large(26, 6) <= 0; cloud_large(26, 7) <= 0; cloud_large(26, 8) <= 0; cloud_large(26, 9) <= 0; cloud_large(26, 10) <= 0; cloud_large(26, 11) <= 0; cloud_large(26, 12) <= 0; cloud_large(26, 13) <= 0; cloud_large(26, 14) <= 0; cloud_large(26, 15) <= 0; cloud_large(26, 16) <= 0; cloud_large(26, 17) <= 0; cloud_large(26, 18) <= 0; cloud_large(26, 19) <= 0; cloud_large(26, 20) <= 0; cloud_large(26, 21) <= 0; cloud_large(26, 22) <= 0; cloud_large(26, 23) <= 0; cloud_large(26, 24) <= 0; cloud_large(26, 25) <= 0; cloud_large(26, 26) <= 0; cloud_large(26, 27) <= 0; cloud_large(26, 28) <= 0; cloud_large(26, 29) <= 0; cloud_large(26, 30) <= 0; cloud_large(26, 31) <= 0; cloud_large(26, 32) <= 0; cloud_large(26, 33) <= 0; cloud_large(26, 34) <= 0; cloud_large(26, 35) <= 0; cloud_large(26, 36) <= 0; cloud_large(26, 37) <= 0; cloud_large(26, 38) <= 0; cloud_large(26, 39) <= 0; cloud_large(26, 40) <= 0; cloud_large(26, 41) <= 0; cloud_large(26, 42) <= 0; cloud_large(26, 43) <= 0; cloud_large(26, 44) <= 0; cloud_large(26, 45) <= 0; cloud_large(26, 46) <= 0; cloud_large(26, 47) <= 0; cloud_large(26, 48) <= 1; cloud_large(26, 49) <= 1; cloud_large(26, 50) <= 1; cloud_large(26, 51) <= 1; 
cloud_large(27, 0) <= 1; cloud_large(27, 1) <= 1; cloud_large(27, 2) <= 1; cloud_large(27, 3) <= 1; cloud_large(27, 4) <= 0; cloud_large(27, 5) <= 0; cloud_large(27, 6) <= 0; cloud_large(27, 7) <= 0; cloud_large(27, 8) <= 0; cloud_large(27, 9) <= 0; cloud_large(27, 10) <= 0; cloud_large(27, 11) <= 0; cloud_large(27, 12) <= 0; cloud_large(27, 13) <= 0; cloud_large(27, 14) <= 0; cloud_large(27, 15) <= 0; cloud_large(27, 16) <= 0; cloud_large(27, 17) <= 0; cloud_large(27, 18) <= 0; cloud_large(27, 19) <= 0; cloud_large(27, 20) <= 0; cloud_large(27, 21) <= 0; cloud_large(27, 22) <= 0; cloud_large(27, 23) <= 0; cloud_large(27, 24) <= 0; cloud_large(27, 25) <= 0; cloud_large(27, 26) <= 0; cloud_large(27, 27) <= 0; cloud_large(27, 28) <= 0; cloud_large(27, 29) <= 0; cloud_large(27, 30) <= 0; cloud_large(27, 31) <= 0; cloud_large(27, 32) <= 0; cloud_large(27, 33) <= 0; cloud_large(27, 34) <= 0; cloud_large(27, 35) <= 0; cloud_large(27, 36) <= 0; cloud_large(27, 37) <= 0; cloud_large(27, 38) <= 0; cloud_large(27, 39) <= 0; cloud_large(27, 40) <= 0; cloud_large(27, 41) <= 0; cloud_large(27, 42) <= 0; cloud_large(27, 43) <= 0; cloud_large(27, 44) <= 0; cloud_large(27, 45) <= 0; cloud_large(27, 46) <= 0; cloud_large(27, 47) <= 0; cloud_large(27, 48) <= 1; cloud_large(27, 49) <= 1; cloud_large(27, 50) <= 1; cloud_large(27, 51) <= 1; 
cloud_large(28, 0) <= 2; cloud_large(28, 1) <= 2; cloud_large(28, 2) <= 2; cloud_large(28, 3) <= 2; cloud_large(28, 4) <= 1; cloud_large(28, 5) <= 1; cloud_large(28, 6) <= 1; cloud_large(28, 7) <= 1; cloud_large(28, 8) <= 0; cloud_large(28, 9) <= 0; cloud_large(28, 10) <= 0; cloud_large(28, 11) <= 0; cloud_large(28, 12) <= 0; cloud_large(28, 13) <= 0; cloud_large(28, 14) <= 0; cloud_large(28, 15) <= 0; cloud_large(28, 16) <= 0; cloud_large(28, 17) <= 0; cloud_large(28, 18) <= 0; cloud_large(28, 19) <= 0; cloud_large(28, 20) <= 0; cloud_large(28, 21) <= 0; cloud_large(28, 22) <= 0; cloud_large(28, 23) <= 0; cloud_large(28, 24) <= 0; cloud_large(28, 25) <= 0; cloud_large(28, 26) <= 0; cloud_large(28, 27) <= 0; cloud_large(28, 28) <= 0; cloud_large(28, 29) <= 0; cloud_large(28, 30) <= 0; cloud_large(28, 31) <= 0; cloud_large(28, 32) <= 0; cloud_large(28, 33) <= 0; cloud_large(28, 34) <= 0; cloud_large(28, 35) <= 0; cloud_large(28, 36) <= 0; cloud_large(28, 37) <= 0; cloud_large(28, 38) <= 0; cloud_large(28, 39) <= 0; cloud_large(28, 40) <= 0; cloud_large(28, 41) <= 0; cloud_large(28, 42) <= 0; cloud_large(28, 43) <= 0; cloud_large(28, 44) <= 1; cloud_large(28, 45) <= 1; cloud_large(28, 46) <= 1; cloud_large(28, 47) <= 1; cloud_large(28, 48) <= 2; cloud_large(28, 49) <= 2; cloud_large(28, 50) <= 2; cloud_large(28, 51) <= 2; 
cloud_large(29, 0) <= 2; cloud_large(29, 1) <= 2; cloud_large(29, 2) <= 2; cloud_large(29, 3) <= 2; cloud_large(29, 4) <= 1; cloud_large(29, 5) <= 1; cloud_large(29, 6) <= 1; cloud_large(29, 7) <= 1; cloud_large(29, 8) <= 0; cloud_large(29, 9) <= 0; cloud_large(29, 10) <= 0; cloud_large(29, 11) <= 0; cloud_large(29, 12) <= 0; cloud_large(29, 13) <= 0; cloud_large(29, 14) <= 0; cloud_large(29, 15) <= 0; cloud_large(29, 16) <= 0; cloud_large(29, 17) <= 0; cloud_large(29, 18) <= 0; cloud_large(29, 19) <= 0; cloud_large(29, 20) <= 0; cloud_large(29, 21) <= 0; cloud_large(29, 22) <= 0; cloud_large(29, 23) <= 0; cloud_large(29, 24) <= 0; cloud_large(29, 25) <= 0; cloud_large(29, 26) <= 0; cloud_large(29, 27) <= 0; cloud_large(29, 28) <= 0; cloud_large(29, 29) <= 0; cloud_large(29, 30) <= 0; cloud_large(29, 31) <= 0; cloud_large(29, 32) <= 0; cloud_large(29, 33) <= 0; cloud_large(29, 34) <= 0; cloud_large(29, 35) <= 0; cloud_large(29, 36) <= 0; cloud_large(29, 37) <= 0; cloud_large(29, 38) <= 0; cloud_large(29, 39) <= 0; cloud_large(29, 40) <= 0; cloud_large(29, 41) <= 0; cloud_large(29, 42) <= 0; cloud_large(29, 43) <= 0; cloud_large(29, 44) <= 1; cloud_large(29, 45) <= 1; cloud_large(29, 46) <= 1; cloud_large(29, 47) <= 1; cloud_large(29, 48) <= 2; cloud_large(29, 49) <= 2; cloud_large(29, 50) <= 2; cloud_large(29, 51) <= 2; 
cloud_large(30, 0) <= 2; cloud_large(30, 1) <= 2; cloud_large(30, 2) <= 2; cloud_large(30, 3) <= 2; cloud_large(30, 4) <= 1; cloud_large(30, 5) <= 1; cloud_large(30, 6) <= 1; cloud_large(30, 7) <= 1; cloud_large(30, 8) <= 0; cloud_large(30, 9) <= 0; cloud_large(30, 10) <= 0; cloud_large(30, 11) <= 0; cloud_large(30, 12) <= 0; cloud_large(30, 13) <= 0; cloud_large(30, 14) <= 0; cloud_large(30, 15) <= 0; cloud_large(30, 16) <= 0; cloud_large(30, 17) <= 0; cloud_large(30, 18) <= 0; cloud_large(30, 19) <= 0; cloud_large(30, 20) <= 0; cloud_large(30, 21) <= 0; cloud_large(30, 22) <= 0; cloud_large(30, 23) <= 0; cloud_large(30, 24) <= 0; cloud_large(30, 25) <= 0; cloud_large(30, 26) <= 0; cloud_large(30, 27) <= 0; cloud_large(30, 28) <= 0; cloud_large(30, 29) <= 0; cloud_large(30, 30) <= 0; cloud_large(30, 31) <= 0; cloud_large(30, 32) <= 0; cloud_large(30, 33) <= 0; cloud_large(30, 34) <= 0; cloud_large(30, 35) <= 0; cloud_large(30, 36) <= 0; cloud_large(30, 37) <= 0; cloud_large(30, 38) <= 0; cloud_large(30, 39) <= 0; cloud_large(30, 40) <= 0; cloud_large(30, 41) <= 0; cloud_large(30, 42) <= 0; cloud_large(30, 43) <= 0; cloud_large(30, 44) <= 1; cloud_large(30, 45) <= 1; cloud_large(30, 46) <= 1; cloud_large(30, 47) <= 1; cloud_large(30, 48) <= 2; cloud_large(30, 49) <= 2; cloud_large(30, 50) <= 2; cloud_large(30, 51) <= 2; 
cloud_large(31, 0) <= 2; cloud_large(31, 1) <= 2; cloud_large(31, 2) <= 2; cloud_large(31, 3) <= 2; cloud_large(31, 4) <= 1; cloud_large(31, 5) <= 1; cloud_large(31, 6) <= 1; cloud_large(31, 7) <= 1; cloud_large(31, 8) <= 0; cloud_large(31, 9) <= 0; cloud_large(31, 10) <= 0; cloud_large(31, 11) <= 0; cloud_large(31, 12) <= 0; cloud_large(31, 13) <= 0; cloud_large(31, 14) <= 0; cloud_large(31, 15) <= 0; cloud_large(31, 16) <= 0; cloud_large(31, 17) <= 0; cloud_large(31, 18) <= 0; cloud_large(31, 19) <= 0; cloud_large(31, 20) <= 0; cloud_large(31, 21) <= 0; cloud_large(31, 22) <= 0; cloud_large(31, 23) <= 0; cloud_large(31, 24) <= 0; cloud_large(31, 25) <= 0; cloud_large(31, 26) <= 0; cloud_large(31, 27) <= 0; cloud_large(31, 28) <= 0; cloud_large(31, 29) <= 0; cloud_large(31, 30) <= 0; cloud_large(31, 31) <= 0; cloud_large(31, 32) <= 0; cloud_large(31, 33) <= 0; cloud_large(31, 34) <= 0; cloud_large(31, 35) <= 0; cloud_large(31, 36) <= 0; cloud_large(31, 37) <= 0; cloud_large(31, 38) <= 0; cloud_large(31, 39) <= 0; cloud_large(31, 40) <= 0; cloud_large(31, 41) <= 0; cloud_large(31, 42) <= 0; cloud_large(31, 43) <= 0; cloud_large(31, 44) <= 1; cloud_large(31, 45) <= 1; cloud_large(31, 46) <= 1; cloud_large(31, 47) <= 1; cloud_large(31, 48) <= 2; cloud_large(31, 49) <= 2; cloud_large(31, 50) <= 2; cloud_large(31, 51) <= 2; 
cloud_large(32, 0) <= 2; cloud_large(32, 1) <= 2; cloud_large(32, 2) <= 2; cloud_large(32, 3) <= 2; cloud_large(32, 4) <= 2; cloud_large(32, 5) <= 2; cloud_large(32, 6) <= 2; cloud_large(32, 7) <= 2; cloud_large(32, 8) <= 1; cloud_large(32, 9) <= 1; cloud_large(32, 10) <= 1; cloud_large(32, 11) <= 1; cloud_large(32, 12) <= 1; cloud_large(32, 13) <= 1; cloud_large(32, 14) <= 1; cloud_large(32, 15) <= 1; cloud_large(32, 16) <= 1; cloud_large(32, 17) <= 1; cloud_large(32, 18) <= 1; cloud_large(32, 19) <= 1; cloud_large(32, 20) <= 1; cloud_large(32, 21) <= 1; cloud_large(32, 22) <= 1; cloud_large(32, 23) <= 1; cloud_large(32, 24) <= 1; cloud_large(32, 25) <= 1; cloud_large(32, 26) <= 1; cloud_large(32, 27) <= 1; cloud_large(32, 28) <= 1; cloud_large(32, 29) <= 1; cloud_large(32, 30) <= 1; cloud_large(32, 31) <= 1; cloud_large(32, 32) <= 1; cloud_large(32, 33) <= 1; cloud_large(32, 34) <= 1; cloud_large(32, 35) <= 1; cloud_large(32, 36) <= 1; cloud_large(32, 37) <= 1; cloud_large(32, 38) <= 1; cloud_large(32, 39) <= 1; cloud_large(32, 40) <= 1; cloud_large(32, 41) <= 1; cloud_large(32, 42) <= 1; cloud_large(32, 43) <= 1; cloud_large(32, 44) <= 2; cloud_large(32, 45) <= 2; cloud_large(32, 46) <= 2; cloud_large(32, 47) <= 2; cloud_large(32, 48) <= 2; cloud_large(32, 49) <= 2; cloud_large(32, 50) <= 2; cloud_large(32, 51) <= 2; 
cloud_large(33, 0) <= 2; cloud_large(33, 1) <= 2; cloud_large(33, 2) <= 2; cloud_large(33, 3) <= 2; cloud_large(33, 4) <= 2; cloud_large(33, 5) <= 2; cloud_large(33, 6) <= 2; cloud_large(33, 7) <= 2; cloud_large(33, 8) <= 1; cloud_large(33, 9) <= 1; cloud_large(33, 10) <= 1; cloud_large(33, 11) <= 1; cloud_large(33, 12) <= 1; cloud_large(33, 13) <= 1; cloud_large(33, 14) <= 1; cloud_large(33, 15) <= 1; cloud_large(33, 16) <= 1; cloud_large(33, 17) <= 1; cloud_large(33, 18) <= 1; cloud_large(33, 19) <= 1; cloud_large(33, 20) <= 1; cloud_large(33, 21) <= 1; cloud_large(33, 22) <= 1; cloud_large(33, 23) <= 1; cloud_large(33, 24) <= 1; cloud_large(33, 25) <= 1; cloud_large(33, 26) <= 1; cloud_large(33, 27) <= 1; cloud_large(33, 28) <= 1; cloud_large(33, 29) <= 1; cloud_large(33, 30) <= 1; cloud_large(33, 31) <= 1; cloud_large(33, 32) <= 1; cloud_large(33, 33) <= 1; cloud_large(33, 34) <= 1; cloud_large(33, 35) <= 1; cloud_large(33, 36) <= 1; cloud_large(33, 37) <= 1; cloud_large(33, 38) <= 1; cloud_large(33, 39) <= 1; cloud_large(33, 40) <= 1; cloud_large(33, 41) <= 1; cloud_large(33, 42) <= 1; cloud_large(33, 43) <= 1; cloud_large(33, 44) <= 2; cloud_large(33, 45) <= 2; cloud_large(33, 46) <= 2; cloud_large(33, 47) <= 2; cloud_large(33, 48) <= 2; cloud_large(33, 49) <= 2; cloud_large(33, 50) <= 2; cloud_large(33, 51) <= 2; 
cloud_large(34, 0) <= 2; cloud_large(34, 1) <= 2; cloud_large(34, 2) <= 2; cloud_large(34, 3) <= 2; cloud_large(34, 4) <= 2; cloud_large(34, 5) <= 2; cloud_large(34, 6) <= 2; cloud_large(34, 7) <= 2; cloud_large(34, 8) <= 1; cloud_large(34, 9) <= 1; cloud_large(34, 10) <= 1; cloud_large(34, 11) <= 1; cloud_large(34, 12) <= 1; cloud_large(34, 13) <= 1; cloud_large(34, 14) <= 1; cloud_large(34, 15) <= 1; cloud_large(34, 16) <= 1; cloud_large(34, 17) <= 1; cloud_large(34, 18) <= 1; cloud_large(34, 19) <= 1; cloud_large(34, 20) <= 1; cloud_large(34, 21) <= 1; cloud_large(34, 22) <= 1; cloud_large(34, 23) <= 1; cloud_large(34, 24) <= 1; cloud_large(34, 25) <= 1; cloud_large(34, 26) <= 1; cloud_large(34, 27) <= 1; cloud_large(34, 28) <= 1; cloud_large(34, 29) <= 1; cloud_large(34, 30) <= 1; cloud_large(34, 31) <= 1; cloud_large(34, 32) <= 1; cloud_large(34, 33) <= 1; cloud_large(34, 34) <= 1; cloud_large(34, 35) <= 1; cloud_large(34, 36) <= 1; cloud_large(34, 37) <= 1; cloud_large(34, 38) <= 1; cloud_large(34, 39) <= 1; cloud_large(34, 40) <= 1; cloud_large(34, 41) <= 1; cloud_large(34, 42) <= 1; cloud_large(34, 43) <= 1; cloud_large(34, 44) <= 2; cloud_large(34, 45) <= 2; cloud_large(34, 46) <= 2; cloud_large(34, 47) <= 2; cloud_large(34, 48) <= 2; cloud_large(34, 49) <= 2; cloud_large(34, 50) <= 2; cloud_large(34, 51) <= 2; 
cloud_large(35, 0) <= 2; cloud_large(35, 1) <= 2; cloud_large(35, 2) <= 2; cloud_large(35, 3) <= 2; cloud_large(35, 4) <= 2; cloud_large(35, 5) <= 2; cloud_large(35, 6) <= 2; cloud_large(35, 7) <= 2; cloud_large(35, 8) <= 1; cloud_large(35, 9) <= 1; cloud_large(35, 10) <= 1; cloud_large(35, 11) <= 1; cloud_large(35, 12) <= 1; cloud_large(35, 13) <= 1; cloud_large(35, 14) <= 1; cloud_large(35, 15) <= 1; cloud_large(35, 16) <= 1; cloud_large(35, 17) <= 1; cloud_large(35, 18) <= 1; cloud_large(35, 19) <= 1; cloud_large(35, 20) <= 1; cloud_large(35, 21) <= 1; cloud_large(35, 22) <= 1; cloud_large(35, 23) <= 1; cloud_large(35, 24) <= 1; cloud_large(35, 25) <= 1; cloud_large(35, 26) <= 1; cloud_large(35, 27) <= 1; cloud_large(35, 28) <= 1; cloud_large(35, 29) <= 1; cloud_large(35, 30) <= 1; cloud_large(35, 31) <= 1; cloud_large(35, 32) <= 1; cloud_large(35, 33) <= 1; cloud_large(35, 34) <= 1; cloud_large(35, 35) <= 1; cloud_large(35, 36) <= 1; cloud_large(35, 37) <= 1; cloud_large(35, 38) <= 1; cloud_large(35, 39) <= 1; cloud_large(35, 40) <= 1; cloud_large(35, 41) <= 1; cloud_large(35, 42) <= 1; cloud_large(35, 43) <= 1; cloud_large(35, 44) <= 2; cloud_large(35, 45) <= 2; cloud_large(35, 46) <= 2; cloud_large(35, 47) <= 2; cloud_large(35, 48) <= 2; cloud_large(35, 49) <= 2; cloud_large(35, 50) <= 2; cloud_large(35, 51) <= 2; 

cloud_small(0, 0) <= 2; cloud_small(0, 1) <= 2; cloud_small(0, 2) <= 2; cloud_small(0, 3) <= 2; cloud_small(0, 4) <= 2; cloud_small(0, 5) <= 2; cloud_small(0, 6) <= 2; cloud_small(0, 7) <= 2; cloud_small(0, 8) <= 2; cloud_small(0, 9) <= 2; cloud_small(0, 10) <= 2; cloud_small(0, 11) <= 2; cloud_small(0, 12) <= 2; cloud_small(0, 13) <= 2; cloud_small(0, 14) <= 2; cloud_small(0, 15) <= 1; cloud_small(0, 16) <= 1; cloud_small(0, 17) <= 1; cloud_small(0, 18) <= 1; cloud_small(0, 19) <= 1; cloud_small(0, 20) <= 1; cloud_small(0, 21) <= 1; cloud_small(0, 22) <= 1; cloud_small(0, 23) <= 1; cloud_small(0, 24) <= 2; cloud_small(0, 25) <= 2; cloud_small(0, 26) <= 2; cloud_small(0, 27) <= 2; cloud_small(0, 28) <= 2; cloud_small(0, 29) <= 2; cloud_small(0, 30) <= 2; cloud_small(0, 31) <= 2; cloud_small(0, 32) <= 2; cloud_small(0, 33) <= 2; cloud_small(0, 34) <= 2; cloud_small(0, 35) <= 2; cloud_small(0, 36) <= 2; cloud_small(0, 37) <= 2; cloud_small(0, 38) <= 2; 
cloud_small(1, 0) <= 2; cloud_small(1, 1) <= 2; cloud_small(1, 2) <= 2; cloud_small(1, 3) <= 2; cloud_small(1, 4) <= 2; cloud_small(1, 5) <= 2; cloud_small(1, 6) <= 2; cloud_small(1, 7) <= 2; cloud_small(1, 8) <= 2; cloud_small(1, 9) <= 2; cloud_small(1, 10) <= 2; cloud_small(1, 11) <= 2; cloud_small(1, 12) <= 2; cloud_small(1, 13) <= 2; cloud_small(1, 14) <= 2; cloud_small(1, 15) <= 1; cloud_small(1, 16) <= 1; cloud_small(1, 17) <= 1; cloud_small(1, 18) <= 1; cloud_small(1, 19) <= 1; cloud_small(1, 20) <= 1; cloud_small(1, 21) <= 1; cloud_small(1, 22) <= 1; cloud_small(1, 23) <= 1; cloud_small(1, 24) <= 2; cloud_small(1, 25) <= 2; cloud_small(1, 26) <= 2; cloud_small(1, 27) <= 2; cloud_small(1, 28) <= 2; cloud_small(1, 29) <= 2; cloud_small(1, 30) <= 2; cloud_small(1, 31) <= 2; cloud_small(1, 32) <= 2; cloud_small(1, 33) <= 2; cloud_small(1, 34) <= 2; cloud_small(1, 35) <= 2; cloud_small(1, 36) <= 2; cloud_small(1, 37) <= 2; cloud_small(1, 38) <= 2; 
cloud_small(2, 0) <= 2; cloud_small(2, 1) <= 2; cloud_small(2, 2) <= 2; cloud_small(2, 3) <= 2; cloud_small(2, 4) <= 2; cloud_small(2, 5) <= 2; cloud_small(2, 6) <= 2; cloud_small(2, 7) <= 2; cloud_small(2, 8) <= 2; cloud_small(2, 9) <= 2; cloud_small(2, 10) <= 2; cloud_small(2, 11) <= 2; cloud_small(2, 12) <= 2; cloud_small(2, 13) <= 2; cloud_small(2, 14) <= 2; cloud_small(2, 15) <= 1; cloud_small(2, 16) <= 1; cloud_small(2, 17) <= 1; cloud_small(2, 18) <= 1; cloud_small(2, 19) <= 1; cloud_small(2, 20) <= 1; cloud_small(2, 21) <= 1; cloud_small(2, 22) <= 1; cloud_small(2, 23) <= 1; cloud_small(2, 24) <= 2; cloud_small(2, 25) <= 2; cloud_small(2, 26) <= 2; cloud_small(2, 27) <= 2; cloud_small(2, 28) <= 2; cloud_small(2, 29) <= 2; cloud_small(2, 30) <= 2; cloud_small(2, 31) <= 2; cloud_small(2, 32) <= 2; cloud_small(2, 33) <= 2; cloud_small(2, 34) <= 2; cloud_small(2, 35) <= 2; cloud_small(2, 36) <= 2; cloud_small(2, 37) <= 2; cloud_small(2, 38) <= 2; 
cloud_small(3, 0) <= 2; cloud_small(3, 1) <= 2; cloud_small(3, 2) <= 2; cloud_small(3, 3) <= 2; cloud_small(3, 4) <= 2; cloud_small(3, 5) <= 2; cloud_small(3, 6) <= 2; cloud_small(3, 7) <= 2; cloud_small(3, 8) <= 2; cloud_small(3, 9) <= 2; cloud_small(3, 10) <= 2; cloud_small(3, 11) <= 2; cloud_small(3, 12) <= 1; cloud_small(3, 13) <= 1; cloud_small(3, 14) <= 1; cloud_small(3, 15) <= 0; cloud_small(3, 16) <= 0; cloud_small(3, 17) <= 0; cloud_small(3, 18) <= 0; cloud_small(3, 19) <= 0; cloud_small(3, 20) <= 0; cloud_small(3, 21) <= 0; cloud_small(3, 22) <= 0; cloud_small(3, 23) <= 0; cloud_small(3, 24) <= 1; cloud_small(3, 25) <= 1; cloud_small(3, 26) <= 1; cloud_small(3, 27) <= 2; cloud_small(3, 28) <= 2; cloud_small(3, 29) <= 2; cloud_small(3, 30) <= 2; cloud_small(3, 31) <= 2; cloud_small(3, 32) <= 2; cloud_small(3, 33) <= 2; cloud_small(3, 34) <= 2; cloud_small(3, 35) <= 2; cloud_small(3, 36) <= 2; cloud_small(3, 37) <= 2; cloud_small(3, 38) <= 2; 
cloud_small(4, 0) <= 2; cloud_small(4, 1) <= 2; cloud_small(4, 2) <= 2; cloud_small(4, 3) <= 2; cloud_small(4, 4) <= 2; cloud_small(4, 5) <= 2; cloud_small(4, 6) <= 2; cloud_small(4, 7) <= 2; cloud_small(4, 8) <= 2; cloud_small(4, 9) <= 2; cloud_small(4, 10) <= 2; cloud_small(4, 11) <= 2; cloud_small(4, 12) <= 1; cloud_small(4, 13) <= 1; cloud_small(4, 14) <= 1; cloud_small(4, 15) <= 0; cloud_small(4, 16) <= 0; cloud_small(4, 17) <= 0; cloud_small(4, 18) <= 0; cloud_small(4, 19) <= 0; cloud_small(4, 20) <= 0; cloud_small(4, 21) <= 0; cloud_small(4, 22) <= 0; cloud_small(4, 23) <= 0; cloud_small(4, 24) <= 1; cloud_small(4, 25) <= 1; cloud_small(4, 26) <= 1; cloud_small(4, 27) <= 2; cloud_small(4, 28) <= 2; cloud_small(4, 29) <= 2; cloud_small(4, 30) <= 2; cloud_small(4, 31) <= 2; cloud_small(4, 32) <= 2; cloud_small(4, 33) <= 2; cloud_small(4, 34) <= 2; cloud_small(4, 35) <= 2; cloud_small(4, 36) <= 2; cloud_small(4, 37) <= 2; cloud_small(4, 38) <= 2; 
cloud_small(5, 0) <= 2; cloud_small(5, 1) <= 2; cloud_small(5, 2) <= 2; cloud_small(5, 3) <= 2; cloud_small(5, 4) <= 2; cloud_small(5, 5) <= 2; cloud_small(5, 6) <= 2; cloud_small(5, 7) <= 2; cloud_small(5, 8) <= 2; cloud_small(5, 9) <= 2; cloud_small(5, 10) <= 2; cloud_small(5, 11) <= 2; cloud_small(5, 12) <= 1; cloud_small(5, 13) <= 1; cloud_small(5, 14) <= 1; cloud_small(5, 15) <= 0; cloud_small(5, 16) <= 0; cloud_small(5, 17) <= 0; cloud_small(5, 18) <= 0; cloud_small(5, 19) <= 0; cloud_small(5, 20) <= 0; cloud_small(5, 21) <= 0; cloud_small(5, 22) <= 0; cloud_small(5, 23) <= 0; cloud_small(5, 24) <= 1; cloud_small(5, 25) <= 1; cloud_small(5, 26) <= 1; cloud_small(5, 27) <= 2; cloud_small(5, 28) <= 2; cloud_small(5, 29) <= 2; cloud_small(5, 30) <= 2; cloud_small(5, 31) <= 2; cloud_small(5, 32) <= 2; cloud_small(5, 33) <= 2; cloud_small(5, 34) <= 2; cloud_small(5, 35) <= 2; cloud_small(5, 36) <= 2; cloud_small(5, 37) <= 2; cloud_small(5, 38) <= 2; 
cloud_small(6, 0) <= 2; cloud_small(6, 1) <= 2; cloud_small(6, 2) <= 2; cloud_small(6, 3) <= 2; cloud_small(6, 4) <= 2; cloud_small(6, 5) <= 2; cloud_small(6, 6) <= 1; cloud_small(6, 7) <= 1; cloud_small(6, 8) <= 1; cloud_small(6, 9) <= 1; cloud_small(6, 10) <= 1; cloud_small(6, 11) <= 1; cloud_small(6, 12) <= 0; cloud_small(6, 13) <= 0; cloud_small(6, 14) <= 0; cloud_small(6, 15) <= 0; cloud_small(6, 16) <= 0; cloud_small(6, 17) <= 0; cloud_small(6, 18) <= 0; cloud_small(6, 19) <= 0; cloud_small(6, 20) <= 0; cloud_small(6, 21) <= 0; cloud_small(6, 22) <= 0; cloud_small(6, 23) <= 0; cloud_small(6, 24) <= 0; cloud_small(6, 25) <= 0; cloud_small(6, 26) <= 0; cloud_small(6, 27) <= 1; cloud_small(6, 28) <= 1; cloud_small(6, 29) <= 1; cloud_small(6, 30) <= 2; cloud_small(6, 31) <= 2; cloud_small(6, 32) <= 2; cloud_small(6, 33) <= 2; cloud_small(6, 34) <= 2; cloud_small(6, 35) <= 2; cloud_small(6, 36) <= 2; cloud_small(6, 37) <= 2; cloud_small(6, 38) <= 2; 
cloud_small(7, 0) <= 2; cloud_small(7, 1) <= 2; cloud_small(7, 2) <= 2; cloud_small(7, 3) <= 2; cloud_small(7, 4) <= 2; cloud_small(7, 5) <= 2; cloud_small(7, 6) <= 1; cloud_small(7, 7) <= 1; cloud_small(7, 8) <= 1; cloud_small(7, 9) <= 1; cloud_small(7, 10) <= 1; cloud_small(7, 11) <= 1; cloud_small(7, 12) <= 0; cloud_small(7, 13) <= 0; cloud_small(7, 14) <= 0; cloud_small(7, 15) <= 0; cloud_small(7, 16) <= 0; cloud_small(7, 17) <= 0; cloud_small(7, 18) <= 0; cloud_small(7, 19) <= 0; cloud_small(7, 20) <= 0; cloud_small(7, 21) <= 0; cloud_small(7, 22) <= 0; cloud_small(7, 23) <= 0; cloud_small(7, 24) <= 0; cloud_small(7, 25) <= 0; cloud_small(7, 26) <= 0; cloud_small(7, 27) <= 1; cloud_small(7, 28) <= 1; cloud_small(7, 29) <= 1; cloud_small(7, 30) <= 2; cloud_small(7, 31) <= 2; cloud_small(7, 32) <= 2; cloud_small(7, 33) <= 2; cloud_small(7, 34) <= 2; cloud_small(7, 35) <= 2; cloud_small(7, 36) <= 2; cloud_small(7, 37) <= 2; cloud_small(7, 38) <= 2; 
cloud_small(8, 0) <= 2; cloud_small(8, 1) <= 2; cloud_small(8, 2) <= 2; cloud_small(8, 3) <= 2; cloud_small(8, 4) <= 2; cloud_small(8, 5) <= 2; cloud_small(8, 6) <= 1; cloud_small(8, 7) <= 1; cloud_small(8, 8) <= 1; cloud_small(8, 9) <= 1; cloud_small(8, 10) <= 1; cloud_small(8, 11) <= 1; cloud_small(8, 12) <= 0; cloud_small(8, 13) <= 0; cloud_small(8, 14) <= 0; cloud_small(8, 15) <= 0; cloud_small(8, 16) <= 0; cloud_small(8, 17) <= 0; cloud_small(8, 18) <= 0; cloud_small(8, 19) <= 0; cloud_small(8, 20) <= 0; cloud_small(8, 21) <= 0; cloud_small(8, 22) <= 0; cloud_small(8, 23) <= 0; cloud_small(8, 24) <= 0; cloud_small(8, 25) <= 0; cloud_small(8, 26) <= 0; cloud_small(8, 27) <= 1; cloud_small(8, 28) <= 1; cloud_small(8, 29) <= 1; cloud_small(8, 30) <= 2; cloud_small(8, 31) <= 2; cloud_small(8, 32) <= 2; cloud_small(8, 33) <= 2; cloud_small(8, 34) <= 2; cloud_small(8, 35) <= 2; cloud_small(8, 36) <= 2; cloud_small(8, 37) <= 2; cloud_small(8, 38) <= 2; 
cloud_small(9, 0) <= 2; cloud_small(9, 1) <= 2; cloud_small(9, 2) <= 2; cloud_small(9, 3) <= 1; cloud_small(9, 4) <= 1; cloud_small(9, 5) <= 1; cloud_small(9, 6) <= 0; cloud_small(9, 7) <= 0; cloud_small(9, 8) <= 0; cloud_small(9, 9) <= 0; cloud_small(9, 10) <= 0; cloud_small(9, 11) <= 0; cloud_small(9, 12) <= 0; cloud_small(9, 13) <= 0; cloud_small(9, 14) <= 0; cloud_small(9, 15) <= 0; cloud_small(9, 16) <= 0; cloud_small(9, 17) <= 0; cloud_small(9, 18) <= 0; cloud_small(9, 19) <= 0; cloud_small(9, 20) <= 0; cloud_small(9, 21) <= 0; cloud_small(9, 22) <= 0; cloud_small(9, 23) <= 0; cloud_small(9, 24) <= 0; cloud_small(9, 25) <= 0; cloud_small(9, 26) <= 0; cloud_small(9, 27) <= 0; cloud_small(9, 28) <= 0; cloud_small(9, 29) <= 0; cloud_small(9, 30) <= 1; cloud_small(9, 31) <= 1; cloud_small(9, 32) <= 1; cloud_small(9, 33) <= 1; cloud_small(9, 34) <= 1; cloud_small(9, 35) <= 1; cloud_small(9, 36) <= 2; cloud_small(9, 37) <= 2; cloud_small(9, 38) <= 2; 
cloud_small(10, 0) <= 2; cloud_small(10, 1) <= 2; cloud_small(10, 2) <= 2; cloud_small(10, 3) <= 1; cloud_small(10, 4) <= 1; cloud_small(10, 5) <= 1; cloud_small(10, 6) <= 0; cloud_small(10, 7) <= 0; cloud_small(10, 8) <= 0; cloud_small(10, 9) <= 0; cloud_small(10, 10) <= 0; cloud_small(10, 11) <= 0; cloud_small(10, 12) <= 0; cloud_small(10, 13) <= 0; cloud_small(10, 14) <= 0; cloud_small(10, 15) <= 0; cloud_small(10, 16) <= 0; cloud_small(10, 17) <= 0; cloud_small(10, 18) <= 0; cloud_small(10, 19) <= 0; cloud_small(10, 20) <= 0; cloud_small(10, 21) <= 0; cloud_small(10, 22) <= 0; cloud_small(10, 23) <= 0; cloud_small(10, 24) <= 0; cloud_small(10, 25) <= 0; cloud_small(10, 26) <= 0; cloud_small(10, 27) <= 0; cloud_small(10, 28) <= 0; cloud_small(10, 29) <= 0; cloud_small(10, 30) <= 1; cloud_small(10, 31) <= 1; cloud_small(10, 32) <= 1; cloud_small(10, 33) <= 1; cloud_small(10, 34) <= 1; cloud_small(10, 35) <= 1; cloud_small(10, 36) <= 2; cloud_small(10, 37) <= 2; cloud_small(10, 38) <= 2; 
cloud_small(11, 0) <= 2; cloud_small(11, 1) <= 2; cloud_small(11, 2) <= 2; cloud_small(11, 3) <= 1; cloud_small(11, 4) <= 1; cloud_small(11, 5) <= 1; cloud_small(11, 6) <= 0; cloud_small(11, 7) <= 0; cloud_small(11, 8) <= 0; cloud_small(11, 9) <= 0; cloud_small(11, 10) <= 0; cloud_small(11, 11) <= 0; cloud_small(11, 12) <= 0; cloud_small(11, 13) <= 0; cloud_small(11, 14) <= 0; cloud_small(11, 15) <= 0; cloud_small(11, 16) <= 0; cloud_small(11, 17) <= 0; cloud_small(11, 18) <= 0; cloud_small(11, 19) <= 0; cloud_small(11, 20) <= 0; cloud_small(11, 21) <= 0; cloud_small(11, 22) <= 0; cloud_small(11, 23) <= 0; cloud_small(11, 24) <= 0; cloud_small(11, 25) <= 0; cloud_small(11, 26) <= 0; cloud_small(11, 27) <= 0; cloud_small(11, 28) <= 0; cloud_small(11, 29) <= 0; cloud_small(11, 30) <= 1; cloud_small(11, 31) <= 1; cloud_small(11, 32) <= 1; cloud_small(11, 33) <= 1; cloud_small(11, 34) <= 1; cloud_small(11, 35) <= 1; cloud_small(11, 36) <= 2; cloud_small(11, 37) <= 2; cloud_small(11, 38) <= 2; 
cloud_small(12, 0) <= 1; cloud_small(12, 1) <= 1; cloud_small(12, 2) <= 1; cloud_small(12, 3) <= 0; cloud_small(12, 4) <= 0; cloud_small(12, 5) <= 0; cloud_small(12, 6) <= 0; cloud_small(12, 7) <= 0; cloud_small(12, 8) <= 0; cloud_small(12, 9) <= 0; cloud_small(12, 10) <= 0; cloud_small(12, 11) <= 0; cloud_small(12, 12) <= 0; cloud_small(12, 13) <= 0; cloud_small(12, 14) <= 0; cloud_small(12, 15) <= 0; cloud_small(12, 16) <= 0; cloud_small(12, 17) <= 0; cloud_small(12, 18) <= 0; cloud_small(12, 19) <= 0; cloud_small(12, 20) <= 0; cloud_small(12, 21) <= 0; cloud_small(12, 22) <= 0; cloud_small(12, 23) <= 0; cloud_small(12, 24) <= 0; cloud_small(12, 25) <= 0; cloud_small(12, 26) <= 0; cloud_small(12, 27) <= 0; cloud_small(12, 28) <= 0; cloud_small(12, 29) <= 0; cloud_small(12, 30) <= 0; cloud_small(12, 31) <= 0; cloud_small(12, 32) <= 0; cloud_small(12, 33) <= 0; cloud_small(12, 34) <= 0; cloud_small(12, 35) <= 0; cloud_small(12, 36) <= 1; cloud_small(12, 37) <= 1; cloud_small(12, 38) <= 1; 
cloud_small(13, 0) <= 1; cloud_small(13, 1) <= 1; cloud_small(13, 2) <= 1; cloud_small(13, 3) <= 0; cloud_small(13, 4) <= 0; cloud_small(13, 5) <= 0; cloud_small(13, 6) <= 0; cloud_small(13, 7) <= 0; cloud_small(13, 8) <= 0; cloud_small(13, 9) <= 0; cloud_small(13, 10) <= 0; cloud_small(13, 11) <= 0; cloud_small(13, 12) <= 0; cloud_small(13, 13) <= 0; cloud_small(13, 14) <= 0; cloud_small(13, 15) <= 0; cloud_small(13, 16) <= 0; cloud_small(13, 17) <= 0; cloud_small(13, 18) <= 0; cloud_small(13, 19) <= 0; cloud_small(13, 20) <= 0; cloud_small(13, 21) <= 0; cloud_small(13, 22) <= 0; cloud_small(13, 23) <= 0; cloud_small(13, 24) <= 0; cloud_small(13, 25) <= 0; cloud_small(13, 26) <= 0; cloud_small(13, 27) <= 0; cloud_small(13, 28) <= 0; cloud_small(13, 29) <= 0; cloud_small(13, 30) <= 0; cloud_small(13, 31) <= 0; cloud_small(13, 32) <= 0; cloud_small(13, 33) <= 0; cloud_small(13, 34) <= 0; cloud_small(13, 35) <= 0; cloud_small(13, 36) <= 1; cloud_small(13, 37) <= 1; cloud_small(13, 38) <= 1; 
cloud_small(14, 0) <= 1; cloud_small(14, 1) <= 1; cloud_small(14, 2) <= 1; cloud_small(14, 3) <= 0; cloud_small(14, 4) <= 0; cloud_small(14, 5) <= 0; cloud_small(14, 6) <= 0; cloud_small(14, 7) <= 0; cloud_small(14, 8) <= 0; cloud_small(14, 9) <= 0; cloud_small(14, 10) <= 0; cloud_small(14, 11) <= 0; cloud_small(14, 12) <= 0; cloud_small(14, 13) <= 0; cloud_small(14, 14) <= 0; cloud_small(14, 15) <= 0; cloud_small(14, 16) <= 0; cloud_small(14, 17) <= 0; cloud_small(14, 18) <= 0; cloud_small(14, 19) <= 0; cloud_small(14, 20) <= 0; cloud_small(14, 21) <= 0; cloud_small(14, 22) <= 0; cloud_small(14, 23) <= 0; cloud_small(14, 24) <= 0; cloud_small(14, 25) <= 0; cloud_small(14, 26) <= 0; cloud_small(14, 27) <= 0; cloud_small(14, 28) <= 0; cloud_small(14, 29) <= 0; cloud_small(14, 30) <= 0; cloud_small(14, 31) <= 0; cloud_small(14, 32) <= 0; cloud_small(14, 33) <= 0; cloud_small(14, 34) <= 0; cloud_small(14, 35) <= 0; cloud_small(14, 36) <= 1; cloud_small(14, 37) <= 1; cloud_small(14, 38) <= 1; 
cloud_small(15, 0) <= 1; cloud_small(15, 1) <= 1; cloud_small(15, 2) <= 1; cloud_small(15, 3) <= 0; cloud_small(15, 4) <= 0; cloud_small(15, 5) <= 0; cloud_small(15, 6) <= 0; cloud_small(15, 7) <= 0; cloud_small(15, 8) <= 0; cloud_small(15, 9) <= 0; cloud_small(15, 10) <= 0; cloud_small(15, 11) <= 0; cloud_small(15, 12) <= 0; cloud_small(15, 13) <= 0; cloud_small(15, 14) <= 0; cloud_small(15, 15) <= 0; cloud_small(15, 16) <= 0; cloud_small(15, 17) <= 0; cloud_small(15, 18) <= 0; cloud_small(15, 19) <= 0; cloud_small(15, 20) <= 0; cloud_small(15, 21) <= 0; cloud_small(15, 22) <= 0; cloud_small(15, 23) <= 0; cloud_small(15, 24) <= 0; cloud_small(15, 25) <= 0; cloud_small(15, 26) <= 0; cloud_small(15, 27) <= 0; cloud_small(15, 28) <= 0; cloud_small(15, 29) <= 0; cloud_small(15, 30) <= 0; cloud_small(15, 31) <= 0; cloud_small(15, 32) <= 0; cloud_small(15, 33) <= 0; cloud_small(15, 34) <= 0; cloud_small(15, 35) <= 0; cloud_small(15, 36) <= 1; cloud_small(15, 37) <= 1; cloud_small(15, 38) <= 1; 
cloud_small(16, 0) <= 1; cloud_small(16, 1) <= 1; cloud_small(16, 2) <= 1; cloud_small(16, 3) <= 0; cloud_small(16, 4) <= 0; cloud_small(16, 5) <= 0; cloud_small(16, 6) <= 0; cloud_small(16, 7) <= 0; cloud_small(16, 8) <= 0; cloud_small(16, 9) <= 0; cloud_small(16, 10) <= 0; cloud_small(16, 11) <= 0; cloud_small(16, 12) <= 0; cloud_small(16, 13) <= 0; cloud_small(16, 14) <= 0; cloud_small(16, 15) <= 0; cloud_small(16, 16) <= 0; cloud_small(16, 17) <= 0; cloud_small(16, 18) <= 0; cloud_small(16, 19) <= 0; cloud_small(16, 20) <= 0; cloud_small(16, 21) <= 0; cloud_small(16, 22) <= 0; cloud_small(16, 23) <= 0; cloud_small(16, 24) <= 0; cloud_small(16, 25) <= 0; cloud_small(16, 26) <= 0; cloud_small(16, 27) <= 0; cloud_small(16, 28) <= 0; cloud_small(16, 29) <= 0; cloud_small(16, 30) <= 0; cloud_small(16, 31) <= 0; cloud_small(16, 32) <= 0; cloud_small(16, 33) <= 0; cloud_small(16, 34) <= 0; cloud_small(16, 35) <= 0; cloud_small(16, 36) <= 1; cloud_small(16, 37) <= 1; cloud_small(16, 38) <= 1; 
cloud_small(17, 0) <= 1; cloud_small(17, 1) <= 1; cloud_small(17, 2) <= 1; cloud_small(17, 3) <= 0; cloud_small(17, 4) <= 0; cloud_small(17, 5) <= 0; cloud_small(17, 6) <= 0; cloud_small(17, 7) <= 0; cloud_small(17, 8) <= 0; cloud_small(17, 9) <= 0; cloud_small(17, 10) <= 0; cloud_small(17, 11) <= 0; cloud_small(17, 12) <= 0; cloud_small(17, 13) <= 0; cloud_small(17, 14) <= 0; cloud_small(17, 15) <= 0; cloud_small(17, 16) <= 0; cloud_small(17, 17) <= 0; cloud_small(17, 18) <= 0; cloud_small(17, 19) <= 0; cloud_small(17, 20) <= 0; cloud_small(17, 21) <= 0; cloud_small(17, 22) <= 0; cloud_small(17, 23) <= 0; cloud_small(17, 24) <= 0; cloud_small(17, 25) <= 0; cloud_small(17, 26) <= 0; cloud_small(17, 27) <= 0; cloud_small(17, 28) <= 0; cloud_small(17, 29) <= 0; cloud_small(17, 30) <= 0; cloud_small(17, 31) <= 0; cloud_small(17, 32) <= 0; cloud_small(17, 33) <= 0; cloud_small(17, 34) <= 0; cloud_small(17, 35) <= 0; cloud_small(17, 36) <= 1; cloud_small(17, 37) <= 1; cloud_small(17, 38) <= 1; 
cloud_small(18, 0) <= 1; cloud_small(18, 1) <= 1; cloud_small(18, 2) <= 1; cloud_small(18, 3) <= 0; cloud_small(18, 4) <= 0; cloud_small(18, 5) <= 0; cloud_small(18, 6) <= 0; cloud_small(18, 7) <= 0; cloud_small(18, 8) <= 0; cloud_small(18, 9) <= 0; cloud_small(18, 10) <= 0; cloud_small(18, 11) <= 0; cloud_small(18, 12) <= 0; cloud_small(18, 13) <= 0; cloud_small(18, 14) <= 0; cloud_small(18, 15) <= 0; cloud_small(18, 16) <= 0; cloud_small(18, 17) <= 0; cloud_small(18, 18) <= 0; cloud_small(18, 19) <= 0; cloud_small(18, 20) <= 0; cloud_small(18, 21) <= 0; cloud_small(18, 22) <= 0; cloud_small(18, 23) <= 0; cloud_small(18, 24) <= 0; cloud_small(18, 25) <= 0; cloud_small(18, 26) <= 0; cloud_small(18, 27) <= 0; cloud_small(18, 28) <= 0; cloud_small(18, 29) <= 0; cloud_small(18, 30) <= 0; cloud_small(18, 31) <= 0; cloud_small(18, 32) <= 0; cloud_small(18, 33) <= 0; cloud_small(18, 34) <= 0; cloud_small(18, 35) <= 0; cloud_small(18, 36) <= 1; cloud_small(18, 37) <= 1; cloud_small(18, 38) <= 1; 
cloud_small(19, 0) <= 1; cloud_small(19, 1) <= 1; cloud_small(19, 2) <= 1; cloud_small(19, 3) <= 0; cloud_small(19, 4) <= 0; cloud_small(19, 5) <= 0; cloud_small(19, 6) <= 0; cloud_small(19, 7) <= 0; cloud_small(19, 8) <= 0; cloud_small(19, 9) <= 0; cloud_small(19, 10) <= 0; cloud_small(19, 11) <= 0; cloud_small(19, 12) <= 0; cloud_small(19, 13) <= 0; cloud_small(19, 14) <= 0; cloud_small(19, 15) <= 0; cloud_small(19, 16) <= 0; cloud_small(19, 17) <= 0; cloud_small(19, 18) <= 0; cloud_small(19, 19) <= 0; cloud_small(19, 20) <= 0; cloud_small(19, 21) <= 0; cloud_small(19, 22) <= 0; cloud_small(19, 23) <= 0; cloud_small(19, 24) <= 0; cloud_small(19, 25) <= 0; cloud_small(19, 26) <= 0; cloud_small(19, 27) <= 0; cloud_small(19, 28) <= 0; cloud_small(19, 29) <= 0; cloud_small(19, 30) <= 0; cloud_small(19, 31) <= 0; cloud_small(19, 32) <= 0; cloud_small(19, 33) <= 0; cloud_small(19, 34) <= 0; cloud_small(19, 35) <= 0; cloud_small(19, 36) <= 1; cloud_small(19, 37) <= 1; cloud_small(19, 38) <= 1; 
cloud_small(20, 0) <= 1; cloud_small(20, 1) <= 1; cloud_small(20, 2) <= 1; cloud_small(20, 3) <= 0; cloud_small(20, 4) <= 0; cloud_small(20, 5) <= 0; cloud_small(20, 6) <= 0; cloud_small(20, 7) <= 0; cloud_small(20, 8) <= 0; cloud_small(20, 9) <= 0; cloud_small(20, 10) <= 0; cloud_small(20, 11) <= 0; cloud_small(20, 12) <= 0; cloud_small(20, 13) <= 0; cloud_small(20, 14) <= 0; cloud_small(20, 15) <= 0; cloud_small(20, 16) <= 0; cloud_small(20, 17) <= 0; cloud_small(20, 18) <= 0; cloud_small(20, 19) <= 0; cloud_small(20, 20) <= 0; cloud_small(20, 21) <= 0; cloud_small(20, 22) <= 0; cloud_small(20, 23) <= 0; cloud_small(20, 24) <= 0; cloud_small(20, 25) <= 0; cloud_small(20, 26) <= 0; cloud_small(20, 27) <= 0; cloud_small(20, 28) <= 0; cloud_small(20, 29) <= 0; cloud_small(20, 30) <= 0; cloud_small(20, 31) <= 0; cloud_small(20, 32) <= 0; cloud_small(20, 33) <= 0; cloud_small(20, 34) <= 0; cloud_small(20, 35) <= 0; cloud_small(20, 36) <= 1; cloud_small(20, 37) <= 1; cloud_small(20, 38) <= 1; 
cloud_small(21, 0) <= 2; cloud_small(21, 1) <= 2; cloud_small(21, 2) <= 2; cloud_small(21, 3) <= 1; cloud_small(21, 4) <= 1; cloud_small(21, 5) <= 1; cloud_small(21, 6) <= 0; cloud_small(21, 7) <= 0; cloud_small(21, 8) <= 0; cloud_small(21, 9) <= 0; cloud_small(21, 10) <= 0; cloud_small(21, 11) <= 0; cloud_small(21, 12) <= 0; cloud_small(21, 13) <= 0; cloud_small(21, 14) <= 0; cloud_small(21, 15) <= 0; cloud_small(21, 16) <= 0; cloud_small(21, 17) <= 0; cloud_small(21, 18) <= 0; cloud_small(21, 19) <= 0; cloud_small(21, 20) <= 0; cloud_small(21, 21) <= 0; cloud_small(21, 22) <= 0; cloud_small(21, 23) <= 0; cloud_small(21, 24) <= 0; cloud_small(21, 25) <= 0; cloud_small(21, 26) <= 0; cloud_small(21, 27) <= 0; cloud_small(21, 28) <= 0; cloud_small(21, 29) <= 0; cloud_small(21, 30) <= 0; cloud_small(21, 31) <= 0; cloud_small(21, 32) <= 0; cloud_small(21, 33) <= 1; cloud_small(21, 34) <= 1; cloud_small(21, 35) <= 1; cloud_small(21, 36) <= 2; cloud_small(21, 37) <= 2; cloud_small(21, 38) <= 2; 
cloud_small(22, 0) <= 2; cloud_small(22, 1) <= 2; cloud_small(22, 2) <= 2; cloud_small(22, 3) <= 1; cloud_small(22, 4) <= 1; cloud_small(22, 5) <= 1; cloud_small(22, 6) <= 0; cloud_small(22, 7) <= 0; cloud_small(22, 8) <= 0; cloud_small(22, 9) <= 0; cloud_small(22, 10) <= 0; cloud_small(22, 11) <= 0; cloud_small(22, 12) <= 0; cloud_small(22, 13) <= 0; cloud_small(22, 14) <= 0; cloud_small(22, 15) <= 0; cloud_small(22, 16) <= 0; cloud_small(22, 17) <= 0; cloud_small(22, 18) <= 0; cloud_small(22, 19) <= 0; cloud_small(22, 20) <= 0; cloud_small(22, 21) <= 0; cloud_small(22, 22) <= 0; cloud_small(22, 23) <= 0; cloud_small(22, 24) <= 0; cloud_small(22, 25) <= 0; cloud_small(22, 26) <= 0; cloud_small(22, 27) <= 0; cloud_small(22, 28) <= 0; cloud_small(22, 29) <= 0; cloud_small(22, 30) <= 0; cloud_small(22, 31) <= 0; cloud_small(22, 32) <= 0; cloud_small(22, 33) <= 1; cloud_small(22, 34) <= 1; cloud_small(22, 35) <= 1; cloud_small(22, 36) <= 2; cloud_small(22, 37) <= 2; cloud_small(22, 38) <= 2; 
cloud_small(23, 0) <= 2; cloud_small(23, 1) <= 2; cloud_small(23, 2) <= 2; cloud_small(23, 3) <= 1; cloud_small(23, 4) <= 1; cloud_small(23, 5) <= 1; cloud_small(23, 6) <= 0; cloud_small(23, 7) <= 0; cloud_small(23, 8) <= 0; cloud_small(23, 9) <= 0; cloud_small(23, 10) <= 0; cloud_small(23, 11) <= 0; cloud_small(23, 12) <= 0; cloud_small(23, 13) <= 0; cloud_small(23, 14) <= 0; cloud_small(23, 15) <= 0; cloud_small(23, 16) <= 0; cloud_small(23, 17) <= 0; cloud_small(23, 18) <= 0; cloud_small(23, 19) <= 0; cloud_small(23, 20) <= 0; cloud_small(23, 21) <= 0; cloud_small(23, 22) <= 0; cloud_small(23, 23) <= 0; cloud_small(23, 24) <= 0; cloud_small(23, 25) <= 0; cloud_small(23, 26) <= 0; cloud_small(23, 27) <= 0; cloud_small(23, 28) <= 0; cloud_small(23, 29) <= 0; cloud_small(23, 30) <= 0; cloud_small(23, 31) <= 0; cloud_small(23, 32) <= 0; cloud_small(23, 33) <= 1; cloud_small(23, 34) <= 1; cloud_small(23, 35) <= 1; cloud_small(23, 36) <= 2; cloud_small(23, 37) <= 2; cloud_small(23, 38) <= 2; 
cloud_small(24, 0) <= 2; cloud_small(24, 1) <= 2; cloud_small(24, 2) <= 2; cloud_small(24, 3) <= 2; cloud_small(24, 4) <= 2; cloud_small(24, 5) <= 2; cloud_small(24, 6) <= 1; cloud_small(24, 7) <= 1; cloud_small(24, 8) <= 1; cloud_small(24, 9) <= 1; cloud_small(24, 10) <= 1; cloud_small(24, 11) <= 1; cloud_small(24, 12) <= 1; cloud_small(24, 13) <= 1; cloud_small(24, 14) <= 1; cloud_small(24, 15) <= 1; cloud_small(24, 16) <= 1; cloud_small(24, 17) <= 1; cloud_small(24, 18) <= 1; cloud_small(24, 19) <= 1; cloud_small(24, 20) <= 1; cloud_small(24, 21) <= 1; cloud_small(24, 22) <= 1; cloud_small(24, 23) <= 1; cloud_small(24, 24) <= 1; cloud_small(24, 25) <= 1; cloud_small(24, 26) <= 1; cloud_small(24, 27) <= 1; cloud_small(24, 28) <= 1; cloud_small(24, 29) <= 1; cloud_small(24, 30) <= 1; cloud_small(24, 31) <= 1; cloud_small(24, 32) <= 1; cloud_small(24, 33) <= 2; cloud_small(24, 34) <= 2; cloud_small(24, 35) <= 2; cloud_small(24, 36) <= 2; cloud_small(24, 37) <= 2; cloud_small(24, 38) <= 2; 
cloud_small(25, 0) <= 2; cloud_small(25, 1) <= 2; cloud_small(25, 2) <= 2; cloud_small(25, 3) <= 2; cloud_small(25, 4) <= 2; cloud_small(25, 5) <= 2; cloud_small(25, 6) <= 1; cloud_small(25, 7) <= 1; cloud_small(25, 8) <= 1; cloud_small(25, 9) <= 1; cloud_small(25, 10) <= 1; cloud_small(25, 11) <= 1; cloud_small(25, 12) <= 1; cloud_small(25, 13) <= 1; cloud_small(25, 14) <= 1; cloud_small(25, 15) <= 1; cloud_small(25, 16) <= 1; cloud_small(25, 17) <= 1; cloud_small(25, 18) <= 1; cloud_small(25, 19) <= 1; cloud_small(25, 20) <= 1; cloud_small(25, 21) <= 1; cloud_small(25, 22) <= 1; cloud_small(25, 23) <= 1; cloud_small(25, 24) <= 1; cloud_small(25, 25) <= 1; cloud_small(25, 26) <= 1; cloud_small(25, 27) <= 1; cloud_small(25, 28) <= 1; cloud_small(25, 29) <= 1; cloud_small(25, 30) <= 1; cloud_small(25, 31) <= 1; cloud_small(25, 32) <= 1; cloud_small(25, 33) <= 2; cloud_small(25, 34) <= 2; cloud_small(25, 35) <= 2; cloud_small(25, 36) <= 2; cloud_small(25, 37) <= 2; cloud_small(25, 38) <= 2; 
cloud_small(26, 0) <= 2; cloud_small(26, 1) <= 2; cloud_small(26, 2) <= 2; cloud_small(26, 3) <= 2; cloud_small(26, 4) <= 2; cloud_small(26, 5) <= 2; cloud_small(26, 6) <= 1; cloud_small(26, 7) <= 1; cloud_small(26, 8) <= 1; cloud_small(26, 9) <= 1; cloud_small(26, 10) <= 1; cloud_small(26, 11) <= 1; cloud_small(26, 12) <= 1; cloud_small(26, 13) <= 1; cloud_small(26, 14) <= 1; cloud_small(26, 15) <= 1; cloud_small(26, 16) <= 1; cloud_small(26, 17) <= 1; cloud_small(26, 18) <= 1; cloud_small(26, 19) <= 1; cloud_small(26, 20) <= 1; cloud_small(26, 21) <= 1; cloud_small(26, 22) <= 1; cloud_small(26, 23) <= 1; cloud_small(26, 24) <= 1; cloud_small(26, 25) <= 1; cloud_small(26, 26) <= 1; cloud_small(26, 27) <= 1; cloud_small(26, 28) <= 1; cloud_small(26, 29) <= 1; cloud_small(26, 30) <= 1; cloud_small(26, 31) <= 1; cloud_small(26, 32) <= 1; cloud_small(26, 33) <= 2; cloud_small(26, 34) <= 2; cloud_small(26, 35) <= 2; cloud_small(26, 36) <= 2; cloud_small(26, 37) <= 2; cloud_small(26, 38) <= 2; 

cloud_xl(0, 0) <= 2; cloud_xl(0, 1) <= 2; cloud_xl(0, 2) <= 2; cloud_xl(0, 3) <= 2; cloud_xl(0, 4) <= 2; cloud_xl(0, 5) <= 2; cloud_xl(0, 6) <= 2; cloud_xl(0, 7) <= 2; cloud_xl(0, 8) <= 2; cloud_xl(0, 9) <= 2; cloud_xl(0, 10) <= 2; cloud_xl(0, 11) <= 2; cloud_xl(0, 12) <= 2; cloud_xl(0, 13) <= 2; cloud_xl(0, 14) <= 2; cloud_xl(0, 15) <= 2; cloud_xl(0, 16) <= 2; cloud_xl(0, 17) <= 2; cloud_xl(0, 18) <= 2; cloud_xl(0, 19) <= 2; cloud_xl(0, 20) <= 2; cloud_xl(0, 21) <= 2; cloud_xl(0, 22) <= 2; cloud_xl(0, 23) <= 2; cloud_xl(0, 24) <= 2; cloud_xl(0, 25) <= 2; cloud_xl(0, 26) <= 2; cloud_xl(0, 27) <= 2; cloud_xl(0, 28) <= 2; cloud_xl(0, 29) <= 2; cloud_xl(0, 30) <= 1; cloud_xl(0, 31) <= 1; cloud_xl(0, 32) <= 1; cloud_xl(0, 33) <= 1; cloud_xl(0, 34) <= 1; cloud_xl(0, 35) <= 1; cloud_xl(0, 36) <= 1; cloud_xl(0, 37) <= 1; cloud_xl(0, 38) <= 1; cloud_xl(0, 39) <= 1; cloud_xl(0, 40) <= 1; cloud_xl(0, 41) <= 1; cloud_xl(0, 42) <= 1; cloud_xl(0, 43) <= 1; cloud_xl(0, 44) <= 1; cloud_xl(0, 45) <= 1; cloud_xl(0, 46) <= 1; cloud_xl(0, 47) <= 1; cloud_xl(0, 48) <= 2; cloud_xl(0, 49) <= 2; cloud_xl(0, 50) <= 2; cloud_xl(0, 51) <= 2; cloud_xl(0, 52) <= 2; cloud_xl(0, 53) <= 2; cloud_xl(0, 54) <= 2; cloud_xl(0, 55) <= 2; cloud_xl(0, 56) <= 2; cloud_xl(0, 57) <= 2; cloud_xl(0, 58) <= 2; cloud_xl(0, 59) <= 2; cloud_xl(0, 60) <= 2; cloud_xl(0, 61) <= 2; cloud_xl(0, 62) <= 2; cloud_xl(0, 63) <= 2; cloud_xl(0, 64) <= 2; cloud_xl(0, 65) <= 2; cloud_xl(0, 66) <= 2; cloud_xl(0, 67) <= 2; cloud_xl(0, 68) <= 2; cloud_xl(0, 69) <= 2; cloud_xl(0, 70) <= 2; cloud_xl(0, 71) <= 2; cloud_xl(0, 72) <= 2; cloud_xl(0, 73) <= 2; cloud_xl(0, 74) <= 2; cloud_xl(0, 75) <= 2; cloud_xl(0, 76) <= 2; cloud_xl(0, 77) <= 2; 
cloud_xl(1, 0) <= 2; cloud_xl(1, 1) <= 2; cloud_xl(1, 2) <= 2; cloud_xl(1, 3) <= 2; cloud_xl(1, 4) <= 2; cloud_xl(1, 5) <= 2; cloud_xl(1, 6) <= 2; cloud_xl(1, 7) <= 2; cloud_xl(1, 8) <= 2; cloud_xl(1, 9) <= 2; cloud_xl(1, 10) <= 2; cloud_xl(1, 11) <= 2; cloud_xl(1, 12) <= 2; cloud_xl(1, 13) <= 2; cloud_xl(1, 14) <= 2; cloud_xl(1, 15) <= 2; cloud_xl(1, 16) <= 2; cloud_xl(1, 17) <= 2; cloud_xl(1, 18) <= 2; cloud_xl(1, 19) <= 2; cloud_xl(1, 20) <= 2; cloud_xl(1, 21) <= 2; cloud_xl(1, 22) <= 2; cloud_xl(1, 23) <= 2; cloud_xl(1, 24) <= 2; cloud_xl(1, 25) <= 2; cloud_xl(1, 26) <= 2; cloud_xl(1, 27) <= 2; cloud_xl(1, 28) <= 2; cloud_xl(1, 29) <= 2; cloud_xl(1, 30) <= 1; cloud_xl(1, 31) <= 1; cloud_xl(1, 32) <= 1; cloud_xl(1, 33) <= 1; cloud_xl(1, 34) <= 1; cloud_xl(1, 35) <= 1; cloud_xl(1, 36) <= 1; cloud_xl(1, 37) <= 1; cloud_xl(1, 38) <= 1; cloud_xl(1, 39) <= 1; cloud_xl(1, 40) <= 1; cloud_xl(1, 41) <= 1; cloud_xl(1, 42) <= 1; cloud_xl(1, 43) <= 1; cloud_xl(1, 44) <= 1; cloud_xl(1, 45) <= 1; cloud_xl(1, 46) <= 1; cloud_xl(1, 47) <= 1; cloud_xl(1, 48) <= 2; cloud_xl(1, 49) <= 2; cloud_xl(1, 50) <= 2; cloud_xl(1, 51) <= 2; cloud_xl(1, 52) <= 2; cloud_xl(1, 53) <= 2; cloud_xl(1, 54) <= 2; cloud_xl(1, 55) <= 2; cloud_xl(1, 56) <= 2; cloud_xl(1, 57) <= 2; cloud_xl(1, 58) <= 2; cloud_xl(1, 59) <= 2; cloud_xl(1, 60) <= 2; cloud_xl(1, 61) <= 2; cloud_xl(1, 62) <= 2; cloud_xl(1, 63) <= 2; cloud_xl(1, 64) <= 2; cloud_xl(1, 65) <= 2; cloud_xl(1, 66) <= 2; cloud_xl(1, 67) <= 2; cloud_xl(1, 68) <= 2; cloud_xl(1, 69) <= 2; cloud_xl(1, 70) <= 2; cloud_xl(1, 71) <= 2; cloud_xl(1, 72) <= 2; cloud_xl(1, 73) <= 2; cloud_xl(1, 74) <= 2; cloud_xl(1, 75) <= 2; cloud_xl(1, 76) <= 2; cloud_xl(1, 77) <= 2; 
cloud_xl(2, 0) <= 2; cloud_xl(2, 1) <= 2; cloud_xl(2, 2) <= 2; cloud_xl(2, 3) <= 2; cloud_xl(2, 4) <= 2; cloud_xl(2, 5) <= 2; cloud_xl(2, 6) <= 2; cloud_xl(2, 7) <= 2; cloud_xl(2, 8) <= 2; cloud_xl(2, 9) <= 2; cloud_xl(2, 10) <= 2; cloud_xl(2, 11) <= 2; cloud_xl(2, 12) <= 2; cloud_xl(2, 13) <= 2; cloud_xl(2, 14) <= 2; cloud_xl(2, 15) <= 2; cloud_xl(2, 16) <= 2; cloud_xl(2, 17) <= 2; cloud_xl(2, 18) <= 2; cloud_xl(2, 19) <= 2; cloud_xl(2, 20) <= 2; cloud_xl(2, 21) <= 2; cloud_xl(2, 22) <= 2; cloud_xl(2, 23) <= 2; cloud_xl(2, 24) <= 2; cloud_xl(2, 25) <= 2; cloud_xl(2, 26) <= 2; cloud_xl(2, 27) <= 2; cloud_xl(2, 28) <= 2; cloud_xl(2, 29) <= 2; cloud_xl(2, 30) <= 1; cloud_xl(2, 31) <= 1; cloud_xl(2, 32) <= 1; cloud_xl(2, 33) <= 1; cloud_xl(2, 34) <= 1; cloud_xl(2, 35) <= 1; cloud_xl(2, 36) <= 1; cloud_xl(2, 37) <= 1; cloud_xl(2, 38) <= 1; cloud_xl(2, 39) <= 1; cloud_xl(2, 40) <= 1; cloud_xl(2, 41) <= 1; cloud_xl(2, 42) <= 1; cloud_xl(2, 43) <= 1; cloud_xl(2, 44) <= 1; cloud_xl(2, 45) <= 1; cloud_xl(2, 46) <= 1; cloud_xl(2, 47) <= 1; cloud_xl(2, 48) <= 2; cloud_xl(2, 49) <= 2; cloud_xl(2, 50) <= 2; cloud_xl(2, 51) <= 2; cloud_xl(2, 52) <= 2; cloud_xl(2, 53) <= 2; cloud_xl(2, 54) <= 2; cloud_xl(2, 55) <= 2; cloud_xl(2, 56) <= 2; cloud_xl(2, 57) <= 2; cloud_xl(2, 58) <= 2; cloud_xl(2, 59) <= 2; cloud_xl(2, 60) <= 2; cloud_xl(2, 61) <= 2; cloud_xl(2, 62) <= 2; cloud_xl(2, 63) <= 2; cloud_xl(2, 64) <= 2; cloud_xl(2, 65) <= 2; cloud_xl(2, 66) <= 2; cloud_xl(2, 67) <= 2; cloud_xl(2, 68) <= 2; cloud_xl(2, 69) <= 2; cloud_xl(2, 70) <= 2; cloud_xl(2, 71) <= 2; cloud_xl(2, 72) <= 2; cloud_xl(2, 73) <= 2; cloud_xl(2, 74) <= 2; cloud_xl(2, 75) <= 2; cloud_xl(2, 76) <= 2; cloud_xl(2, 77) <= 2; 
cloud_xl(3, 0) <= 2; cloud_xl(3, 1) <= 2; cloud_xl(3, 2) <= 2; cloud_xl(3, 3) <= 2; cloud_xl(3, 4) <= 2; cloud_xl(3, 5) <= 2; cloud_xl(3, 6) <= 2; cloud_xl(3, 7) <= 2; cloud_xl(3, 8) <= 2; cloud_xl(3, 9) <= 2; cloud_xl(3, 10) <= 2; cloud_xl(3, 11) <= 2; cloud_xl(3, 12) <= 2; cloud_xl(3, 13) <= 2; cloud_xl(3, 14) <= 2; cloud_xl(3, 15) <= 2; cloud_xl(3, 16) <= 2; cloud_xl(3, 17) <= 2; cloud_xl(3, 18) <= 2; cloud_xl(3, 19) <= 2; cloud_xl(3, 20) <= 2; cloud_xl(3, 21) <= 2; cloud_xl(3, 22) <= 2; cloud_xl(3, 23) <= 2; cloud_xl(3, 24) <= 2; cloud_xl(3, 25) <= 2; cloud_xl(3, 26) <= 2; cloud_xl(3, 27) <= 2; cloud_xl(3, 28) <= 2; cloud_xl(3, 29) <= 2; cloud_xl(3, 30) <= 1; cloud_xl(3, 31) <= 1; cloud_xl(3, 32) <= 1; cloud_xl(3, 33) <= 1; cloud_xl(3, 34) <= 1; cloud_xl(3, 35) <= 1; cloud_xl(3, 36) <= 1; cloud_xl(3, 37) <= 1; cloud_xl(3, 38) <= 1; cloud_xl(3, 39) <= 1; cloud_xl(3, 40) <= 1; cloud_xl(3, 41) <= 1; cloud_xl(3, 42) <= 1; cloud_xl(3, 43) <= 1; cloud_xl(3, 44) <= 1; cloud_xl(3, 45) <= 1; cloud_xl(3, 46) <= 1; cloud_xl(3, 47) <= 1; cloud_xl(3, 48) <= 2; cloud_xl(3, 49) <= 2; cloud_xl(3, 50) <= 2; cloud_xl(3, 51) <= 2; cloud_xl(3, 52) <= 2; cloud_xl(3, 53) <= 2; cloud_xl(3, 54) <= 2; cloud_xl(3, 55) <= 2; cloud_xl(3, 56) <= 2; cloud_xl(3, 57) <= 2; cloud_xl(3, 58) <= 2; cloud_xl(3, 59) <= 2; cloud_xl(3, 60) <= 2; cloud_xl(3, 61) <= 2; cloud_xl(3, 62) <= 2; cloud_xl(3, 63) <= 2; cloud_xl(3, 64) <= 2; cloud_xl(3, 65) <= 2; cloud_xl(3, 66) <= 2; cloud_xl(3, 67) <= 2; cloud_xl(3, 68) <= 2; cloud_xl(3, 69) <= 2; cloud_xl(3, 70) <= 2; cloud_xl(3, 71) <= 2; cloud_xl(3, 72) <= 2; cloud_xl(3, 73) <= 2; cloud_xl(3, 74) <= 2; cloud_xl(3, 75) <= 2; cloud_xl(3, 76) <= 2; cloud_xl(3, 77) <= 2; 
cloud_xl(4, 0) <= 2; cloud_xl(4, 1) <= 2; cloud_xl(4, 2) <= 2; cloud_xl(4, 3) <= 2; cloud_xl(4, 4) <= 2; cloud_xl(4, 5) <= 2; cloud_xl(4, 6) <= 2; cloud_xl(4, 7) <= 2; cloud_xl(4, 8) <= 2; cloud_xl(4, 9) <= 2; cloud_xl(4, 10) <= 2; cloud_xl(4, 11) <= 2; cloud_xl(4, 12) <= 2; cloud_xl(4, 13) <= 2; cloud_xl(4, 14) <= 2; cloud_xl(4, 15) <= 2; cloud_xl(4, 16) <= 2; cloud_xl(4, 17) <= 2; cloud_xl(4, 18) <= 2; cloud_xl(4, 19) <= 2; cloud_xl(4, 20) <= 2; cloud_xl(4, 21) <= 2; cloud_xl(4, 22) <= 2; cloud_xl(4, 23) <= 2; cloud_xl(4, 24) <= 2; cloud_xl(4, 25) <= 2; cloud_xl(4, 26) <= 2; cloud_xl(4, 27) <= 2; cloud_xl(4, 28) <= 2; cloud_xl(4, 29) <= 2; cloud_xl(4, 30) <= 1; cloud_xl(4, 31) <= 1; cloud_xl(4, 32) <= 1; cloud_xl(4, 33) <= 1; cloud_xl(4, 34) <= 1; cloud_xl(4, 35) <= 1; cloud_xl(4, 36) <= 1; cloud_xl(4, 37) <= 1; cloud_xl(4, 38) <= 1; cloud_xl(4, 39) <= 1; cloud_xl(4, 40) <= 1; cloud_xl(4, 41) <= 1; cloud_xl(4, 42) <= 1; cloud_xl(4, 43) <= 1; cloud_xl(4, 44) <= 1; cloud_xl(4, 45) <= 1; cloud_xl(4, 46) <= 1; cloud_xl(4, 47) <= 1; cloud_xl(4, 48) <= 2; cloud_xl(4, 49) <= 2; cloud_xl(4, 50) <= 2; cloud_xl(4, 51) <= 2; cloud_xl(4, 52) <= 2; cloud_xl(4, 53) <= 2; cloud_xl(4, 54) <= 2; cloud_xl(4, 55) <= 2; cloud_xl(4, 56) <= 2; cloud_xl(4, 57) <= 2; cloud_xl(4, 58) <= 2; cloud_xl(4, 59) <= 2; cloud_xl(4, 60) <= 2; cloud_xl(4, 61) <= 2; cloud_xl(4, 62) <= 2; cloud_xl(4, 63) <= 2; cloud_xl(4, 64) <= 2; cloud_xl(4, 65) <= 2; cloud_xl(4, 66) <= 2; cloud_xl(4, 67) <= 2; cloud_xl(4, 68) <= 2; cloud_xl(4, 69) <= 2; cloud_xl(4, 70) <= 2; cloud_xl(4, 71) <= 2; cloud_xl(4, 72) <= 2; cloud_xl(4, 73) <= 2; cloud_xl(4, 74) <= 2; cloud_xl(4, 75) <= 2; cloud_xl(4, 76) <= 2; cloud_xl(4, 77) <= 2; 
cloud_xl(5, 0) <= 2; cloud_xl(5, 1) <= 2; cloud_xl(5, 2) <= 2; cloud_xl(5, 3) <= 2; cloud_xl(5, 4) <= 2; cloud_xl(5, 5) <= 2; cloud_xl(5, 6) <= 2; cloud_xl(5, 7) <= 2; cloud_xl(5, 8) <= 2; cloud_xl(5, 9) <= 2; cloud_xl(5, 10) <= 2; cloud_xl(5, 11) <= 2; cloud_xl(5, 12) <= 2; cloud_xl(5, 13) <= 2; cloud_xl(5, 14) <= 2; cloud_xl(5, 15) <= 2; cloud_xl(5, 16) <= 2; cloud_xl(5, 17) <= 2; cloud_xl(5, 18) <= 2; cloud_xl(5, 19) <= 2; cloud_xl(5, 20) <= 2; cloud_xl(5, 21) <= 2; cloud_xl(5, 22) <= 2; cloud_xl(5, 23) <= 2; cloud_xl(5, 24) <= 2; cloud_xl(5, 25) <= 2; cloud_xl(5, 26) <= 2; cloud_xl(5, 27) <= 2; cloud_xl(5, 28) <= 2; cloud_xl(5, 29) <= 2; cloud_xl(5, 30) <= 1; cloud_xl(5, 31) <= 1; cloud_xl(5, 32) <= 1; cloud_xl(5, 33) <= 1; cloud_xl(5, 34) <= 1; cloud_xl(5, 35) <= 1; cloud_xl(5, 36) <= 1; cloud_xl(5, 37) <= 1; cloud_xl(5, 38) <= 1; cloud_xl(5, 39) <= 1; cloud_xl(5, 40) <= 1; cloud_xl(5, 41) <= 1; cloud_xl(5, 42) <= 1; cloud_xl(5, 43) <= 1; cloud_xl(5, 44) <= 1; cloud_xl(5, 45) <= 1; cloud_xl(5, 46) <= 1; cloud_xl(5, 47) <= 1; cloud_xl(5, 48) <= 2; cloud_xl(5, 49) <= 2; cloud_xl(5, 50) <= 2; cloud_xl(5, 51) <= 2; cloud_xl(5, 52) <= 2; cloud_xl(5, 53) <= 2; cloud_xl(5, 54) <= 2; cloud_xl(5, 55) <= 2; cloud_xl(5, 56) <= 2; cloud_xl(5, 57) <= 2; cloud_xl(5, 58) <= 2; cloud_xl(5, 59) <= 2; cloud_xl(5, 60) <= 2; cloud_xl(5, 61) <= 2; cloud_xl(5, 62) <= 2; cloud_xl(5, 63) <= 2; cloud_xl(5, 64) <= 2; cloud_xl(5, 65) <= 2; cloud_xl(5, 66) <= 2; cloud_xl(5, 67) <= 2; cloud_xl(5, 68) <= 2; cloud_xl(5, 69) <= 2; cloud_xl(5, 70) <= 2; cloud_xl(5, 71) <= 2; cloud_xl(5, 72) <= 2; cloud_xl(5, 73) <= 2; cloud_xl(5, 74) <= 2; cloud_xl(5, 75) <= 2; cloud_xl(5, 76) <= 2; cloud_xl(5, 77) <= 2; 
cloud_xl(6, 0) <= 2; cloud_xl(6, 1) <= 2; cloud_xl(6, 2) <= 2; cloud_xl(6, 3) <= 2; cloud_xl(6, 4) <= 2; cloud_xl(6, 5) <= 2; cloud_xl(6, 6) <= 2; cloud_xl(6, 7) <= 2; cloud_xl(6, 8) <= 2; cloud_xl(6, 9) <= 2; cloud_xl(6, 10) <= 2; cloud_xl(6, 11) <= 2; cloud_xl(6, 12) <= 2; cloud_xl(6, 13) <= 2; cloud_xl(6, 14) <= 2; cloud_xl(6, 15) <= 2; cloud_xl(6, 16) <= 2; cloud_xl(6, 17) <= 2; cloud_xl(6, 18) <= 2; cloud_xl(6, 19) <= 2; cloud_xl(6, 20) <= 2; cloud_xl(6, 21) <= 2; cloud_xl(6, 22) <= 2; cloud_xl(6, 23) <= 2; cloud_xl(6, 24) <= 1; cloud_xl(6, 25) <= 1; cloud_xl(6, 26) <= 1; cloud_xl(6, 27) <= 1; cloud_xl(6, 28) <= 1; cloud_xl(6, 29) <= 1; cloud_xl(6, 30) <= 0; cloud_xl(6, 31) <= 0; cloud_xl(6, 32) <= 0; cloud_xl(6, 33) <= 0; cloud_xl(6, 34) <= 0; cloud_xl(6, 35) <= 0; cloud_xl(6, 36) <= 0; cloud_xl(6, 37) <= 0; cloud_xl(6, 38) <= 0; cloud_xl(6, 39) <= 0; cloud_xl(6, 40) <= 0; cloud_xl(6, 41) <= 0; cloud_xl(6, 42) <= 0; cloud_xl(6, 43) <= 0; cloud_xl(6, 44) <= 0; cloud_xl(6, 45) <= 0; cloud_xl(6, 46) <= 0; cloud_xl(6, 47) <= 0; cloud_xl(6, 48) <= 1; cloud_xl(6, 49) <= 1; cloud_xl(6, 50) <= 1; cloud_xl(6, 51) <= 1; cloud_xl(6, 52) <= 1; cloud_xl(6, 53) <= 1; cloud_xl(6, 54) <= 2; cloud_xl(6, 55) <= 2; cloud_xl(6, 56) <= 2; cloud_xl(6, 57) <= 2; cloud_xl(6, 58) <= 2; cloud_xl(6, 59) <= 2; cloud_xl(6, 60) <= 2; cloud_xl(6, 61) <= 2; cloud_xl(6, 62) <= 2; cloud_xl(6, 63) <= 2; cloud_xl(6, 64) <= 2; cloud_xl(6, 65) <= 2; cloud_xl(6, 66) <= 2; cloud_xl(6, 67) <= 2; cloud_xl(6, 68) <= 2; cloud_xl(6, 69) <= 2; cloud_xl(6, 70) <= 2; cloud_xl(6, 71) <= 2; cloud_xl(6, 72) <= 2; cloud_xl(6, 73) <= 2; cloud_xl(6, 74) <= 2; cloud_xl(6, 75) <= 2; cloud_xl(6, 76) <= 2; cloud_xl(6, 77) <= 2; 
cloud_xl(7, 0) <= 2; cloud_xl(7, 1) <= 2; cloud_xl(7, 2) <= 2; cloud_xl(7, 3) <= 2; cloud_xl(7, 4) <= 2; cloud_xl(7, 5) <= 2; cloud_xl(7, 6) <= 2; cloud_xl(7, 7) <= 2; cloud_xl(7, 8) <= 2; cloud_xl(7, 9) <= 2; cloud_xl(7, 10) <= 2; cloud_xl(7, 11) <= 2; cloud_xl(7, 12) <= 2; cloud_xl(7, 13) <= 2; cloud_xl(7, 14) <= 2; cloud_xl(7, 15) <= 2; cloud_xl(7, 16) <= 2; cloud_xl(7, 17) <= 2; cloud_xl(7, 18) <= 2; cloud_xl(7, 19) <= 2; cloud_xl(7, 20) <= 2; cloud_xl(7, 21) <= 2; cloud_xl(7, 22) <= 2; cloud_xl(7, 23) <= 2; cloud_xl(7, 24) <= 1; cloud_xl(7, 25) <= 1; cloud_xl(7, 26) <= 1; cloud_xl(7, 27) <= 1; cloud_xl(7, 28) <= 1; cloud_xl(7, 29) <= 1; cloud_xl(7, 30) <= 0; cloud_xl(7, 31) <= 0; cloud_xl(7, 32) <= 0; cloud_xl(7, 33) <= 0; cloud_xl(7, 34) <= 0; cloud_xl(7, 35) <= 0; cloud_xl(7, 36) <= 0; cloud_xl(7, 37) <= 0; cloud_xl(7, 38) <= 0; cloud_xl(7, 39) <= 0; cloud_xl(7, 40) <= 0; cloud_xl(7, 41) <= 0; cloud_xl(7, 42) <= 0; cloud_xl(7, 43) <= 0; cloud_xl(7, 44) <= 0; cloud_xl(7, 45) <= 0; cloud_xl(7, 46) <= 0; cloud_xl(7, 47) <= 0; cloud_xl(7, 48) <= 1; cloud_xl(7, 49) <= 1; cloud_xl(7, 50) <= 1; cloud_xl(7, 51) <= 1; cloud_xl(7, 52) <= 1; cloud_xl(7, 53) <= 1; cloud_xl(7, 54) <= 2; cloud_xl(7, 55) <= 2; cloud_xl(7, 56) <= 2; cloud_xl(7, 57) <= 2; cloud_xl(7, 58) <= 2; cloud_xl(7, 59) <= 2; cloud_xl(7, 60) <= 2; cloud_xl(7, 61) <= 2; cloud_xl(7, 62) <= 2; cloud_xl(7, 63) <= 2; cloud_xl(7, 64) <= 2; cloud_xl(7, 65) <= 2; cloud_xl(7, 66) <= 2; cloud_xl(7, 67) <= 2; cloud_xl(7, 68) <= 2; cloud_xl(7, 69) <= 2; cloud_xl(7, 70) <= 2; cloud_xl(7, 71) <= 2; cloud_xl(7, 72) <= 2; cloud_xl(7, 73) <= 2; cloud_xl(7, 74) <= 2; cloud_xl(7, 75) <= 2; cloud_xl(7, 76) <= 2; cloud_xl(7, 77) <= 2; 
cloud_xl(8, 0) <= 2; cloud_xl(8, 1) <= 2; cloud_xl(8, 2) <= 2; cloud_xl(8, 3) <= 2; cloud_xl(8, 4) <= 2; cloud_xl(8, 5) <= 2; cloud_xl(8, 6) <= 2; cloud_xl(8, 7) <= 2; cloud_xl(8, 8) <= 2; cloud_xl(8, 9) <= 2; cloud_xl(8, 10) <= 2; cloud_xl(8, 11) <= 2; cloud_xl(8, 12) <= 2; cloud_xl(8, 13) <= 2; cloud_xl(8, 14) <= 2; cloud_xl(8, 15) <= 2; cloud_xl(8, 16) <= 2; cloud_xl(8, 17) <= 2; cloud_xl(8, 18) <= 2; cloud_xl(8, 19) <= 2; cloud_xl(8, 20) <= 2; cloud_xl(8, 21) <= 2; cloud_xl(8, 22) <= 2; cloud_xl(8, 23) <= 2; cloud_xl(8, 24) <= 1; cloud_xl(8, 25) <= 1; cloud_xl(8, 26) <= 1; cloud_xl(8, 27) <= 1; cloud_xl(8, 28) <= 1; cloud_xl(8, 29) <= 1; cloud_xl(8, 30) <= 0; cloud_xl(8, 31) <= 0; cloud_xl(8, 32) <= 0; cloud_xl(8, 33) <= 0; cloud_xl(8, 34) <= 0; cloud_xl(8, 35) <= 0; cloud_xl(8, 36) <= 0; cloud_xl(8, 37) <= 0; cloud_xl(8, 38) <= 0; cloud_xl(8, 39) <= 0; cloud_xl(8, 40) <= 0; cloud_xl(8, 41) <= 0; cloud_xl(8, 42) <= 0; cloud_xl(8, 43) <= 0; cloud_xl(8, 44) <= 0; cloud_xl(8, 45) <= 0; cloud_xl(8, 46) <= 0; cloud_xl(8, 47) <= 0; cloud_xl(8, 48) <= 1; cloud_xl(8, 49) <= 1; cloud_xl(8, 50) <= 1; cloud_xl(8, 51) <= 1; cloud_xl(8, 52) <= 1; cloud_xl(8, 53) <= 1; cloud_xl(8, 54) <= 2; cloud_xl(8, 55) <= 2; cloud_xl(8, 56) <= 2; cloud_xl(8, 57) <= 2; cloud_xl(8, 58) <= 2; cloud_xl(8, 59) <= 2; cloud_xl(8, 60) <= 2; cloud_xl(8, 61) <= 2; cloud_xl(8, 62) <= 2; cloud_xl(8, 63) <= 2; cloud_xl(8, 64) <= 2; cloud_xl(8, 65) <= 2; cloud_xl(8, 66) <= 2; cloud_xl(8, 67) <= 2; cloud_xl(8, 68) <= 2; cloud_xl(8, 69) <= 2; cloud_xl(8, 70) <= 2; cloud_xl(8, 71) <= 2; cloud_xl(8, 72) <= 2; cloud_xl(8, 73) <= 2; cloud_xl(8, 74) <= 2; cloud_xl(8, 75) <= 2; cloud_xl(8, 76) <= 2; cloud_xl(8, 77) <= 2; 
cloud_xl(9, 0) <= 2; cloud_xl(9, 1) <= 2; cloud_xl(9, 2) <= 2; cloud_xl(9, 3) <= 2; cloud_xl(9, 4) <= 2; cloud_xl(9, 5) <= 2; cloud_xl(9, 6) <= 2; cloud_xl(9, 7) <= 2; cloud_xl(9, 8) <= 2; cloud_xl(9, 9) <= 2; cloud_xl(9, 10) <= 2; cloud_xl(9, 11) <= 2; cloud_xl(9, 12) <= 2; cloud_xl(9, 13) <= 2; cloud_xl(9, 14) <= 2; cloud_xl(9, 15) <= 2; cloud_xl(9, 16) <= 2; cloud_xl(9, 17) <= 2; cloud_xl(9, 18) <= 2; cloud_xl(9, 19) <= 2; cloud_xl(9, 20) <= 2; cloud_xl(9, 21) <= 2; cloud_xl(9, 22) <= 2; cloud_xl(9, 23) <= 2; cloud_xl(9, 24) <= 1; cloud_xl(9, 25) <= 1; cloud_xl(9, 26) <= 1; cloud_xl(9, 27) <= 1; cloud_xl(9, 28) <= 1; cloud_xl(9, 29) <= 1; cloud_xl(9, 30) <= 0; cloud_xl(9, 31) <= 0; cloud_xl(9, 32) <= 0; cloud_xl(9, 33) <= 0; cloud_xl(9, 34) <= 0; cloud_xl(9, 35) <= 0; cloud_xl(9, 36) <= 0; cloud_xl(9, 37) <= 0; cloud_xl(9, 38) <= 0; cloud_xl(9, 39) <= 0; cloud_xl(9, 40) <= 0; cloud_xl(9, 41) <= 0; cloud_xl(9, 42) <= 0; cloud_xl(9, 43) <= 0; cloud_xl(9, 44) <= 0; cloud_xl(9, 45) <= 0; cloud_xl(9, 46) <= 0; cloud_xl(9, 47) <= 0; cloud_xl(9, 48) <= 1; cloud_xl(9, 49) <= 1; cloud_xl(9, 50) <= 1; cloud_xl(9, 51) <= 1; cloud_xl(9, 52) <= 1; cloud_xl(9, 53) <= 1; cloud_xl(9, 54) <= 2; cloud_xl(9, 55) <= 2; cloud_xl(9, 56) <= 2; cloud_xl(9, 57) <= 2; cloud_xl(9, 58) <= 2; cloud_xl(9, 59) <= 2; cloud_xl(9, 60) <= 2; cloud_xl(9, 61) <= 2; cloud_xl(9, 62) <= 2; cloud_xl(9, 63) <= 2; cloud_xl(9, 64) <= 2; cloud_xl(9, 65) <= 2; cloud_xl(9, 66) <= 2; cloud_xl(9, 67) <= 2; cloud_xl(9, 68) <= 2; cloud_xl(9, 69) <= 2; cloud_xl(9, 70) <= 2; cloud_xl(9, 71) <= 2; cloud_xl(9, 72) <= 2; cloud_xl(9, 73) <= 2; cloud_xl(9, 74) <= 2; cloud_xl(9, 75) <= 2; cloud_xl(9, 76) <= 2; cloud_xl(9, 77) <= 2; 
cloud_xl(10, 0) <= 2; cloud_xl(10, 1) <= 2; cloud_xl(10, 2) <= 2; cloud_xl(10, 3) <= 2; cloud_xl(10, 4) <= 2; cloud_xl(10, 5) <= 2; cloud_xl(10, 6) <= 2; cloud_xl(10, 7) <= 2; cloud_xl(10, 8) <= 2; cloud_xl(10, 9) <= 2; cloud_xl(10, 10) <= 2; cloud_xl(10, 11) <= 2; cloud_xl(10, 12) <= 2; cloud_xl(10, 13) <= 2; cloud_xl(10, 14) <= 2; cloud_xl(10, 15) <= 2; cloud_xl(10, 16) <= 2; cloud_xl(10, 17) <= 2; cloud_xl(10, 18) <= 2; cloud_xl(10, 19) <= 2; cloud_xl(10, 20) <= 2; cloud_xl(10, 21) <= 2; cloud_xl(10, 22) <= 2; cloud_xl(10, 23) <= 2; cloud_xl(10, 24) <= 1; cloud_xl(10, 25) <= 1; cloud_xl(10, 26) <= 1; cloud_xl(10, 27) <= 1; cloud_xl(10, 28) <= 1; cloud_xl(10, 29) <= 1; cloud_xl(10, 30) <= 0; cloud_xl(10, 31) <= 0; cloud_xl(10, 32) <= 0; cloud_xl(10, 33) <= 0; cloud_xl(10, 34) <= 0; cloud_xl(10, 35) <= 0; cloud_xl(10, 36) <= 0; cloud_xl(10, 37) <= 0; cloud_xl(10, 38) <= 0; cloud_xl(10, 39) <= 0; cloud_xl(10, 40) <= 0; cloud_xl(10, 41) <= 0; cloud_xl(10, 42) <= 0; cloud_xl(10, 43) <= 0; cloud_xl(10, 44) <= 0; cloud_xl(10, 45) <= 0; cloud_xl(10, 46) <= 0; cloud_xl(10, 47) <= 0; cloud_xl(10, 48) <= 1; cloud_xl(10, 49) <= 1; cloud_xl(10, 50) <= 1; cloud_xl(10, 51) <= 1; cloud_xl(10, 52) <= 1; cloud_xl(10, 53) <= 1; cloud_xl(10, 54) <= 2; cloud_xl(10, 55) <= 2; cloud_xl(10, 56) <= 2; cloud_xl(10, 57) <= 2; cloud_xl(10, 58) <= 2; cloud_xl(10, 59) <= 2; cloud_xl(10, 60) <= 2; cloud_xl(10, 61) <= 2; cloud_xl(10, 62) <= 2; cloud_xl(10, 63) <= 2; cloud_xl(10, 64) <= 2; cloud_xl(10, 65) <= 2; cloud_xl(10, 66) <= 2; cloud_xl(10, 67) <= 2; cloud_xl(10, 68) <= 2; cloud_xl(10, 69) <= 2; cloud_xl(10, 70) <= 2; cloud_xl(10, 71) <= 2; cloud_xl(10, 72) <= 2; cloud_xl(10, 73) <= 2; cloud_xl(10, 74) <= 2; cloud_xl(10, 75) <= 2; cloud_xl(10, 76) <= 2; cloud_xl(10, 77) <= 2; 
cloud_xl(11, 0) <= 2; cloud_xl(11, 1) <= 2; cloud_xl(11, 2) <= 2; cloud_xl(11, 3) <= 2; cloud_xl(11, 4) <= 2; cloud_xl(11, 5) <= 2; cloud_xl(11, 6) <= 2; cloud_xl(11, 7) <= 2; cloud_xl(11, 8) <= 2; cloud_xl(11, 9) <= 2; cloud_xl(11, 10) <= 2; cloud_xl(11, 11) <= 2; cloud_xl(11, 12) <= 2; cloud_xl(11, 13) <= 2; cloud_xl(11, 14) <= 2; cloud_xl(11, 15) <= 2; cloud_xl(11, 16) <= 2; cloud_xl(11, 17) <= 2; cloud_xl(11, 18) <= 2; cloud_xl(11, 19) <= 2; cloud_xl(11, 20) <= 2; cloud_xl(11, 21) <= 2; cloud_xl(11, 22) <= 2; cloud_xl(11, 23) <= 2; cloud_xl(11, 24) <= 1; cloud_xl(11, 25) <= 1; cloud_xl(11, 26) <= 1; cloud_xl(11, 27) <= 1; cloud_xl(11, 28) <= 1; cloud_xl(11, 29) <= 1; cloud_xl(11, 30) <= 0; cloud_xl(11, 31) <= 0; cloud_xl(11, 32) <= 0; cloud_xl(11, 33) <= 0; cloud_xl(11, 34) <= 0; cloud_xl(11, 35) <= 0; cloud_xl(11, 36) <= 0; cloud_xl(11, 37) <= 0; cloud_xl(11, 38) <= 0; cloud_xl(11, 39) <= 0; cloud_xl(11, 40) <= 0; cloud_xl(11, 41) <= 0; cloud_xl(11, 42) <= 0; cloud_xl(11, 43) <= 0; cloud_xl(11, 44) <= 0; cloud_xl(11, 45) <= 0; cloud_xl(11, 46) <= 0; cloud_xl(11, 47) <= 0; cloud_xl(11, 48) <= 1; cloud_xl(11, 49) <= 1; cloud_xl(11, 50) <= 1; cloud_xl(11, 51) <= 1; cloud_xl(11, 52) <= 1; cloud_xl(11, 53) <= 1; cloud_xl(11, 54) <= 2; cloud_xl(11, 55) <= 2; cloud_xl(11, 56) <= 2; cloud_xl(11, 57) <= 2; cloud_xl(11, 58) <= 2; cloud_xl(11, 59) <= 2; cloud_xl(11, 60) <= 2; cloud_xl(11, 61) <= 2; cloud_xl(11, 62) <= 2; cloud_xl(11, 63) <= 2; cloud_xl(11, 64) <= 2; cloud_xl(11, 65) <= 2; cloud_xl(11, 66) <= 2; cloud_xl(11, 67) <= 2; cloud_xl(11, 68) <= 2; cloud_xl(11, 69) <= 2; cloud_xl(11, 70) <= 2; cloud_xl(11, 71) <= 2; cloud_xl(11, 72) <= 2; cloud_xl(11, 73) <= 2; cloud_xl(11, 74) <= 2; cloud_xl(11, 75) <= 2; cloud_xl(11, 76) <= 2; cloud_xl(11, 77) <= 2; 
cloud_xl(12, 0) <= 2; cloud_xl(12, 1) <= 2; cloud_xl(12, 2) <= 2; cloud_xl(12, 3) <= 2; cloud_xl(12, 4) <= 2; cloud_xl(12, 5) <= 2; cloud_xl(12, 6) <= 2; cloud_xl(12, 7) <= 2; cloud_xl(12, 8) <= 2; cloud_xl(12, 9) <= 2; cloud_xl(12, 10) <= 2; cloud_xl(12, 11) <= 2; cloud_xl(12, 12) <= 1; cloud_xl(12, 13) <= 1; cloud_xl(12, 14) <= 1; cloud_xl(12, 15) <= 1; cloud_xl(12, 16) <= 1; cloud_xl(12, 17) <= 1; cloud_xl(12, 18) <= 1; cloud_xl(12, 19) <= 1; cloud_xl(12, 20) <= 1; cloud_xl(12, 21) <= 1; cloud_xl(12, 22) <= 1; cloud_xl(12, 23) <= 1; cloud_xl(12, 24) <= 0; cloud_xl(12, 25) <= 0; cloud_xl(12, 26) <= 0; cloud_xl(12, 27) <= 0; cloud_xl(12, 28) <= 0; cloud_xl(12, 29) <= 0; cloud_xl(12, 30) <= 0; cloud_xl(12, 31) <= 0; cloud_xl(12, 32) <= 0; cloud_xl(12, 33) <= 0; cloud_xl(12, 34) <= 0; cloud_xl(12, 35) <= 0; cloud_xl(12, 36) <= 0; cloud_xl(12, 37) <= 0; cloud_xl(12, 38) <= 0; cloud_xl(12, 39) <= 0; cloud_xl(12, 40) <= 0; cloud_xl(12, 41) <= 0; cloud_xl(12, 42) <= 0; cloud_xl(12, 43) <= 0; cloud_xl(12, 44) <= 0; cloud_xl(12, 45) <= 0; cloud_xl(12, 46) <= 0; cloud_xl(12, 47) <= 0; cloud_xl(12, 48) <= 0; cloud_xl(12, 49) <= 0; cloud_xl(12, 50) <= 0; cloud_xl(12, 51) <= 0; cloud_xl(12, 52) <= 0; cloud_xl(12, 53) <= 0; cloud_xl(12, 54) <= 1; cloud_xl(12, 55) <= 1; cloud_xl(12, 56) <= 1; cloud_xl(12, 57) <= 1; cloud_xl(12, 58) <= 1; cloud_xl(12, 59) <= 1; cloud_xl(12, 60) <= 2; cloud_xl(12, 61) <= 2; cloud_xl(12, 62) <= 2; cloud_xl(12, 63) <= 2; cloud_xl(12, 64) <= 2; cloud_xl(12, 65) <= 2; cloud_xl(12, 66) <= 2; cloud_xl(12, 67) <= 2; cloud_xl(12, 68) <= 2; cloud_xl(12, 69) <= 2; cloud_xl(12, 70) <= 2; cloud_xl(12, 71) <= 2; cloud_xl(12, 72) <= 2; cloud_xl(12, 73) <= 2; cloud_xl(12, 74) <= 2; cloud_xl(12, 75) <= 2; cloud_xl(12, 76) <= 2; cloud_xl(12, 77) <= 2; 
cloud_xl(13, 0) <= 2; cloud_xl(13, 1) <= 2; cloud_xl(13, 2) <= 2; cloud_xl(13, 3) <= 2; cloud_xl(13, 4) <= 2; cloud_xl(13, 5) <= 2; cloud_xl(13, 6) <= 2; cloud_xl(13, 7) <= 2; cloud_xl(13, 8) <= 2; cloud_xl(13, 9) <= 2; cloud_xl(13, 10) <= 2; cloud_xl(13, 11) <= 2; cloud_xl(13, 12) <= 1; cloud_xl(13, 13) <= 1; cloud_xl(13, 14) <= 1; cloud_xl(13, 15) <= 1; cloud_xl(13, 16) <= 1; cloud_xl(13, 17) <= 1; cloud_xl(13, 18) <= 1; cloud_xl(13, 19) <= 1; cloud_xl(13, 20) <= 1; cloud_xl(13, 21) <= 1; cloud_xl(13, 22) <= 1; cloud_xl(13, 23) <= 1; cloud_xl(13, 24) <= 0; cloud_xl(13, 25) <= 0; cloud_xl(13, 26) <= 0; cloud_xl(13, 27) <= 0; cloud_xl(13, 28) <= 0; cloud_xl(13, 29) <= 0; cloud_xl(13, 30) <= 0; cloud_xl(13, 31) <= 0; cloud_xl(13, 32) <= 0; cloud_xl(13, 33) <= 0; cloud_xl(13, 34) <= 0; cloud_xl(13, 35) <= 0; cloud_xl(13, 36) <= 0; cloud_xl(13, 37) <= 0; cloud_xl(13, 38) <= 0; cloud_xl(13, 39) <= 0; cloud_xl(13, 40) <= 0; cloud_xl(13, 41) <= 0; cloud_xl(13, 42) <= 0; cloud_xl(13, 43) <= 0; cloud_xl(13, 44) <= 0; cloud_xl(13, 45) <= 0; cloud_xl(13, 46) <= 0; cloud_xl(13, 47) <= 0; cloud_xl(13, 48) <= 0; cloud_xl(13, 49) <= 0; cloud_xl(13, 50) <= 0; cloud_xl(13, 51) <= 0; cloud_xl(13, 52) <= 0; cloud_xl(13, 53) <= 0; cloud_xl(13, 54) <= 1; cloud_xl(13, 55) <= 1; cloud_xl(13, 56) <= 1; cloud_xl(13, 57) <= 1; cloud_xl(13, 58) <= 1; cloud_xl(13, 59) <= 1; cloud_xl(13, 60) <= 2; cloud_xl(13, 61) <= 2; cloud_xl(13, 62) <= 2; cloud_xl(13, 63) <= 2; cloud_xl(13, 64) <= 2; cloud_xl(13, 65) <= 2; cloud_xl(13, 66) <= 2; cloud_xl(13, 67) <= 2; cloud_xl(13, 68) <= 2; cloud_xl(13, 69) <= 2; cloud_xl(13, 70) <= 2; cloud_xl(13, 71) <= 2; cloud_xl(13, 72) <= 2; cloud_xl(13, 73) <= 2; cloud_xl(13, 74) <= 2; cloud_xl(13, 75) <= 2; cloud_xl(13, 76) <= 2; cloud_xl(13, 77) <= 2; 
cloud_xl(14, 0) <= 2; cloud_xl(14, 1) <= 2; cloud_xl(14, 2) <= 2; cloud_xl(14, 3) <= 2; cloud_xl(14, 4) <= 2; cloud_xl(14, 5) <= 2; cloud_xl(14, 6) <= 2; cloud_xl(14, 7) <= 2; cloud_xl(14, 8) <= 2; cloud_xl(14, 9) <= 2; cloud_xl(14, 10) <= 2; cloud_xl(14, 11) <= 2; cloud_xl(14, 12) <= 1; cloud_xl(14, 13) <= 1; cloud_xl(14, 14) <= 1; cloud_xl(14, 15) <= 1; cloud_xl(14, 16) <= 1; cloud_xl(14, 17) <= 1; cloud_xl(14, 18) <= 1; cloud_xl(14, 19) <= 1; cloud_xl(14, 20) <= 1; cloud_xl(14, 21) <= 1; cloud_xl(14, 22) <= 1; cloud_xl(14, 23) <= 1; cloud_xl(14, 24) <= 0; cloud_xl(14, 25) <= 0; cloud_xl(14, 26) <= 0; cloud_xl(14, 27) <= 0; cloud_xl(14, 28) <= 0; cloud_xl(14, 29) <= 0; cloud_xl(14, 30) <= 0; cloud_xl(14, 31) <= 0; cloud_xl(14, 32) <= 0; cloud_xl(14, 33) <= 0; cloud_xl(14, 34) <= 0; cloud_xl(14, 35) <= 0; cloud_xl(14, 36) <= 0; cloud_xl(14, 37) <= 0; cloud_xl(14, 38) <= 0; cloud_xl(14, 39) <= 0; cloud_xl(14, 40) <= 0; cloud_xl(14, 41) <= 0; cloud_xl(14, 42) <= 0; cloud_xl(14, 43) <= 0; cloud_xl(14, 44) <= 0; cloud_xl(14, 45) <= 0; cloud_xl(14, 46) <= 0; cloud_xl(14, 47) <= 0; cloud_xl(14, 48) <= 0; cloud_xl(14, 49) <= 0; cloud_xl(14, 50) <= 0; cloud_xl(14, 51) <= 0; cloud_xl(14, 52) <= 0; cloud_xl(14, 53) <= 0; cloud_xl(14, 54) <= 1; cloud_xl(14, 55) <= 1; cloud_xl(14, 56) <= 1; cloud_xl(14, 57) <= 1; cloud_xl(14, 58) <= 1; cloud_xl(14, 59) <= 1; cloud_xl(14, 60) <= 2; cloud_xl(14, 61) <= 2; cloud_xl(14, 62) <= 2; cloud_xl(14, 63) <= 2; cloud_xl(14, 64) <= 2; cloud_xl(14, 65) <= 2; cloud_xl(14, 66) <= 2; cloud_xl(14, 67) <= 2; cloud_xl(14, 68) <= 2; cloud_xl(14, 69) <= 2; cloud_xl(14, 70) <= 2; cloud_xl(14, 71) <= 2; cloud_xl(14, 72) <= 2; cloud_xl(14, 73) <= 2; cloud_xl(14, 74) <= 2; cloud_xl(14, 75) <= 2; cloud_xl(14, 76) <= 2; cloud_xl(14, 77) <= 2; 
cloud_xl(15, 0) <= 2; cloud_xl(15, 1) <= 2; cloud_xl(15, 2) <= 2; cloud_xl(15, 3) <= 2; cloud_xl(15, 4) <= 2; cloud_xl(15, 5) <= 2; cloud_xl(15, 6) <= 2; cloud_xl(15, 7) <= 2; cloud_xl(15, 8) <= 2; cloud_xl(15, 9) <= 2; cloud_xl(15, 10) <= 2; cloud_xl(15, 11) <= 2; cloud_xl(15, 12) <= 1; cloud_xl(15, 13) <= 1; cloud_xl(15, 14) <= 1; cloud_xl(15, 15) <= 1; cloud_xl(15, 16) <= 1; cloud_xl(15, 17) <= 1; cloud_xl(15, 18) <= 1; cloud_xl(15, 19) <= 1; cloud_xl(15, 20) <= 1; cloud_xl(15, 21) <= 1; cloud_xl(15, 22) <= 1; cloud_xl(15, 23) <= 1; cloud_xl(15, 24) <= 0; cloud_xl(15, 25) <= 0; cloud_xl(15, 26) <= 0; cloud_xl(15, 27) <= 0; cloud_xl(15, 28) <= 0; cloud_xl(15, 29) <= 0; cloud_xl(15, 30) <= 0; cloud_xl(15, 31) <= 0; cloud_xl(15, 32) <= 0; cloud_xl(15, 33) <= 0; cloud_xl(15, 34) <= 0; cloud_xl(15, 35) <= 0; cloud_xl(15, 36) <= 0; cloud_xl(15, 37) <= 0; cloud_xl(15, 38) <= 0; cloud_xl(15, 39) <= 0; cloud_xl(15, 40) <= 0; cloud_xl(15, 41) <= 0; cloud_xl(15, 42) <= 0; cloud_xl(15, 43) <= 0; cloud_xl(15, 44) <= 0; cloud_xl(15, 45) <= 0; cloud_xl(15, 46) <= 0; cloud_xl(15, 47) <= 0; cloud_xl(15, 48) <= 0; cloud_xl(15, 49) <= 0; cloud_xl(15, 50) <= 0; cloud_xl(15, 51) <= 0; cloud_xl(15, 52) <= 0; cloud_xl(15, 53) <= 0; cloud_xl(15, 54) <= 1; cloud_xl(15, 55) <= 1; cloud_xl(15, 56) <= 1; cloud_xl(15, 57) <= 1; cloud_xl(15, 58) <= 1; cloud_xl(15, 59) <= 1; cloud_xl(15, 60) <= 2; cloud_xl(15, 61) <= 2; cloud_xl(15, 62) <= 2; cloud_xl(15, 63) <= 2; cloud_xl(15, 64) <= 2; cloud_xl(15, 65) <= 2; cloud_xl(15, 66) <= 2; cloud_xl(15, 67) <= 2; cloud_xl(15, 68) <= 2; cloud_xl(15, 69) <= 2; cloud_xl(15, 70) <= 2; cloud_xl(15, 71) <= 2; cloud_xl(15, 72) <= 2; cloud_xl(15, 73) <= 2; cloud_xl(15, 74) <= 2; cloud_xl(15, 75) <= 2; cloud_xl(15, 76) <= 2; cloud_xl(15, 77) <= 2; 
cloud_xl(16, 0) <= 2; cloud_xl(16, 1) <= 2; cloud_xl(16, 2) <= 2; cloud_xl(16, 3) <= 2; cloud_xl(16, 4) <= 2; cloud_xl(16, 5) <= 2; cloud_xl(16, 6) <= 2; cloud_xl(16, 7) <= 2; cloud_xl(16, 8) <= 2; cloud_xl(16, 9) <= 2; cloud_xl(16, 10) <= 2; cloud_xl(16, 11) <= 2; cloud_xl(16, 12) <= 1; cloud_xl(16, 13) <= 1; cloud_xl(16, 14) <= 1; cloud_xl(16, 15) <= 1; cloud_xl(16, 16) <= 1; cloud_xl(16, 17) <= 1; cloud_xl(16, 18) <= 1; cloud_xl(16, 19) <= 1; cloud_xl(16, 20) <= 1; cloud_xl(16, 21) <= 1; cloud_xl(16, 22) <= 1; cloud_xl(16, 23) <= 1; cloud_xl(16, 24) <= 0; cloud_xl(16, 25) <= 0; cloud_xl(16, 26) <= 0; cloud_xl(16, 27) <= 0; cloud_xl(16, 28) <= 0; cloud_xl(16, 29) <= 0; cloud_xl(16, 30) <= 0; cloud_xl(16, 31) <= 0; cloud_xl(16, 32) <= 0; cloud_xl(16, 33) <= 0; cloud_xl(16, 34) <= 0; cloud_xl(16, 35) <= 0; cloud_xl(16, 36) <= 0; cloud_xl(16, 37) <= 0; cloud_xl(16, 38) <= 0; cloud_xl(16, 39) <= 0; cloud_xl(16, 40) <= 0; cloud_xl(16, 41) <= 0; cloud_xl(16, 42) <= 0; cloud_xl(16, 43) <= 0; cloud_xl(16, 44) <= 0; cloud_xl(16, 45) <= 0; cloud_xl(16, 46) <= 0; cloud_xl(16, 47) <= 0; cloud_xl(16, 48) <= 0; cloud_xl(16, 49) <= 0; cloud_xl(16, 50) <= 0; cloud_xl(16, 51) <= 0; cloud_xl(16, 52) <= 0; cloud_xl(16, 53) <= 0; cloud_xl(16, 54) <= 1; cloud_xl(16, 55) <= 1; cloud_xl(16, 56) <= 1; cloud_xl(16, 57) <= 1; cloud_xl(16, 58) <= 1; cloud_xl(16, 59) <= 1; cloud_xl(16, 60) <= 2; cloud_xl(16, 61) <= 2; cloud_xl(16, 62) <= 2; cloud_xl(16, 63) <= 2; cloud_xl(16, 64) <= 2; cloud_xl(16, 65) <= 2; cloud_xl(16, 66) <= 2; cloud_xl(16, 67) <= 2; cloud_xl(16, 68) <= 2; cloud_xl(16, 69) <= 2; cloud_xl(16, 70) <= 2; cloud_xl(16, 71) <= 2; cloud_xl(16, 72) <= 2; cloud_xl(16, 73) <= 2; cloud_xl(16, 74) <= 2; cloud_xl(16, 75) <= 2; cloud_xl(16, 76) <= 2; cloud_xl(16, 77) <= 2; 
cloud_xl(17, 0) <= 2; cloud_xl(17, 1) <= 2; cloud_xl(17, 2) <= 2; cloud_xl(17, 3) <= 2; cloud_xl(17, 4) <= 2; cloud_xl(17, 5) <= 2; cloud_xl(17, 6) <= 2; cloud_xl(17, 7) <= 2; cloud_xl(17, 8) <= 2; cloud_xl(17, 9) <= 2; cloud_xl(17, 10) <= 2; cloud_xl(17, 11) <= 2; cloud_xl(17, 12) <= 1; cloud_xl(17, 13) <= 1; cloud_xl(17, 14) <= 1; cloud_xl(17, 15) <= 1; cloud_xl(17, 16) <= 1; cloud_xl(17, 17) <= 1; cloud_xl(17, 18) <= 1; cloud_xl(17, 19) <= 1; cloud_xl(17, 20) <= 1; cloud_xl(17, 21) <= 1; cloud_xl(17, 22) <= 1; cloud_xl(17, 23) <= 1; cloud_xl(17, 24) <= 0; cloud_xl(17, 25) <= 0; cloud_xl(17, 26) <= 0; cloud_xl(17, 27) <= 0; cloud_xl(17, 28) <= 0; cloud_xl(17, 29) <= 0; cloud_xl(17, 30) <= 0; cloud_xl(17, 31) <= 0; cloud_xl(17, 32) <= 0; cloud_xl(17, 33) <= 0; cloud_xl(17, 34) <= 0; cloud_xl(17, 35) <= 0; cloud_xl(17, 36) <= 0; cloud_xl(17, 37) <= 0; cloud_xl(17, 38) <= 0; cloud_xl(17, 39) <= 0; cloud_xl(17, 40) <= 0; cloud_xl(17, 41) <= 0; cloud_xl(17, 42) <= 0; cloud_xl(17, 43) <= 0; cloud_xl(17, 44) <= 0; cloud_xl(17, 45) <= 0; cloud_xl(17, 46) <= 0; cloud_xl(17, 47) <= 0; cloud_xl(17, 48) <= 0; cloud_xl(17, 49) <= 0; cloud_xl(17, 50) <= 0; cloud_xl(17, 51) <= 0; cloud_xl(17, 52) <= 0; cloud_xl(17, 53) <= 0; cloud_xl(17, 54) <= 1; cloud_xl(17, 55) <= 1; cloud_xl(17, 56) <= 1; cloud_xl(17, 57) <= 1; cloud_xl(17, 58) <= 1; cloud_xl(17, 59) <= 1; cloud_xl(17, 60) <= 2; cloud_xl(17, 61) <= 2; cloud_xl(17, 62) <= 2; cloud_xl(17, 63) <= 2; cloud_xl(17, 64) <= 2; cloud_xl(17, 65) <= 2; cloud_xl(17, 66) <= 2; cloud_xl(17, 67) <= 2; cloud_xl(17, 68) <= 2; cloud_xl(17, 69) <= 2; cloud_xl(17, 70) <= 2; cloud_xl(17, 71) <= 2; cloud_xl(17, 72) <= 2; cloud_xl(17, 73) <= 2; cloud_xl(17, 74) <= 2; cloud_xl(17, 75) <= 2; cloud_xl(17, 76) <= 2; cloud_xl(17, 77) <= 2; 
cloud_xl(18, 0) <= 2; cloud_xl(18, 1) <= 2; cloud_xl(18, 2) <= 2; cloud_xl(18, 3) <= 2; cloud_xl(18, 4) <= 2; cloud_xl(18, 5) <= 2; cloud_xl(18, 6) <= 1; cloud_xl(18, 7) <= 1; cloud_xl(18, 8) <= 1; cloud_xl(18, 9) <= 1; cloud_xl(18, 10) <= 1; cloud_xl(18, 11) <= 1; cloud_xl(18, 12) <= 0; cloud_xl(18, 13) <= 0; cloud_xl(18, 14) <= 0; cloud_xl(18, 15) <= 0; cloud_xl(18, 16) <= 0; cloud_xl(18, 17) <= 0; cloud_xl(18, 18) <= 0; cloud_xl(18, 19) <= 0; cloud_xl(18, 20) <= 0; cloud_xl(18, 21) <= 0; cloud_xl(18, 22) <= 0; cloud_xl(18, 23) <= 0; cloud_xl(18, 24) <= 0; cloud_xl(18, 25) <= 0; cloud_xl(18, 26) <= 0; cloud_xl(18, 27) <= 0; cloud_xl(18, 28) <= 0; cloud_xl(18, 29) <= 0; cloud_xl(18, 30) <= 0; cloud_xl(18, 31) <= 0; cloud_xl(18, 32) <= 0; cloud_xl(18, 33) <= 0; cloud_xl(18, 34) <= 0; cloud_xl(18, 35) <= 0; cloud_xl(18, 36) <= 0; cloud_xl(18, 37) <= 0; cloud_xl(18, 38) <= 0; cloud_xl(18, 39) <= 0; cloud_xl(18, 40) <= 0; cloud_xl(18, 41) <= 0; cloud_xl(18, 42) <= 0; cloud_xl(18, 43) <= 0; cloud_xl(18, 44) <= 0; cloud_xl(18, 45) <= 0; cloud_xl(18, 46) <= 0; cloud_xl(18, 47) <= 0; cloud_xl(18, 48) <= 0; cloud_xl(18, 49) <= 0; cloud_xl(18, 50) <= 0; cloud_xl(18, 51) <= 0; cloud_xl(18, 52) <= 0; cloud_xl(18, 53) <= 0; cloud_xl(18, 54) <= 0; cloud_xl(18, 55) <= 0; cloud_xl(18, 56) <= 0; cloud_xl(18, 57) <= 0; cloud_xl(18, 58) <= 0; cloud_xl(18, 59) <= 0; cloud_xl(18, 60) <= 1; cloud_xl(18, 61) <= 1; cloud_xl(18, 62) <= 1; cloud_xl(18, 63) <= 1; cloud_xl(18, 64) <= 1; cloud_xl(18, 65) <= 1; cloud_xl(18, 66) <= 1; cloud_xl(18, 67) <= 1; cloud_xl(18, 68) <= 1; cloud_xl(18, 69) <= 1; cloud_xl(18, 70) <= 1; cloud_xl(18, 71) <= 1; cloud_xl(18, 72) <= 2; cloud_xl(18, 73) <= 2; cloud_xl(18, 74) <= 2; cloud_xl(18, 75) <= 2; cloud_xl(18, 76) <= 2; cloud_xl(18, 77) <= 2; 
cloud_xl(19, 0) <= 2; cloud_xl(19, 1) <= 2; cloud_xl(19, 2) <= 2; cloud_xl(19, 3) <= 2; cloud_xl(19, 4) <= 2; cloud_xl(19, 5) <= 2; cloud_xl(19, 6) <= 1; cloud_xl(19, 7) <= 1; cloud_xl(19, 8) <= 1; cloud_xl(19, 9) <= 1; cloud_xl(19, 10) <= 1; cloud_xl(19, 11) <= 1; cloud_xl(19, 12) <= 0; cloud_xl(19, 13) <= 0; cloud_xl(19, 14) <= 0; cloud_xl(19, 15) <= 0; cloud_xl(19, 16) <= 0; cloud_xl(19, 17) <= 0; cloud_xl(19, 18) <= 0; cloud_xl(19, 19) <= 0; cloud_xl(19, 20) <= 0; cloud_xl(19, 21) <= 0; cloud_xl(19, 22) <= 0; cloud_xl(19, 23) <= 0; cloud_xl(19, 24) <= 0; cloud_xl(19, 25) <= 0; cloud_xl(19, 26) <= 0; cloud_xl(19, 27) <= 0; cloud_xl(19, 28) <= 0; cloud_xl(19, 29) <= 0; cloud_xl(19, 30) <= 0; cloud_xl(19, 31) <= 0; cloud_xl(19, 32) <= 0; cloud_xl(19, 33) <= 0; cloud_xl(19, 34) <= 0; cloud_xl(19, 35) <= 0; cloud_xl(19, 36) <= 0; cloud_xl(19, 37) <= 0; cloud_xl(19, 38) <= 0; cloud_xl(19, 39) <= 0; cloud_xl(19, 40) <= 0; cloud_xl(19, 41) <= 0; cloud_xl(19, 42) <= 0; cloud_xl(19, 43) <= 0; cloud_xl(19, 44) <= 0; cloud_xl(19, 45) <= 0; cloud_xl(19, 46) <= 0; cloud_xl(19, 47) <= 0; cloud_xl(19, 48) <= 0; cloud_xl(19, 49) <= 0; cloud_xl(19, 50) <= 0; cloud_xl(19, 51) <= 0; cloud_xl(19, 52) <= 0; cloud_xl(19, 53) <= 0; cloud_xl(19, 54) <= 0; cloud_xl(19, 55) <= 0; cloud_xl(19, 56) <= 0; cloud_xl(19, 57) <= 0; cloud_xl(19, 58) <= 0; cloud_xl(19, 59) <= 0; cloud_xl(19, 60) <= 1; cloud_xl(19, 61) <= 1; cloud_xl(19, 62) <= 1; cloud_xl(19, 63) <= 1; cloud_xl(19, 64) <= 1; cloud_xl(19, 65) <= 1; cloud_xl(19, 66) <= 1; cloud_xl(19, 67) <= 1; cloud_xl(19, 68) <= 1; cloud_xl(19, 69) <= 1; cloud_xl(19, 70) <= 1; cloud_xl(19, 71) <= 1; cloud_xl(19, 72) <= 2; cloud_xl(19, 73) <= 2; cloud_xl(19, 74) <= 2; cloud_xl(19, 75) <= 2; cloud_xl(19, 76) <= 2; cloud_xl(19, 77) <= 2; 
cloud_xl(20, 0) <= 2; cloud_xl(20, 1) <= 2; cloud_xl(20, 2) <= 2; cloud_xl(20, 3) <= 2; cloud_xl(20, 4) <= 2; cloud_xl(20, 5) <= 2; cloud_xl(20, 6) <= 1; cloud_xl(20, 7) <= 1; cloud_xl(20, 8) <= 1; cloud_xl(20, 9) <= 1; cloud_xl(20, 10) <= 1; cloud_xl(20, 11) <= 1; cloud_xl(20, 12) <= 0; cloud_xl(20, 13) <= 0; cloud_xl(20, 14) <= 0; cloud_xl(20, 15) <= 0; cloud_xl(20, 16) <= 0; cloud_xl(20, 17) <= 0; cloud_xl(20, 18) <= 0; cloud_xl(20, 19) <= 0; cloud_xl(20, 20) <= 0; cloud_xl(20, 21) <= 0; cloud_xl(20, 22) <= 0; cloud_xl(20, 23) <= 0; cloud_xl(20, 24) <= 0; cloud_xl(20, 25) <= 0; cloud_xl(20, 26) <= 0; cloud_xl(20, 27) <= 0; cloud_xl(20, 28) <= 0; cloud_xl(20, 29) <= 0; cloud_xl(20, 30) <= 0; cloud_xl(20, 31) <= 0; cloud_xl(20, 32) <= 0; cloud_xl(20, 33) <= 0; cloud_xl(20, 34) <= 0; cloud_xl(20, 35) <= 0; cloud_xl(20, 36) <= 0; cloud_xl(20, 37) <= 0; cloud_xl(20, 38) <= 0; cloud_xl(20, 39) <= 0; cloud_xl(20, 40) <= 0; cloud_xl(20, 41) <= 0; cloud_xl(20, 42) <= 0; cloud_xl(20, 43) <= 0; cloud_xl(20, 44) <= 0; cloud_xl(20, 45) <= 0; cloud_xl(20, 46) <= 0; cloud_xl(20, 47) <= 0; cloud_xl(20, 48) <= 0; cloud_xl(20, 49) <= 0; cloud_xl(20, 50) <= 0; cloud_xl(20, 51) <= 0; cloud_xl(20, 52) <= 0; cloud_xl(20, 53) <= 0; cloud_xl(20, 54) <= 0; cloud_xl(20, 55) <= 0; cloud_xl(20, 56) <= 0; cloud_xl(20, 57) <= 0; cloud_xl(20, 58) <= 0; cloud_xl(20, 59) <= 0; cloud_xl(20, 60) <= 1; cloud_xl(20, 61) <= 1; cloud_xl(20, 62) <= 1; cloud_xl(20, 63) <= 1; cloud_xl(20, 64) <= 1; cloud_xl(20, 65) <= 1; cloud_xl(20, 66) <= 1; cloud_xl(20, 67) <= 1; cloud_xl(20, 68) <= 1; cloud_xl(20, 69) <= 1; cloud_xl(20, 70) <= 1; cloud_xl(20, 71) <= 1; cloud_xl(20, 72) <= 2; cloud_xl(20, 73) <= 2; cloud_xl(20, 74) <= 2; cloud_xl(20, 75) <= 2; cloud_xl(20, 76) <= 2; cloud_xl(20, 77) <= 2; 
cloud_xl(21, 0) <= 2; cloud_xl(21, 1) <= 2; cloud_xl(21, 2) <= 2; cloud_xl(21, 3) <= 2; cloud_xl(21, 4) <= 2; cloud_xl(21, 5) <= 2; cloud_xl(21, 6) <= 1; cloud_xl(21, 7) <= 1; cloud_xl(21, 8) <= 1; cloud_xl(21, 9) <= 1; cloud_xl(21, 10) <= 1; cloud_xl(21, 11) <= 1; cloud_xl(21, 12) <= 0; cloud_xl(21, 13) <= 0; cloud_xl(21, 14) <= 0; cloud_xl(21, 15) <= 0; cloud_xl(21, 16) <= 0; cloud_xl(21, 17) <= 0; cloud_xl(21, 18) <= 0; cloud_xl(21, 19) <= 0; cloud_xl(21, 20) <= 0; cloud_xl(21, 21) <= 0; cloud_xl(21, 22) <= 0; cloud_xl(21, 23) <= 0; cloud_xl(21, 24) <= 0; cloud_xl(21, 25) <= 0; cloud_xl(21, 26) <= 0; cloud_xl(21, 27) <= 0; cloud_xl(21, 28) <= 0; cloud_xl(21, 29) <= 0; cloud_xl(21, 30) <= 0; cloud_xl(21, 31) <= 0; cloud_xl(21, 32) <= 0; cloud_xl(21, 33) <= 0; cloud_xl(21, 34) <= 0; cloud_xl(21, 35) <= 0; cloud_xl(21, 36) <= 0; cloud_xl(21, 37) <= 0; cloud_xl(21, 38) <= 0; cloud_xl(21, 39) <= 0; cloud_xl(21, 40) <= 0; cloud_xl(21, 41) <= 0; cloud_xl(21, 42) <= 0; cloud_xl(21, 43) <= 0; cloud_xl(21, 44) <= 0; cloud_xl(21, 45) <= 0; cloud_xl(21, 46) <= 0; cloud_xl(21, 47) <= 0; cloud_xl(21, 48) <= 0; cloud_xl(21, 49) <= 0; cloud_xl(21, 50) <= 0; cloud_xl(21, 51) <= 0; cloud_xl(21, 52) <= 0; cloud_xl(21, 53) <= 0; cloud_xl(21, 54) <= 0; cloud_xl(21, 55) <= 0; cloud_xl(21, 56) <= 0; cloud_xl(21, 57) <= 0; cloud_xl(21, 58) <= 0; cloud_xl(21, 59) <= 0; cloud_xl(21, 60) <= 1; cloud_xl(21, 61) <= 1; cloud_xl(21, 62) <= 1; cloud_xl(21, 63) <= 1; cloud_xl(21, 64) <= 1; cloud_xl(21, 65) <= 1; cloud_xl(21, 66) <= 1; cloud_xl(21, 67) <= 1; cloud_xl(21, 68) <= 1; cloud_xl(21, 69) <= 1; cloud_xl(21, 70) <= 1; cloud_xl(21, 71) <= 1; cloud_xl(21, 72) <= 2; cloud_xl(21, 73) <= 2; cloud_xl(21, 74) <= 2; cloud_xl(21, 75) <= 2; cloud_xl(21, 76) <= 2; cloud_xl(21, 77) <= 2; 
cloud_xl(22, 0) <= 2; cloud_xl(22, 1) <= 2; cloud_xl(22, 2) <= 2; cloud_xl(22, 3) <= 2; cloud_xl(22, 4) <= 2; cloud_xl(22, 5) <= 2; cloud_xl(22, 6) <= 1; cloud_xl(22, 7) <= 1; cloud_xl(22, 8) <= 1; cloud_xl(22, 9) <= 1; cloud_xl(22, 10) <= 1; cloud_xl(22, 11) <= 1; cloud_xl(22, 12) <= 0; cloud_xl(22, 13) <= 0; cloud_xl(22, 14) <= 0; cloud_xl(22, 15) <= 0; cloud_xl(22, 16) <= 0; cloud_xl(22, 17) <= 0; cloud_xl(22, 18) <= 0; cloud_xl(22, 19) <= 0; cloud_xl(22, 20) <= 0; cloud_xl(22, 21) <= 0; cloud_xl(22, 22) <= 0; cloud_xl(22, 23) <= 0; cloud_xl(22, 24) <= 0; cloud_xl(22, 25) <= 0; cloud_xl(22, 26) <= 0; cloud_xl(22, 27) <= 0; cloud_xl(22, 28) <= 0; cloud_xl(22, 29) <= 0; cloud_xl(22, 30) <= 0; cloud_xl(22, 31) <= 0; cloud_xl(22, 32) <= 0; cloud_xl(22, 33) <= 0; cloud_xl(22, 34) <= 0; cloud_xl(22, 35) <= 0; cloud_xl(22, 36) <= 0; cloud_xl(22, 37) <= 0; cloud_xl(22, 38) <= 0; cloud_xl(22, 39) <= 0; cloud_xl(22, 40) <= 0; cloud_xl(22, 41) <= 0; cloud_xl(22, 42) <= 0; cloud_xl(22, 43) <= 0; cloud_xl(22, 44) <= 0; cloud_xl(22, 45) <= 0; cloud_xl(22, 46) <= 0; cloud_xl(22, 47) <= 0; cloud_xl(22, 48) <= 0; cloud_xl(22, 49) <= 0; cloud_xl(22, 50) <= 0; cloud_xl(22, 51) <= 0; cloud_xl(22, 52) <= 0; cloud_xl(22, 53) <= 0; cloud_xl(22, 54) <= 0; cloud_xl(22, 55) <= 0; cloud_xl(22, 56) <= 0; cloud_xl(22, 57) <= 0; cloud_xl(22, 58) <= 0; cloud_xl(22, 59) <= 0; cloud_xl(22, 60) <= 1; cloud_xl(22, 61) <= 1; cloud_xl(22, 62) <= 1; cloud_xl(22, 63) <= 1; cloud_xl(22, 64) <= 1; cloud_xl(22, 65) <= 1; cloud_xl(22, 66) <= 1; cloud_xl(22, 67) <= 1; cloud_xl(22, 68) <= 1; cloud_xl(22, 69) <= 1; cloud_xl(22, 70) <= 1; cloud_xl(22, 71) <= 1; cloud_xl(22, 72) <= 2; cloud_xl(22, 73) <= 2; cloud_xl(22, 74) <= 2; cloud_xl(22, 75) <= 2; cloud_xl(22, 76) <= 2; cloud_xl(22, 77) <= 2; 
cloud_xl(23, 0) <= 2; cloud_xl(23, 1) <= 2; cloud_xl(23, 2) <= 2; cloud_xl(23, 3) <= 2; cloud_xl(23, 4) <= 2; cloud_xl(23, 5) <= 2; cloud_xl(23, 6) <= 1; cloud_xl(23, 7) <= 1; cloud_xl(23, 8) <= 1; cloud_xl(23, 9) <= 1; cloud_xl(23, 10) <= 1; cloud_xl(23, 11) <= 1; cloud_xl(23, 12) <= 0; cloud_xl(23, 13) <= 0; cloud_xl(23, 14) <= 0; cloud_xl(23, 15) <= 0; cloud_xl(23, 16) <= 0; cloud_xl(23, 17) <= 0; cloud_xl(23, 18) <= 0; cloud_xl(23, 19) <= 0; cloud_xl(23, 20) <= 0; cloud_xl(23, 21) <= 0; cloud_xl(23, 22) <= 0; cloud_xl(23, 23) <= 0; cloud_xl(23, 24) <= 0; cloud_xl(23, 25) <= 0; cloud_xl(23, 26) <= 0; cloud_xl(23, 27) <= 0; cloud_xl(23, 28) <= 0; cloud_xl(23, 29) <= 0; cloud_xl(23, 30) <= 0; cloud_xl(23, 31) <= 0; cloud_xl(23, 32) <= 0; cloud_xl(23, 33) <= 0; cloud_xl(23, 34) <= 0; cloud_xl(23, 35) <= 0; cloud_xl(23, 36) <= 0; cloud_xl(23, 37) <= 0; cloud_xl(23, 38) <= 0; cloud_xl(23, 39) <= 0; cloud_xl(23, 40) <= 0; cloud_xl(23, 41) <= 0; cloud_xl(23, 42) <= 0; cloud_xl(23, 43) <= 0; cloud_xl(23, 44) <= 0; cloud_xl(23, 45) <= 0; cloud_xl(23, 46) <= 0; cloud_xl(23, 47) <= 0; cloud_xl(23, 48) <= 0; cloud_xl(23, 49) <= 0; cloud_xl(23, 50) <= 0; cloud_xl(23, 51) <= 0; cloud_xl(23, 52) <= 0; cloud_xl(23, 53) <= 0; cloud_xl(23, 54) <= 0; cloud_xl(23, 55) <= 0; cloud_xl(23, 56) <= 0; cloud_xl(23, 57) <= 0; cloud_xl(23, 58) <= 0; cloud_xl(23, 59) <= 0; cloud_xl(23, 60) <= 1; cloud_xl(23, 61) <= 1; cloud_xl(23, 62) <= 1; cloud_xl(23, 63) <= 1; cloud_xl(23, 64) <= 1; cloud_xl(23, 65) <= 1; cloud_xl(23, 66) <= 1; cloud_xl(23, 67) <= 1; cloud_xl(23, 68) <= 1; cloud_xl(23, 69) <= 1; cloud_xl(23, 70) <= 1; cloud_xl(23, 71) <= 1; cloud_xl(23, 72) <= 2; cloud_xl(23, 73) <= 2; cloud_xl(23, 74) <= 2; cloud_xl(23, 75) <= 2; cloud_xl(23, 76) <= 2; cloud_xl(23, 77) <= 2; 
cloud_xl(24, 0) <= 1; cloud_xl(24, 1) <= 1; cloud_xl(24, 2) <= 1; cloud_xl(24, 3) <= 1; cloud_xl(24, 4) <= 1; cloud_xl(24, 5) <= 1; cloud_xl(24, 6) <= 0; cloud_xl(24, 7) <= 0; cloud_xl(24, 8) <= 0; cloud_xl(24, 9) <= 0; cloud_xl(24, 10) <= 0; cloud_xl(24, 11) <= 0; cloud_xl(24, 12) <= 0; cloud_xl(24, 13) <= 0; cloud_xl(24, 14) <= 0; cloud_xl(24, 15) <= 0; cloud_xl(24, 16) <= 0; cloud_xl(24, 17) <= 0; cloud_xl(24, 18) <= 0; cloud_xl(24, 19) <= 0; cloud_xl(24, 20) <= 0; cloud_xl(24, 21) <= 0; cloud_xl(24, 22) <= 0; cloud_xl(24, 23) <= 0; cloud_xl(24, 24) <= 0; cloud_xl(24, 25) <= 0; cloud_xl(24, 26) <= 0; cloud_xl(24, 27) <= 0; cloud_xl(24, 28) <= 0; cloud_xl(24, 29) <= 0; cloud_xl(24, 30) <= 0; cloud_xl(24, 31) <= 0; cloud_xl(24, 32) <= 0; cloud_xl(24, 33) <= 0; cloud_xl(24, 34) <= 0; cloud_xl(24, 35) <= 0; cloud_xl(24, 36) <= 0; cloud_xl(24, 37) <= 0; cloud_xl(24, 38) <= 0; cloud_xl(24, 39) <= 0; cloud_xl(24, 40) <= 0; cloud_xl(24, 41) <= 0; cloud_xl(24, 42) <= 0; cloud_xl(24, 43) <= 0; cloud_xl(24, 44) <= 0; cloud_xl(24, 45) <= 0; cloud_xl(24, 46) <= 0; cloud_xl(24, 47) <= 0; cloud_xl(24, 48) <= 0; cloud_xl(24, 49) <= 0; cloud_xl(24, 50) <= 0; cloud_xl(24, 51) <= 0; cloud_xl(24, 52) <= 0; cloud_xl(24, 53) <= 0; cloud_xl(24, 54) <= 0; cloud_xl(24, 55) <= 0; cloud_xl(24, 56) <= 0; cloud_xl(24, 57) <= 0; cloud_xl(24, 58) <= 0; cloud_xl(24, 59) <= 0; cloud_xl(24, 60) <= 0; cloud_xl(24, 61) <= 0; cloud_xl(24, 62) <= 0; cloud_xl(24, 63) <= 0; cloud_xl(24, 64) <= 0; cloud_xl(24, 65) <= 0; cloud_xl(24, 66) <= 0; cloud_xl(24, 67) <= 0; cloud_xl(24, 68) <= 0; cloud_xl(24, 69) <= 0; cloud_xl(24, 70) <= 0; cloud_xl(24, 71) <= 0; cloud_xl(24, 72) <= 1; cloud_xl(24, 73) <= 1; cloud_xl(24, 74) <= 1; cloud_xl(24, 75) <= 1; cloud_xl(24, 76) <= 1; cloud_xl(24, 77) <= 1; 
cloud_xl(25, 0) <= 1; cloud_xl(25, 1) <= 1; cloud_xl(25, 2) <= 1; cloud_xl(25, 3) <= 1; cloud_xl(25, 4) <= 1; cloud_xl(25, 5) <= 1; cloud_xl(25, 6) <= 0; cloud_xl(25, 7) <= 0; cloud_xl(25, 8) <= 0; cloud_xl(25, 9) <= 0; cloud_xl(25, 10) <= 0; cloud_xl(25, 11) <= 0; cloud_xl(25, 12) <= 0; cloud_xl(25, 13) <= 0; cloud_xl(25, 14) <= 0; cloud_xl(25, 15) <= 0; cloud_xl(25, 16) <= 0; cloud_xl(25, 17) <= 0; cloud_xl(25, 18) <= 0; cloud_xl(25, 19) <= 0; cloud_xl(25, 20) <= 0; cloud_xl(25, 21) <= 0; cloud_xl(25, 22) <= 0; cloud_xl(25, 23) <= 0; cloud_xl(25, 24) <= 0; cloud_xl(25, 25) <= 0; cloud_xl(25, 26) <= 0; cloud_xl(25, 27) <= 0; cloud_xl(25, 28) <= 0; cloud_xl(25, 29) <= 0; cloud_xl(25, 30) <= 0; cloud_xl(25, 31) <= 0; cloud_xl(25, 32) <= 0; cloud_xl(25, 33) <= 0; cloud_xl(25, 34) <= 0; cloud_xl(25, 35) <= 0; cloud_xl(25, 36) <= 0; cloud_xl(25, 37) <= 0; cloud_xl(25, 38) <= 0; cloud_xl(25, 39) <= 0; cloud_xl(25, 40) <= 0; cloud_xl(25, 41) <= 0; cloud_xl(25, 42) <= 0; cloud_xl(25, 43) <= 0; cloud_xl(25, 44) <= 0; cloud_xl(25, 45) <= 0; cloud_xl(25, 46) <= 0; cloud_xl(25, 47) <= 0; cloud_xl(25, 48) <= 0; cloud_xl(25, 49) <= 0; cloud_xl(25, 50) <= 0; cloud_xl(25, 51) <= 0; cloud_xl(25, 52) <= 0; cloud_xl(25, 53) <= 0; cloud_xl(25, 54) <= 0; cloud_xl(25, 55) <= 0; cloud_xl(25, 56) <= 0; cloud_xl(25, 57) <= 0; cloud_xl(25, 58) <= 0; cloud_xl(25, 59) <= 0; cloud_xl(25, 60) <= 0; cloud_xl(25, 61) <= 0; cloud_xl(25, 62) <= 0; cloud_xl(25, 63) <= 0; cloud_xl(25, 64) <= 0; cloud_xl(25, 65) <= 0; cloud_xl(25, 66) <= 0; cloud_xl(25, 67) <= 0; cloud_xl(25, 68) <= 0; cloud_xl(25, 69) <= 0; cloud_xl(25, 70) <= 0; cloud_xl(25, 71) <= 0; cloud_xl(25, 72) <= 1; cloud_xl(25, 73) <= 1; cloud_xl(25, 74) <= 1; cloud_xl(25, 75) <= 1; cloud_xl(25, 76) <= 1; cloud_xl(25, 77) <= 1; 
cloud_xl(26, 0) <= 1; cloud_xl(26, 1) <= 1; cloud_xl(26, 2) <= 1; cloud_xl(26, 3) <= 1; cloud_xl(26, 4) <= 1; cloud_xl(26, 5) <= 1; cloud_xl(26, 6) <= 0; cloud_xl(26, 7) <= 0; cloud_xl(26, 8) <= 0; cloud_xl(26, 9) <= 0; cloud_xl(26, 10) <= 0; cloud_xl(26, 11) <= 0; cloud_xl(26, 12) <= 0; cloud_xl(26, 13) <= 0; cloud_xl(26, 14) <= 0; cloud_xl(26, 15) <= 0; cloud_xl(26, 16) <= 0; cloud_xl(26, 17) <= 0; cloud_xl(26, 18) <= 0; cloud_xl(26, 19) <= 0; cloud_xl(26, 20) <= 0; cloud_xl(26, 21) <= 0; cloud_xl(26, 22) <= 0; cloud_xl(26, 23) <= 0; cloud_xl(26, 24) <= 0; cloud_xl(26, 25) <= 0; cloud_xl(26, 26) <= 0; cloud_xl(26, 27) <= 0; cloud_xl(26, 28) <= 0; cloud_xl(26, 29) <= 0; cloud_xl(26, 30) <= 0; cloud_xl(26, 31) <= 0; cloud_xl(26, 32) <= 0; cloud_xl(26, 33) <= 0; cloud_xl(26, 34) <= 0; cloud_xl(26, 35) <= 0; cloud_xl(26, 36) <= 0; cloud_xl(26, 37) <= 0; cloud_xl(26, 38) <= 0; cloud_xl(26, 39) <= 0; cloud_xl(26, 40) <= 0; cloud_xl(26, 41) <= 0; cloud_xl(26, 42) <= 0; cloud_xl(26, 43) <= 0; cloud_xl(26, 44) <= 0; cloud_xl(26, 45) <= 0; cloud_xl(26, 46) <= 0; cloud_xl(26, 47) <= 0; cloud_xl(26, 48) <= 0; cloud_xl(26, 49) <= 0; cloud_xl(26, 50) <= 0; cloud_xl(26, 51) <= 0; cloud_xl(26, 52) <= 0; cloud_xl(26, 53) <= 0; cloud_xl(26, 54) <= 0; cloud_xl(26, 55) <= 0; cloud_xl(26, 56) <= 0; cloud_xl(26, 57) <= 0; cloud_xl(26, 58) <= 0; cloud_xl(26, 59) <= 0; cloud_xl(26, 60) <= 0; cloud_xl(26, 61) <= 0; cloud_xl(26, 62) <= 0; cloud_xl(26, 63) <= 0; cloud_xl(26, 64) <= 0; cloud_xl(26, 65) <= 0; cloud_xl(26, 66) <= 0; cloud_xl(26, 67) <= 0; cloud_xl(26, 68) <= 0; cloud_xl(26, 69) <= 0; cloud_xl(26, 70) <= 0; cloud_xl(26, 71) <= 0; cloud_xl(26, 72) <= 1; cloud_xl(26, 73) <= 1; cloud_xl(26, 74) <= 1; cloud_xl(26, 75) <= 1; cloud_xl(26, 76) <= 1; cloud_xl(26, 77) <= 1; 
cloud_xl(27, 0) <= 1; cloud_xl(27, 1) <= 1; cloud_xl(27, 2) <= 1; cloud_xl(27, 3) <= 1; cloud_xl(27, 4) <= 1; cloud_xl(27, 5) <= 1; cloud_xl(27, 6) <= 0; cloud_xl(27, 7) <= 0; cloud_xl(27, 8) <= 0; cloud_xl(27, 9) <= 0; cloud_xl(27, 10) <= 0; cloud_xl(27, 11) <= 0; cloud_xl(27, 12) <= 0; cloud_xl(27, 13) <= 0; cloud_xl(27, 14) <= 0; cloud_xl(27, 15) <= 0; cloud_xl(27, 16) <= 0; cloud_xl(27, 17) <= 0; cloud_xl(27, 18) <= 0; cloud_xl(27, 19) <= 0; cloud_xl(27, 20) <= 0; cloud_xl(27, 21) <= 0; cloud_xl(27, 22) <= 0; cloud_xl(27, 23) <= 0; cloud_xl(27, 24) <= 0; cloud_xl(27, 25) <= 0; cloud_xl(27, 26) <= 0; cloud_xl(27, 27) <= 0; cloud_xl(27, 28) <= 0; cloud_xl(27, 29) <= 0; cloud_xl(27, 30) <= 0; cloud_xl(27, 31) <= 0; cloud_xl(27, 32) <= 0; cloud_xl(27, 33) <= 0; cloud_xl(27, 34) <= 0; cloud_xl(27, 35) <= 0; cloud_xl(27, 36) <= 0; cloud_xl(27, 37) <= 0; cloud_xl(27, 38) <= 0; cloud_xl(27, 39) <= 0; cloud_xl(27, 40) <= 0; cloud_xl(27, 41) <= 0; cloud_xl(27, 42) <= 0; cloud_xl(27, 43) <= 0; cloud_xl(27, 44) <= 0; cloud_xl(27, 45) <= 0; cloud_xl(27, 46) <= 0; cloud_xl(27, 47) <= 0; cloud_xl(27, 48) <= 0; cloud_xl(27, 49) <= 0; cloud_xl(27, 50) <= 0; cloud_xl(27, 51) <= 0; cloud_xl(27, 52) <= 0; cloud_xl(27, 53) <= 0; cloud_xl(27, 54) <= 0; cloud_xl(27, 55) <= 0; cloud_xl(27, 56) <= 0; cloud_xl(27, 57) <= 0; cloud_xl(27, 58) <= 0; cloud_xl(27, 59) <= 0; cloud_xl(27, 60) <= 0; cloud_xl(27, 61) <= 0; cloud_xl(27, 62) <= 0; cloud_xl(27, 63) <= 0; cloud_xl(27, 64) <= 0; cloud_xl(27, 65) <= 0; cloud_xl(27, 66) <= 0; cloud_xl(27, 67) <= 0; cloud_xl(27, 68) <= 0; cloud_xl(27, 69) <= 0; cloud_xl(27, 70) <= 0; cloud_xl(27, 71) <= 0; cloud_xl(27, 72) <= 1; cloud_xl(27, 73) <= 1; cloud_xl(27, 74) <= 1; cloud_xl(27, 75) <= 1; cloud_xl(27, 76) <= 1; cloud_xl(27, 77) <= 1; 
cloud_xl(28, 0) <= 1; cloud_xl(28, 1) <= 1; cloud_xl(28, 2) <= 1; cloud_xl(28, 3) <= 1; cloud_xl(28, 4) <= 1; cloud_xl(28, 5) <= 1; cloud_xl(28, 6) <= 0; cloud_xl(28, 7) <= 0; cloud_xl(28, 8) <= 0; cloud_xl(28, 9) <= 0; cloud_xl(28, 10) <= 0; cloud_xl(28, 11) <= 0; cloud_xl(28, 12) <= 0; cloud_xl(28, 13) <= 0; cloud_xl(28, 14) <= 0; cloud_xl(28, 15) <= 0; cloud_xl(28, 16) <= 0; cloud_xl(28, 17) <= 0; cloud_xl(28, 18) <= 0; cloud_xl(28, 19) <= 0; cloud_xl(28, 20) <= 0; cloud_xl(28, 21) <= 0; cloud_xl(28, 22) <= 0; cloud_xl(28, 23) <= 0; cloud_xl(28, 24) <= 0; cloud_xl(28, 25) <= 0; cloud_xl(28, 26) <= 0; cloud_xl(28, 27) <= 0; cloud_xl(28, 28) <= 0; cloud_xl(28, 29) <= 0; cloud_xl(28, 30) <= 0; cloud_xl(28, 31) <= 0; cloud_xl(28, 32) <= 0; cloud_xl(28, 33) <= 0; cloud_xl(28, 34) <= 0; cloud_xl(28, 35) <= 0; cloud_xl(28, 36) <= 0; cloud_xl(28, 37) <= 0; cloud_xl(28, 38) <= 0; cloud_xl(28, 39) <= 0; cloud_xl(28, 40) <= 0; cloud_xl(28, 41) <= 0; cloud_xl(28, 42) <= 0; cloud_xl(28, 43) <= 0; cloud_xl(28, 44) <= 0; cloud_xl(28, 45) <= 0; cloud_xl(28, 46) <= 0; cloud_xl(28, 47) <= 0; cloud_xl(28, 48) <= 0; cloud_xl(28, 49) <= 0; cloud_xl(28, 50) <= 0; cloud_xl(28, 51) <= 0; cloud_xl(28, 52) <= 0; cloud_xl(28, 53) <= 0; cloud_xl(28, 54) <= 0; cloud_xl(28, 55) <= 0; cloud_xl(28, 56) <= 0; cloud_xl(28, 57) <= 0; cloud_xl(28, 58) <= 0; cloud_xl(28, 59) <= 0; cloud_xl(28, 60) <= 0; cloud_xl(28, 61) <= 0; cloud_xl(28, 62) <= 0; cloud_xl(28, 63) <= 0; cloud_xl(28, 64) <= 0; cloud_xl(28, 65) <= 0; cloud_xl(28, 66) <= 0; cloud_xl(28, 67) <= 0; cloud_xl(28, 68) <= 0; cloud_xl(28, 69) <= 0; cloud_xl(28, 70) <= 0; cloud_xl(28, 71) <= 0; cloud_xl(28, 72) <= 1; cloud_xl(28, 73) <= 1; cloud_xl(28, 74) <= 1; cloud_xl(28, 75) <= 1; cloud_xl(28, 76) <= 1; cloud_xl(28, 77) <= 1; 
cloud_xl(29, 0) <= 1; cloud_xl(29, 1) <= 1; cloud_xl(29, 2) <= 1; cloud_xl(29, 3) <= 1; cloud_xl(29, 4) <= 1; cloud_xl(29, 5) <= 1; cloud_xl(29, 6) <= 0; cloud_xl(29, 7) <= 0; cloud_xl(29, 8) <= 0; cloud_xl(29, 9) <= 0; cloud_xl(29, 10) <= 0; cloud_xl(29, 11) <= 0; cloud_xl(29, 12) <= 0; cloud_xl(29, 13) <= 0; cloud_xl(29, 14) <= 0; cloud_xl(29, 15) <= 0; cloud_xl(29, 16) <= 0; cloud_xl(29, 17) <= 0; cloud_xl(29, 18) <= 0; cloud_xl(29, 19) <= 0; cloud_xl(29, 20) <= 0; cloud_xl(29, 21) <= 0; cloud_xl(29, 22) <= 0; cloud_xl(29, 23) <= 0; cloud_xl(29, 24) <= 0; cloud_xl(29, 25) <= 0; cloud_xl(29, 26) <= 0; cloud_xl(29, 27) <= 0; cloud_xl(29, 28) <= 0; cloud_xl(29, 29) <= 0; cloud_xl(29, 30) <= 0; cloud_xl(29, 31) <= 0; cloud_xl(29, 32) <= 0; cloud_xl(29, 33) <= 0; cloud_xl(29, 34) <= 0; cloud_xl(29, 35) <= 0; cloud_xl(29, 36) <= 0; cloud_xl(29, 37) <= 0; cloud_xl(29, 38) <= 0; cloud_xl(29, 39) <= 0; cloud_xl(29, 40) <= 0; cloud_xl(29, 41) <= 0; cloud_xl(29, 42) <= 0; cloud_xl(29, 43) <= 0; cloud_xl(29, 44) <= 0; cloud_xl(29, 45) <= 0; cloud_xl(29, 46) <= 0; cloud_xl(29, 47) <= 0; cloud_xl(29, 48) <= 0; cloud_xl(29, 49) <= 0; cloud_xl(29, 50) <= 0; cloud_xl(29, 51) <= 0; cloud_xl(29, 52) <= 0; cloud_xl(29, 53) <= 0; cloud_xl(29, 54) <= 0; cloud_xl(29, 55) <= 0; cloud_xl(29, 56) <= 0; cloud_xl(29, 57) <= 0; cloud_xl(29, 58) <= 0; cloud_xl(29, 59) <= 0; cloud_xl(29, 60) <= 0; cloud_xl(29, 61) <= 0; cloud_xl(29, 62) <= 0; cloud_xl(29, 63) <= 0; cloud_xl(29, 64) <= 0; cloud_xl(29, 65) <= 0; cloud_xl(29, 66) <= 0; cloud_xl(29, 67) <= 0; cloud_xl(29, 68) <= 0; cloud_xl(29, 69) <= 0; cloud_xl(29, 70) <= 0; cloud_xl(29, 71) <= 0; cloud_xl(29, 72) <= 1; cloud_xl(29, 73) <= 1; cloud_xl(29, 74) <= 1; cloud_xl(29, 75) <= 1; cloud_xl(29, 76) <= 1; cloud_xl(29, 77) <= 1; 
cloud_xl(30, 0) <= 1; cloud_xl(30, 1) <= 1; cloud_xl(30, 2) <= 1; cloud_xl(30, 3) <= 1; cloud_xl(30, 4) <= 1; cloud_xl(30, 5) <= 1; cloud_xl(30, 6) <= 0; cloud_xl(30, 7) <= 0; cloud_xl(30, 8) <= 0; cloud_xl(30, 9) <= 0; cloud_xl(30, 10) <= 0; cloud_xl(30, 11) <= 0; cloud_xl(30, 12) <= 0; cloud_xl(30, 13) <= 0; cloud_xl(30, 14) <= 0; cloud_xl(30, 15) <= 0; cloud_xl(30, 16) <= 0; cloud_xl(30, 17) <= 0; cloud_xl(30, 18) <= 0; cloud_xl(30, 19) <= 0; cloud_xl(30, 20) <= 0; cloud_xl(30, 21) <= 0; cloud_xl(30, 22) <= 0; cloud_xl(30, 23) <= 0; cloud_xl(30, 24) <= 0; cloud_xl(30, 25) <= 0; cloud_xl(30, 26) <= 0; cloud_xl(30, 27) <= 0; cloud_xl(30, 28) <= 0; cloud_xl(30, 29) <= 0; cloud_xl(30, 30) <= 0; cloud_xl(30, 31) <= 0; cloud_xl(30, 32) <= 0; cloud_xl(30, 33) <= 0; cloud_xl(30, 34) <= 0; cloud_xl(30, 35) <= 0; cloud_xl(30, 36) <= 0; cloud_xl(30, 37) <= 0; cloud_xl(30, 38) <= 0; cloud_xl(30, 39) <= 0; cloud_xl(30, 40) <= 0; cloud_xl(30, 41) <= 0; cloud_xl(30, 42) <= 0; cloud_xl(30, 43) <= 0; cloud_xl(30, 44) <= 0; cloud_xl(30, 45) <= 0; cloud_xl(30, 46) <= 0; cloud_xl(30, 47) <= 0; cloud_xl(30, 48) <= 0; cloud_xl(30, 49) <= 0; cloud_xl(30, 50) <= 0; cloud_xl(30, 51) <= 0; cloud_xl(30, 52) <= 0; cloud_xl(30, 53) <= 0; cloud_xl(30, 54) <= 0; cloud_xl(30, 55) <= 0; cloud_xl(30, 56) <= 0; cloud_xl(30, 57) <= 0; cloud_xl(30, 58) <= 0; cloud_xl(30, 59) <= 0; cloud_xl(30, 60) <= 0; cloud_xl(30, 61) <= 0; cloud_xl(30, 62) <= 0; cloud_xl(30, 63) <= 0; cloud_xl(30, 64) <= 0; cloud_xl(30, 65) <= 0; cloud_xl(30, 66) <= 0; cloud_xl(30, 67) <= 0; cloud_xl(30, 68) <= 0; cloud_xl(30, 69) <= 0; cloud_xl(30, 70) <= 0; cloud_xl(30, 71) <= 0; cloud_xl(30, 72) <= 1; cloud_xl(30, 73) <= 1; cloud_xl(30, 74) <= 1; cloud_xl(30, 75) <= 1; cloud_xl(30, 76) <= 1; cloud_xl(30, 77) <= 1; 
cloud_xl(31, 0) <= 1; cloud_xl(31, 1) <= 1; cloud_xl(31, 2) <= 1; cloud_xl(31, 3) <= 1; cloud_xl(31, 4) <= 1; cloud_xl(31, 5) <= 1; cloud_xl(31, 6) <= 0; cloud_xl(31, 7) <= 0; cloud_xl(31, 8) <= 0; cloud_xl(31, 9) <= 0; cloud_xl(31, 10) <= 0; cloud_xl(31, 11) <= 0; cloud_xl(31, 12) <= 0; cloud_xl(31, 13) <= 0; cloud_xl(31, 14) <= 0; cloud_xl(31, 15) <= 0; cloud_xl(31, 16) <= 0; cloud_xl(31, 17) <= 0; cloud_xl(31, 18) <= 0; cloud_xl(31, 19) <= 0; cloud_xl(31, 20) <= 0; cloud_xl(31, 21) <= 0; cloud_xl(31, 22) <= 0; cloud_xl(31, 23) <= 0; cloud_xl(31, 24) <= 0; cloud_xl(31, 25) <= 0; cloud_xl(31, 26) <= 0; cloud_xl(31, 27) <= 0; cloud_xl(31, 28) <= 0; cloud_xl(31, 29) <= 0; cloud_xl(31, 30) <= 0; cloud_xl(31, 31) <= 0; cloud_xl(31, 32) <= 0; cloud_xl(31, 33) <= 0; cloud_xl(31, 34) <= 0; cloud_xl(31, 35) <= 0; cloud_xl(31, 36) <= 0; cloud_xl(31, 37) <= 0; cloud_xl(31, 38) <= 0; cloud_xl(31, 39) <= 0; cloud_xl(31, 40) <= 0; cloud_xl(31, 41) <= 0; cloud_xl(31, 42) <= 0; cloud_xl(31, 43) <= 0; cloud_xl(31, 44) <= 0; cloud_xl(31, 45) <= 0; cloud_xl(31, 46) <= 0; cloud_xl(31, 47) <= 0; cloud_xl(31, 48) <= 0; cloud_xl(31, 49) <= 0; cloud_xl(31, 50) <= 0; cloud_xl(31, 51) <= 0; cloud_xl(31, 52) <= 0; cloud_xl(31, 53) <= 0; cloud_xl(31, 54) <= 0; cloud_xl(31, 55) <= 0; cloud_xl(31, 56) <= 0; cloud_xl(31, 57) <= 0; cloud_xl(31, 58) <= 0; cloud_xl(31, 59) <= 0; cloud_xl(31, 60) <= 0; cloud_xl(31, 61) <= 0; cloud_xl(31, 62) <= 0; cloud_xl(31, 63) <= 0; cloud_xl(31, 64) <= 0; cloud_xl(31, 65) <= 0; cloud_xl(31, 66) <= 0; cloud_xl(31, 67) <= 0; cloud_xl(31, 68) <= 0; cloud_xl(31, 69) <= 0; cloud_xl(31, 70) <= 0; cloud_xl(31, 71) <= 0; cloud_xl(31, 72) <= 1; cloud_xl(31, 73) <= 1; cloud_xl(31, 74) <= 1; cloud_xl(31, 75) <= 1; cloud_xl(31, 76) <= 1; cloud_xl(31, 77) <= 1; 
cloud_xl(32, 0) <= 1; cloud_xl(32, 1) <= 1; cloud_xl(32, 2) <= 1; cloud_xl(32, 3) <= 1; cloud_xl(32, 4) <= 1; cloud_xl(32, 5) <= 1; cloud_xl(32, 6) <= 0; cloud_xl(32, 7) <= 0; cloud_xl(32, 8) <= 0; cloud_xl(32, 9) <= 0; cloud_xl(32, 10) <= 0; cloud_xl(32, 11) <= 0; cloud_xl(32, 12) <= 0; cloud_xl(32, 13) <= 0; cloud_xl(32, 14) <= 0; cloud_xl(32, 15) <= 0; cloud_xl(32, 16) <= 0; cloud_xl(32, 17) <= 0; cloud_xl(32, 18) <= 0; cloud_xl(32, 19) <= 0; cloud_xl(32, 20) <= 0; cloud_xl(32, 21) <= 0; cloud_xl(32, 22) <= 0; cloud_xl(32, 23) <= 0; cloud_xl(32, 24) <= 0; cloud_xl(32, 25) <= 0; cloud_xl(32, 26) <= 0; cloud_xl(32, 27) <= 0; cloud_xl(32, 28) <= 0; cloud_xl(32, 29) <= 0; cloud_xl(32, 30) <= 0; cloud_xl(32, 31) <= 0; cloud_xl(32, 32) <= 0; cloud_xl(32, 33) <= 0; cloud_xl(32, 34) <= 0; cloud_xl(32, 35) <= 0; cloud_xl(32, 36) <= 0; cloud_xl(32, 37) <= 0; cloud_xl(32, 38) <= 0; cloud_xl(32, 39) <= 0; cloud_xl(32, 40) <= 0; cloud_xl(32, 41) <= 0; cloud_xl(32, 42) <= 0; cloud_xl(32, 43) <= 0; cloud_xl(32, 44) <= 0; cloud_xl(32, 45) <= 0; cloud_xl(32, 46) <= 0; cloud_xl(32, 47) <= 0; cloud_xl(32, 48) <= 0; cloud_xl(32, 49) <= 0; cloud_xl(32, 50) <= 0; cloud_xl(32, 51) <= 0; cloud_xl(32, 52) <= 0; cloud_xl(32, 53) <= 0; cloud_xl(32, 54) <= 0; cloud_xl(32, 55) <= 0; cloud_xl(32, 56) <= 0; cloud_xl(32, 57) <= 0; cloud_xl(32, 58) <= 0; cloud_xl(32, 59) <= 0; cloud_xl(32, 60) <= 0; cloud_xl(32, 61) <= 0; cloud_xl(32, 62) <= 0; cloud_xl(32, 63) <= 0; cloud_xl(32, 64) <= 0; cloud_xl(32, 65) <= 0; cloud_xl(32, 66) <= 0; cloud_xl(32, 67) <= 0; cloud_xl(32, 68) <= 0; cloud_xl(32, 69) <= 0; cloud_xl(32, 70) <= 0; cloud_xl(32, 71) <= 0; cloud_xl(32, 72) <= 1; cloud_xl(32, 73) <= 1; cloud_xl(32, 74) <= 1; cloud_xl(32, 75) <= 1; cloud_xl(32, 76) <= 1; cloud_xl(32, 77) <= 1; 
cloud_xl(33, 0) <= 1; cloud_xl(33, 1) <= 1; cloud_xl(33, 2) <= 1; cloud_xl(33, 3) <= 1; cloud_xl(33, 4) <= 1; cloud_xl(33, 5) <= 1; cloud_xl(33, 6) <= 0; cloud_xl(33, 7) <= 0; cloud_xl(33, 8) <= 0; cloud_xl(33, 9) <= 0; cloud_xl(33, 10) <= 0; cloud_xl(33, 11) <= 0; cloud_xl(33, 12) <= 0; cloud_xl(33, 13) <= 0; cloud_xl(33, 14) <= 0; cloud_xl(33, 15) <= 0; cloud_xl(33, 16) <= 0; cloud_xl(33, 17) <= 0; cloud_xl(33, 18) <= 0; cloud_xl(33, 19) <= 0; cloud_xl(33, 20) <= 0; cloud_xl(33, 21) <= 0; cloud_xl(33, 22) <= 0; cloud_xl(33, 23) <= 0; cloud_xl(33, 24) <= 0; cloud_xl(33, 25) <= 0; cloud_xl(33, 26) <= 0; cloud_xl(33, 27) <= 0; cloud_xl(33, 28) <= 0; cloud_xl(33, 29) <= 0; cloud_xl(33, 30) <= 0; cloud_xl(33, 31) <= 0; cloud_xl(33, 32) <= 0; cloud_xl(33, 33) <= 0; cloud_xl(33, 34) <= 0; cloud_xl(33, 35) <= 0; cloud_xl(33, 36) <= 0; cloud_xl(33, 37) <= 0; cloud_xl(33, 38) <= 0; cloud_xl(33, 39) <= 0; cloud_xl(33, 40) <= 0; cloud_xl(33, 41) <= 0; cloud_xl(33, 42) <= 0; cloud_xl(33, 43) <= 0; cloud_xl(33, 44) <= 0; cloud_xl(33, 45) <= 0; cloud_xl(33, 46) <= 0; cloud_xl(33, 47) <= 0; cloud_xl(33, 48) <= 0; cloud_xl(33, 49) <= 0; cloud_xl(33, 50) <= 0; cloud_xl(33, 51) <= 0; cloud_xl(33, 52) <= 0; cloud_xl(33, 53) <= 0; cloud_xl(33, 54) <= 0; cloud_xl(33, 55) <= 0; cloud_xl(33, 56) <= 0; cloud_xl(33, 57) <= 0; cloud_xl(33, 58) <= 0; cloud_xl(33, 59) <= 0; cloud_xl(33, 60) <= 0; cloud_xl(33, 61) <= 0; cloud_xl(33, 62) <= 0; cloud_xl(33, 63) <= 0; cloud_xl(33, 64) <= 0; cloud_xl(33, 65) <= 0; cloud_xl(33, 66) <= 0; cloud_xl(33, 67) <= 0; cloud_xl(33, 68) <= 0; cloud_xl(33, 69) <= 0; cloud_xl(33, 70) <= 0; cloud_xl(33, 71) <= 0; cloud_xl(33, 72) <= 1; cloud_xl(33, 73) <= 1; cloud_xl(33, 74) <= 1; cloud_xl(33, 75) <= 1; cloud_xl(33, 76) <= 1; cloud_xl(33, 77) <= 1; 
cloud_xl(34, 0) <= 1; cloud_xl(34, 1) <= 1; cloud_xl(34, 2) <= 1; cloud_xl(34, 3) <= 1; cloud_xl(34, 4) <= 1; cloud_xl(34, 5) <= 1; cloud_xl(34, 6) <= 0; cloud_xl(34, 7) <= 0; cloud_xl(34, 8) <= 0; cloud_xl(34, 9) <= 0; cloud_xl(34, 10) <= 0; cloud_xl(34, 11) <= 0; cloud_xl(34, 12) <= 0; cloud_xl(34, 13) <= 0; cloud_xl(34, 14) <= 0; cloud_xl(34, 15) <= 0; cloud_xl(34, 16) <= 0; cloud_xl(34, 17) <= 0; cloud_xl(34, 18) <= 0; cloud_xl(34, 19) <= 0; cloud_xl(34, 20) <= 0; cloud_xl(34, 21) <= 0; cloud_xl(34, 22) <= 0; cloud_xl(34, 23) <= 0; cloud_xl(34, 24) <= 0; cloud_xl(34, 25) <= 0; cloud_xl(34, 26) <= 0; cloud_xl(34, 27) <= 0; cloud_xl(34, 28) <= 0; cloud_xl(34, 29) <= 0; cloud_xl(34, 30) <= 0; cloud_xl(34, 31) <= 0; cloud_xl(34, 32) <= 0; cloud_xl(34, 33) <= 0; cloud_xl(34, 34) <= 0; cloud_xl(34, 35) <= 0; cloud_xl(34, 36) <= 0; cloud_xl(34, 37) <= 0; cloud_xl(34, 38) <= 0; cloud_xl(34, 39) <= 0; cloud_xl(34, 40) <= 0; cloud_xl(34, 41) <= 0; cloud_xl(34, 42) <= 0; cloud_xl(34, 43) <= 0; cloud_xl(34, 44) <= 0; cloud_xl(34, 45) <= 0; cloud_xl(34, 46) <= 0; cloud_xl(34, 47) <= 0; cloud_xl(34, 48) <= 0; cloud_xl(34, 49) <= 0; cloud_xl(34, 50) <= 0; cloud_xl(34, 51) <= 0; cloud_xl(34, 52) <= 0; cloud_xl(34, 53) <= 0; cloud_xl(34, 54) <= 0; cloud_xl(34, 55) <= 0; cloud_xl(34, 56) <= 0; cloud_xl(34, 57) <= 0; cloud_xl(34, 58) <= 0; cloud_xl(34, 59) <= 0; cloud_xl(34, 60) <= 0; cloud_xl(34, 61) <= 0; cloud_xl(34, 62) <= 0; cloud_xl(34, 63) <= 0; cloud_xl(34, 64) <= 0; cloud_xl(34, 65) <= 0; cloud_xl(34, 66) <= 0; cloud_xl(34, 67) <= 0; cloud_xl(34, 68) <= 0; cloud_xl(34, 69) <= 0; cloud_xl(34, 70) <= 0; cloud_xl(34, 71) <= 0; cloud_xl(34, 72) <= 1; cloud_xl(34, 73) <= 1; cloud_xl(34, 74) <= 1; cloud_xl(34, 75) <= 1; cloud_xl(34, 76) <= 1; cloud_xl(34, 77) <= 1; 
cloud_xl(35, 0) <= 1; cloud_xl(35, 1) <= 1; cloud_xl(35, 2) <= 1; cloud_xl(35, 3) <= 1; cloud_xl(35, 4) <= 1; cloud_xl(35, 5) <= 1; cloud_xl(35, 6) <= 0; cloud_xl(35, 7) <= 0; cloud_xl(35, 8) <= 0; cloud_xl(35, 9) <= 0; cloud_xl(35, 10) <= 0; cloud_xl(35, 11) <= 0; cloud_xl(35, 12) <= 0; cloud_xl(35, 13) <= 0; cloud_xl(35, 14) <= 0; cloud_xl(35, 15) <= 0; cloud_xl(35, 16) <= 0; cloud_xl(35, 17) <= 0; cloud_xl(35, 18) <= 0; cloud_xl(35, 19) <= 0; cloud_xl(35, 20) <= 0; cloud_xl(35, 21) <= 0; cloud_xl(35, 22) <= 0; cloud_xl(35, 23) <= 0; cloud_xl(35, 24) <= 0; cloud_xl(35, 25) <= 0; cloud_xl(35, 26) <= 0; cloud_xl(35, 27) <= 0; cloud_xl(35, 28) <= 0; cloud_xl(35, 29) <= 0; cloud_xl(35, 30) <= 0; cloud_xl(35, 31) <= 0; cloud_xl(35, 32) <= 0; cloud_xl(35, 33) <= 0; cloud_xl(35, 34) <= 0; cloud_xl(35, 35) <= 0; cloud_xl(35, 36) <= 0; cloud_xl(35, 37) <= 0; cloud_xl(35, 38) <= 0; cloud_xl(35, 39) <= 0; cloud_xl(35, 40) <= 0; cloud_xl(35, 41) <= 0; cloud_xl(35, 42) <= 0; cloud_xl(35, 43) <= 0; cloud_xl(35, 44) <= 0; cloud_xl(35, 45) <= 0; cloud_xl(35, 46) <= 0; cloud_xl(35, 47) <= 0; cloud_xl(35, 48) <= 0; cloud_xl(35, 49) <= 0; cloud_xl(35, 50) <= 0; cloud_xl(35, 51) <= 0; cloud_xl(35, 52) <= 0; cloud_xl(35, 53) <= 0; cloud_xl(35, 54) <= 0; cloud_xl(35, 55) <= 0; cloud_xl(35, 56) <= 0; cloud_xl(35, 57) <= 0; cloud_xl(35, 58) <= 0; cloud_xl(35, 59) <= 0; cloud_xl(35, 60) <= 0; cloud_xl(35, 61) <= 0; cloud_xl(35, 62) <= 0; cloud_xl(35, 63) <= 0; cloud_xl(35, 64) <= 0; cloud_xl(35, 65) <= 0; cloud_xl(35, 66) <= 0; cloud_xl(35, 67) <= 0; cloud_xl(35, 68) <= 0; cloud_xl(35, 69) <= 0; cloud_xl(35, 70) <= 0; cloud_xl(35, 71) <= 0; cloud_xl(35, 72) <= 1; cloud_xl(35, 73) <= 1; cloud_xl(35, 74) <= 1; cloud_xl(35, 75) <= 1; cloud_xl(35, 76) <= 1; cloud_xl(35, 77) <= 1; 
cloud_xl(36, 0) <= 1; cloud_xl(36, 1) <= 1; cloud_xl(36, 2) <= 1; cloud_xl(36, 3) <= 1; cloud_xl(36, 4) <= 1; cloud_xl(36, 5) <= 1; cloud_xl(36, 6) <= 0; cloud_xl(36, 7) <= 0; cloud_xl(36, 8) <= 0; cloud_xl(36, 9) <= 0; cloud_xl(36, 10) <= 0; cloud_xl(36, 11) <= 0; cloud_xl(36, 12) <= 0; cloud_xl(36, 13) <= 0; cloud_xl(36, 14) <= 0; cloud_xl(36, 15) <= 0; cloud_xl(36, 16) <= 0; cloud_xl(36, 17) <= 0; cloud_xl(36, 18) <= 0; cloud_xl(36, 19) <= 0; cloud_xl(36, 20) <= 0; cloud_xl(36, 21) <= 0; cloud_xl(36, 22) <= 0; cloud_xl(36, 23) <= 0; cloud_xl(36, 24) <= 0; cloud_xl(36, 25) <= 0; cloud_xl(36, 26) <= 0; cloud_xl(36, 27) <= 0; cloud_xl(36, 28) <= 0; cloud_xl(36, 29) <= 0; cloud_xl(36, 30) <= 0; cloud_xl(36, 31) <= 0; cloud_xl(36, 32) <= 0; cloud_xl(36, 33) <= 0; cloud_xl(36, 34) <= 0; cloud_xl(36, 35) <= 0; cloud_xl(36, 36) <= 0; cloud_xl(36, 37) <= 0; cloud_xl(36, 38) <= 0; cloud_xl(36, 39) <= 0; cloud_xl(36, 40) <= 0; cloud_xl(36, 41) <= 0; cloud_xl(36, 42) <= 0; cloud_xl(36, 43) <= 0; cloud_xl(36, 44) <= 0; cloud_xl(36, 45) <= 0; cloud_xl(36, 46) <= 0; cloud_xl(36, 47) <= 0; cloud_xl(36, 48) <= 0; cloud_xl(36, 49) <= 0; cloud_xl(36, 50) <= 0; cloud_xl(36, 51) <= 0; cloud_xl(36, 52) <= 0; cloud_xl(36, 53) <= 0; cloud_xl(36, 54) <= 0; cloud_xl(36, 55) <= 0; cloud_xl(36, 56) <= 0; cloud_xl(36, 57) <= 0; cloud_xl(36, 58) <= 0; cloud_xl(36, 59) <= 0; cloud_xl(36, 60) <= 0; cloud_xl(36, 61) <= 0; cloud_xl(36, 62) <= 0; cloud_xl(36, 63) <= 0; cloud_xl(36, 64) <= 0; cloud_xl(36, 65) <= 0; cloud_xl(36, 66) <= 0; cloud_xl(36, 67) <= 0; cloud_xl(36, 68) <= 0; cloud_xl(36, 69) <= 0; cloud_xl(36, 70) <= 0; cloud_xl(36, 71) <= 0; cloud_xl(36, 72) <= 1; cloud_xl(36, 73) <= 1; cloud_xl(36, 74) <= 1; cloud_xl(36, 75) <= 1; cloud_xl(36, 76) <= 1; cloud_xl(36, 77) <= 1; 
cloud_xl(37, 0) <= 1; cloud_xl(37, 1) <= 1; cloud_xl(37, 2) <= 1; cloud_xl(37, 3) <= 1; cloud_xl(37, 4) <= 1; cloud_xl(37, 5) <= 1; cloud_xl(37, 6) <= 0; cloud_xl(37, 7) <= 0; cloud_xl(37, 8) <= 0; cloud_xl(37, 9) <= 0; cloud_xl(37, 10) <= 0; cloud_xl(37, 11) <= 0; cloud_xl(37, 12) <= 0; cloud_xl(37, 13) <= 0; cloud_xl(37, 14) <= 0; cloud_xl(37, 15) <= 0; cloud_xl(37, 16) <= 0; cloud_xl(37, 17) <= 0; cloud_xl(37, 18) <= 0; cloud_xl(37, 19) <= 0; cloud_xl(37, 20) <= 0; cloud_xl(37, 21) <= 0; cloud_xl(37, 22) <= 0; cloud_xl(37, 23) <= 0; cloud_xl(37, 24) <= 0; cloud_xl(37, 25) <= 0; cloud_xl(37, 26) <= 0; cloud_xl(37, 27) <= 0; cloud_xl(37, 28) <= 0; cloud_xl(37, 29) <= 0; cloud_xl(37, 30) <= 0; cloud_xl(37, 31) <= 0; cloud_xl(37, 32) <= 0; cloud_xl(37, 33) <= 0; cloud_xl(37, 34) <= 0; cloud_xl(37, 35) <= 0; cloud_xl(37, 36) <= 0; cloud_xl(37, 37) <= 0; cloud_xl(37, 38) <= 0; cloud_xl(37, 39) <= 0; cloud_xl(37, 40) <= 0; cloud_xl(37, 41) <= 0; cloud_xl(37, 42) <= 0; cloud_xl(37, 43) <= 0; cloud_xl(37, 44) <= 0; cloud_xl(37, 45) <= 0; cloud_xl(37, 46) <= 0; cloud_xl(37, 47) <= 0; cloud_xl(37, 48) <= 0; cloud_xl(37, 49) <= 0; cloud_xl(37, 50) <= 0; cloud_xl(37, 51) <= 0; cloud_xl(37, 52) <= 0; cloud_xl(37, 53) <= 0; cloud_xl(37, 54) <= 0; cloud_xl(37, 55) <= 0; cloud_xl(37, 56) <= 0; cloud_xl(37, 57) <= 0; cloud_xl(37, 58) <= 0; cloud_xl(37, 59) <= 0; cloud_xl(37, 60) <= 0; cloud_xl(37, 61) <= 0; cloud_xl(37, 62) <= 0; cloud_xl(37, 63) <= 0; cloud_xl(37, 64) <= 0; cloud_xl(37, 65) <= 0; cloud_xl(37, 66) <= 0; cloud_xl(37, 67) <= 0; cloud_xl(37, 68) <= 0; cloud_xl(37, 69) <= 0; cloud_xl(37, 70) <= 0; cloud_xl(37, 71) <= 0; cloud_xl(37, 72) <= 1; cloud_xl(37, 73) <= 1; cloud_xl(37, 74) <= 1; cloud_xl(37, 75) <= 1; cloud_xl(37, 76) <= 1; cloud_xl(37, 77) <= 1; 
cloud_xl(38, 0) <= 1; cloud_xl(38, 1) <= 1; cloud_xl(38, 2) <= 1; cloud_xl(38, 3) <= 1; cloud_xl(38, 4) <= 1; cloud_xl(38, 5) <= 1; cloud_xl(38, 6) <= 0; cloud_xl(38, 7) <= 0; cloud_xl(38, 8) <= 0; cloud_xl(38, 9) <= 0; cloud_xl(38, 10) <= 0; cloud_xl(38, 11) <= 0; cloud_xl(38, 12) <= 0; cloud_xl(38, 13) <= 0; cloud_xl(38, 14) <= 0; cloud_xl(38, 15) <= 0; cloud_xl(38, 16) <= 0; cloud_xl(38, 17) <= 0; cloud_xl(38, 18) <= 0; cloud_xl(38, 19) <= 0; cloud_xl(38, 20) <= 0; cloud_xl(38, 21) <= 0; cloud_xl(38, 22) <= 0; cloud_xl(38, 23) <= 0; cloud_xl(38, 24) <= 0; cloud_xl(38, 25) <= 0; cloud_xl(38, 26) <= 0; cloud_xl(38, 27) <= 0; cloud_xl(38, 28) <= 0; cloud_xl(38, 29) <= 0; cloud_xl(38, 30) <= 0; cloud_xl(38, 31) <= 0; cloud_xl(38, 32) <= 0; cloud_xl(38, 33) <= 0; cloud_xl(38, 34) <= 0; cloud_xl(38, 35) <= 0; cloud_xl(38, 36) <= 0; cloud_xl(38, 37) <= 0; cloud_xl(38, 38) <= 0; cloud_xl(38, 39) <= 0; cloud_xl(38, 40) <= 0; cloud_xl(38, 41) <= 0; cloud_xl(38, 42) <= 0; cloud_xl(38, 43) <= 0; cloud_xl(38, 44) <= 0; cloud_xl(38, 45) <= 0; cloud_xl(38, 46) <= 0; cloud_xl(38, 47) <= 0; cloud_xl(38, 48) <= 0; cloud_xl(38, 49) <= 0; cloud_xl(38, 50) <= 0; cloud_xl(38, 51) <= 0; cloud_xl(38, 52) <= 0; cloud_xl(38, 53) <= 0; cloud_xl(38, 54) <= 0; cloud_xl(38, 55) <= 0; cloud_xl(38, 56) <= 0; cloud_xl(38, 57) <= 0; cloud_xl(38, 58) <= 0; cloud_xl(38, 59) <= 0; cloud_xl(38, 60) <= 0; cloud_xl(38, 61) <= 0; cloud_xl(38, 62) <= 0; cloud_xl(38, 63) <= 0; cloud_xl(38, 64) <= 0; cloud_xl(38, 65) <= 0; cloud_xl(38, 66) <= 0; cloud_xl(38, 67) <= 0; cloud_xl(38, 68) <= 0; cloud_xl(38, 69) <= 0; cloud_xl(38, 70) <= 0; cloud_xl(38, 71) <= 0; cloud_xl(38, 72) <= 1; cloud_xl(38, 73) <= 1; cloud_xl(38, 74) <= 1; cloud_xl(38, 75) <= 1; cloud_xl(38, 76) <= 1; cloud_xl(38, 77) <= 1; 
cloud_xl(39, 0) <= 1; cloud_xl(39, 1) <= 1; cloud_xl(39, 2) <= 1; cloud_xl(39, 3) <= 1; cloud_xl(39, 4) <= 1; cloud_xl(39, 5) <= 1; cloud_xl(39, 6) <= 0; cloud_xl(39, 7) <= 0; cloud_xl(39, 8) <= 0; cloud_xl(39, 9) <= 0; cloud_xl(39, 10) <= 0; cloud_xl(39, 11) <= 0; cloud_xl(39, 12) <= 0; cloud_xl(39, 13) <= 0; cloud_xl(39, 14) <= 0; cloud_xl(39, 15) <= 0; cloud_xl(39, 16) <= 0; cloud_xl(39, 17) <= 0; cloud_xl(39, 18) <= 0; cloud_xl(39, 19) <= 0; cloud_xl(39, 20) <= 0; cloud_xl(39, 21) <= 0; cloud_xl(39, 22) <= 0; cloud_xl(39, 23) <= 0; cloud_xl(39, 24) <= 0; cloud_xl(39, 25) <= 0; cloud_xl(39, 26) <= 0; cloud_xl(39, 27) <= 0; cloud_xl(39, 28) <= 0; cloud_xl(39, 29) <= 0; cloud_xl(39, 30) <= 0; cloud_xl(39, 31) <= 0; cloud_xl(39, 32) <= 0; cloud_xl(39, 33) <= 0; cloud_xl(39, 34) <= 0; cloud_xl(39, 35) <= 0; cloud_xl(39, 36) <= 0; cloud_xl(39, 37) <= 0; cloud_xl(39, 38) <= 0; cloud_xl(39, 39) <= 0; cloud_xl(39, 40) <= 0; cloud_xl(39, 41) <= 0; cloud_xl(39, 42) <= 0; cloud_xl(39, 43) <= 0; cloud_xl(39, 44) <= 0; cloud_xl(39, 45) <= 0; cloud_xl(39, 46) <= 0; cloud_xl(39, 47) <= 0; cloud_xl(39, 48) <= 0; cloud_xl(39, 49) <= 0; cloud_xl(39, 50) <= 0; cloud_xl(39, 51) <= 0; cloud_xl(39, 52) <= 0; cloud_xl(39, 53) <= 0; cloud_xl(39, 54) <= 0; cloud_xl(39, 55) <= 0; cloud_xl(39, 56) <= 0; cloud_xl(39, 57) <= 0; cloud_xl(39, 58) <= 0; cloud_xl(39, 59) <= 0; cloud_xl(39, 60) <= 0; cloud_xl(39, 61) <= 0; cloud_xl(39, 62) <= 0; cloud_xl(39, 63) <= 0; cloud_xl(39, 64) <= 0; cloud_xl(39, 65) <= 0; cloud_xl(39, 66) <= 0; cloud_xl(39, 67) <= 0; cloud_xl(39, 68) <= 0; cloud_xl(39, 69) <= 0; cloud_xl(39, 70) <= 0; cloud_xl(39, 71) <= 0; cloud_xl(39, 72) <= 1; cloud_xl(39, 73) <= 1; cloud_xl(39, 74) <= 1; cloud_xl(39, 75) <= 1; cloud_xl(39, 76) <= 1; cloud_xl(39, 77) <= 1; 
cloud_xl(40, 0) <= 1; cloud_xl(40, 1) <= 1; cloud_xl(40, 2) <= 1; cloud_xl(40, 3) <= 1; cloud_xl(40, 4) <= 1; cloud_xl(40, 5) <= 1; cloud_xl(40, 6) <= 0; cloud_xl(40, 7) <= 0; cloud_xl(40, 8) <= 0; cloud_xl(40, 9) <= 0; cloud_xl(40, 10) <= 0; cloud_xl(40, 11) <= 0; cloud_xl(40, 12) <= 0; cloud_xl(40, 13) <= 0; cloud_xl(40, 14) <= 0; cloud_xl(40, 15) <= 0; cloud_xl(40, 16) <= 0; cloud_xl(40, 17) <= 0; cloud_xl(40, 18) <= 0; cloud_xl(40, 19) <= 0; cloud_xl(40, 20) <= 0; cloud_xl(40, 21) <= 0; cloud_xl(40, 22) <= 0; cloud_xl(40, 23) <= 0; cloud_xl(40, 24) <= 0; cloud_xl(40, 25) <= 0; cloud_xl(40, 26) <= 0; cloud_xl(40, 27) <= 0; cloud_xl(40, 28) <= 0; cloud_xl(40, 29) <= 0; cloud_xl(40, 30) <= 0; cloud_xl(40, 31) <= 0; cloud_xl(40, 32) <= 0; cloud_xl(40, 33) <= 0; cloud_xl(40, 34) <= 0; cloud_xl(40, 35) <= 0; cloud_xl(40, 36) <= 0; cloud_xl(40, 37) <= 0; cloud_xl(40, 38) <= 0; cloud_xl(40, 39) <= 0; cloud_xl(40, 40) <= 0; cloud_xl(40, 41) <= 0; cloud_xl(40, 42) <= 0; cloud_xl(40, 43) <= 0; cloud_xl(40, 44) <= 0; cloud_xl(40, 45) <= 0; cloud_xl(40, 46) <= 0; cloud_xl(40, 47) <= 0; cloud_xl(40, 48) <= 0; cloud_xl(40, 49) <= 0; cloud_xl(40, 50) <= 0; cloud_xl(40, 51) <= 0; cloud_xl(40, 52) <= 0; cloud_xl(40, 53) <= 0; cloud_xl(40, 54) <= 0; cloud_xl(40, 55) <= 0; cloud_xl(40, 56) <= 0; cloud_xl(40, 57) <= 0; cloud_xl(40, 58) <= 0; cloud_xl(40, 59) <= 0; cloud_xl(40, 60) <= 0; cloud_xl(40, 61) <= 0; cloud_xl(40, 62) <= 0; cloud_xl(40, 63) <= 0; cloud_xl(40, 64) <= 0; cloud_xl(40, 65) <= 0; cloud_xl(40, 66) <= 0; cloud_xl(40, 67) <= 0; cloud_xl(40, 68) <= 0; cloud_xl(40, 69) <= 0; cloud_xl(40, 70) <= 0; cloud_xl(40, 71) <= 0; cloud_xl(40, 72) <= 1; cloud_xl(40, 73) <= 1; cloud_xl(40, 74) <= 1; cloud_xl(40, 75) <= 1; cloud_xl(40, 76) <= 1; cloud_xl(40, 77) <= 1; 
cloud_xl(41, 0) <= 1; cloud_xl(41, 1) <= 1; cloud_xl(41, 2) <= 1; cloud_xl(41, 3) <= 1; cloud_xl(41, 4) <= 1; cloud_xl(41, 5) <= 1; cloud_xl(41, 6) <= 0; cloud_xl(41, 7) <= 0; cloud_xl(41, 8) <= 0; cloud_xl(41, 9) <= 0; cloud_xl(41, 10) <= 0; cloud_xl(41, 11) <= 0; cloud_xl(41, 12) <= 0; cloud_xl(41, 13) <= 0; cloud_xl(41, 14) <= 0; cloud_xl(41, 15) <= 0; cloud_xl(41, 16) <= 0; cloud_xl(41, 17) <= 0; cloud_xl(41, 18) <= 0; cloud_xl(41, 19) <= 0; cloud_xl(41, 20) <= 0; cloud_xl(41, 21) <= 0; cloud_xl(41, 22) <= 0; cloud_xl(41, 23) <= 0; cloud_xl(41, 24) <= 0; cloud_xl(41, 25) <= 0; cloud_xl(41, 26) <= 0; cloud_xl(41, 27) <= 0; cloud_xl(41, 28) <= 0; cloud_xl(41, 29) <= 0; cloud_xl(41, 30) <= 0; cloud_xl(41, 31) <= 0; cloud_xl(41, 32) <= 0; cloud_xl(41, 33) <= 0; cloud_xl(41, 34) <= 0; cloud_xl(41, 35) <= 0; cloud_xl(41, 36) <= 0; cloud_xl(41, 37) <= 0; cloud_xl(41, 38) <= 0; cloud_xl(41, 39) <= 0; cloud_xl(41, 40) <= 0; cloud_xl(41, 41) <= 0; cloud_xl(41, 42) <= 0; cloud_xl(41, 43) <= 0; cloud_xl(41, 44) <= 0; cloud_xl(41, 45) <= 0; cloud_xl(41, 46) <= 0; cloud_xl(41, 47) <= 0; cloud_xl(41, 48) <= 0; cloud_xl(41, 49) <= 0; cloud_xl(41, 50) <= 0; cloud_xl(41, 51) <= 0; cloud_xl(41, 52) <= 0; cloud_xl(41, 53) <= 0; cloud_xl(41, 54) <= 0; cloud_xl(41, 55) <= 0; cloud_xl(41, 56) <= 0; cloud_xl(41, 57) <= 0; cloud_xl(41, 58) <= 0; cloud_xl(41, 59) <= 0; cloud_xl(41, 60) <= 0; cloud_xl(41, 61) <= 0; cloud_xl(41, 62) <= 0; cloud_xl(41, 63) <= 0; cloud_xl(41, 64) <= 0; cloud_xl(41, 65) <= 0; cloud_xl(41, 66) <= 0; cloud_xl(41, 67) <= 0; cloud_xl(41, 68) <= 0; cloud_xl(41, 69) <= 0; cloud_xl(41, 70) <= 0; cloud_xl(41, 71) <= 0; cloud_xl(41, 72) <= 1; cloud_xl(41, 73) <= 1; cloud_xl(41, 74) <= 1; cloud_xl(41, 75) <= 1; cloud_xl(41, 76) <= 1; cloud_xl(41, 77) <= 1; 
cloud_xl(42, 0) <= 2; cloud_xl(42, 1) <= 2; cloud_xl(42, 2) <= 2; cloud_xl(42, 3) <= 2; cloud_xl(42, 4) <= 2; cloud_xl(42, 5) <= 2; cloud_xl(42, 6) <= 1; cloud_xl(42, 7) <= 1; cloud_xl(42, 8) <= 1; cloud_xl(42, 9) <= 1; cloud_xl(42, 10) <= 1; cloud_xl(42, 11) <= 1; cloud_xl(42, 12) <= 0; cloud_xl(42, 13) <= 0; cloud_xl(42, 14) <= 0; cloud_xl(42, 15) <= 0; cloud_xl(42, 16) <= 0; cloud_xl(42, 17) <= 0; cloud_xl(42, 18) <= 0; cloud_xl(42, 19) <= 0; cloud_xl(42, 20) <= 0; cloud_xl(42, 21) <= 0; cloud_xl(42, 22) <= 0; cloud_xl(42, 23) <= 0; cloud_xl(42, 24) <= 0; cloud_xl(42, 25) <= 0; cloud_xl(42, 26) <= 0; cloud_xl(42, 27) <= 0; cloud_xl(42, 28) <= 0; cloud_xl(42, 29) <= 0; cloud_xl(42, 30) <= 0; cloud_xl(42, 31) <= 0; cloud_xl(42, 32) <= 0; cloud_xl(42, 33) <= 0; cloud_xl(42, 34) <= 0; cloud_xl(42, 35) <= 0; cloud_xl(42, 36) <= 0; cloud_xl(42, 37) <= 0; cloud_xl(42, 38) <= 0; cloud_xl(42, 39) <= 0; cloud_xl(42, 40) <= 0; cloud_xl(42, 41) <= 0; cloud_xl(42, 42) <= 0; cloud_xl(42, 43) <= 0; cloud_xl(42, 44) <= 0; cloud_xl(42, 45) <= 0; cloud_xl(42, 46) <= 0; cloud_xl(42, 47) <= 0; cloud_xl(42, 48) <= 0; cloud_xl(42, 49) <= 0; cloud_xl(42, 50) <= 0; cloud_xl(42, 51) <= 0; cloud_xl(42, 52) <= 0; cloud_xl(42, 53) <= 0; cloud_xl(42, 54) <= 0; cloud_xl(42, 55) <= 0; cloud_xl(42, 56) <= 0; cloud_xl(42, 57) <= 0; cloud_xl(42, 58) <= 0; cloud_xl(42, 59) <= 0; cloud_xl(42, 60) <= 0; cloud_xl(42, 61) <= 0; cloud_xl(42, 62) <= 0; cloud_xl(42, 63) <= 0; cloud_xl(42, 64) <= 0; cloud_xl(42, 65) <= 0; cloud_xl(42, 66) <= 1; cloud_xl(42, 67) <= 1; cloud_xl(42, 68) <= 1; cloud_xl(42, 69) <= 1; cloud_xl(42, 70) <= 1; cloud_xl(42, 71) <= 1; cloud_xl(42, 72) <= 2; cloud_xl(42, 73) <= 2; cloud_xl(42, 74) <= 2; cloud_xl(42, 75) <= 2; cloud_xl(42, 76) <= 2; cloud_xl(42, 77) <= 2; 
cloud_xl(43, 0) <= 2; cloud_xl(43, 1) <= 2; cloud_xl(43, 2) <= 2; cloud_xl(43, 3) <= 2; cloud_xl(43, 4) <= 2; cloud_xl(43, 5) <= 2; cloud_xl(43, 6) <= 1; cloud_xl(43, 7) <= 1; cloud_xl(43, 8) <= 1; cloud_xl(43, 9) <= 1; cloud_xl(43, 10) <= 1; cloud_xl(43, 11) <= 1; cloud_xl(43, 12) <= 0; cloud_xl(43, 13) <= 0; cloud_xl(43, 14) <= 0; cloud_xl(43, 15) <= 0; cloud_xl(43, 16) <= 0; cloud_xl(43, 17) <= 0; cloud_xl(43, 18) <= 0; cloud_xl(43, 19) <= 0; cloud_xl(43, 20) <= 0; cloud_xl(43, 21) <= 0; cloud_xl(43, 22) <= 0; cloud_xl(43, 23) <= 0; cloud_xl(43, 24) <= 0; cloud_xl(43, 25) <= 0; cloud_xl(43, 26) <= 0; cloud_xl(43, 27) <= 0; cloud_xl(43, 28) <= 0; cloud_xl(43, 29) <= 0; cloud_xl(43, 30) <= 0; cloud_xl(43, 31) <= 0; cloud_xl(43, 32) <= 0; cloud_xl(43, 33) <= 0; cloud_xl(43, 34) <= 0; cloud_xl(43, 35) <= 0; cloud_xl(43, 36) <= 0; cloud_xl(43, 37) <= 0; cloud_xl(43, 38) <= 0; cloud_xl(43, 39) <= 0; cloud_xl(43, 40) <= 0; cloud_xl(43, 41) <= 0; cloud_xl(43, 42) <= 0; cloud_xl(43, 43) <= 0; cloud_xl(43, 44) <= 0; cloud_xl(43, 45) <= 0; cloud_xl(43, 46) <= 0; cloud_xl(43, 47) <= 0; cloud_xl(43, 48) <= 0; cloud_xl(43, 49) <= 0; cloud_xl(43, 50) <= 0; cloud_xl(43, 51) <= 0; cloud_xl(43, 52) <= 0; cloud_xl(43, 53) <= 0; cloud_xl(43, 54) <= 0; cloud_xl(43, 55) <= 0; cloud_xl(43, 56) <= 0; cloud_xl(43, 57) <= 0; cloud_xl(43, 58) <= 0; cloud_xl(43, 59) <= 0; cloud_xl(43, 60) <= 0; cloud_xl(43, 61) <= 0; cloud_xl(43, 62) <= 0; cloud_xl(43, 63) <= 0; cloud_xl(43, 64) <= 0; cloud_xl(43, 65) <= 0; cloud_xl(43, 66) <= 1; cloud_xl(43, 67) <= 1; cloud_xl(43, 68) <= 1; cloud_xl(43, 69) <= 1; cloud_xl(43, 70) <= 1; cloud_xl(43, 71) <= 1; cloud_xl(43, 72) <= 2; cloud_xl(43, 73) <= 2; cloud_xl(43, 74) <= 2; cloud_xl(43, 75) <= 2; cloud_xl(43, 76) <= 2; cloud_xl(43, 77) <= 2; 
cloud_xl(44, 0) <= 2; cloud_xl(44, 1) <= 2; cloud_xl(44, 2) <= 2; cloud_xl(44, 3) <= 2; cloud_xl(44, 4) <= 2; cloud_xl(44, 5) <= 2; cloud_xl(44, 6) <= 1; cloud_xl(44, 7) <= 1; cloud_xl(44, 8) <= 1; cloud_xl(44, 9) <= 1; cloud_xl(44, 10) <= 1; cloud_xl(44, 11) <= 1; cloud_xl(44, 12) <= 0; cloud_xl(44, 13) <= 0; cloud_xl(44, 14) <= 0; cloud_xl(44, 15) <= 0; cloud_xl(44, 16) <= 0; cloud_xl(44, 17) <= 0; cloud_xl(44, 18) <= 0; cloud_xl(44, 19) <= 0; cloud_xl(44, 20) <= 0; cloud_xl(44, 21) <= 0; cloud_xl(44, 22) <= 0; cloud_xl(44, 23) <= 0; cloud_xl(44, 24) <= 0; cloud_xl(44, 25) <= 0; cloud_xl(44, 26) <= 0; cloud_xl(44, 27) <= 0; cloud_xl(44, 28) <= 0; cloud_xl(44, 29) <= 0; cloud_xl(44, 30) <= 0; cloud_xl(44, 31) <= 0; cloud_xl(44, 32) <= 0; cloud_xl(44, 33) <= 0; cloud_xl(44, 34) <= 0; cloud_xl(44, 35) <= 0; cloud_xl(44, 36) <= 0; cloud_xl(44, 37) <= 0; cloud_xl(44, 38) <= 0; cloud_xl(44, 39) <= 0; cloud_xl(44, 40) <= 0; cloud_xl(44, 41) <= 0; cloud_xl(44, 42) <= 0; cloud_xl(44, 43) <= 0; cloud_xl(44, 44) <= 0; cloud_xl(44, 45) <= 0; cloud_xl(44, 46) <= 0; cloud_xl(44, 47) <= 0; cloud_xl(44, 48) <= 0; cloud_xl(44, 49) <= 0; cloud_xl(44, 50) <= 0; cloud_xl(44, 51) <= 0; cloud_xl(44, 52) <= 0; cloud_xl(44, 53) <= 0; cloud_xl(44, 54) <= 0; cloud_xl(44, 55) <= 0; cloud_xl(44, 56) <= 0; cloud_xl(44, 57) <= 0; cloud_xl(44, 58) <= 0; cloud_xl(44, 59) <= 0; cloud_xl(44, 60) <= 0; cloud_xl(44, 61) <= 0; cloud_xl(44, 62) <= 0; cloud_xl(44, 63) <= 0; cloud_xl(44, 64) <= 0; cloud_xl(44, 65) <= 0; cloud_xl(44, 66) <= 1; cloud_xl(44, 67) <= 1; cloud_xl(44, 68) <= 1; cloud_xl(44, 69) <= 1; cloud_xl(44, 70) <= 1; cloud_xl(44, 71) <= 1; cloud_xl(44, 72) <= 2; cloud_xl(44, 73) <= 2; cloud_xl(44, 74) <= 2; cloud_xl(44, 75) <= 2; cloud_xl(44, 76) <= 2; cloud_xl(44, 77) <= 2; 
cloud_xl(45, 0) <= 2; cloud_xl(45, 1) <= 2; cloud_xl(45, 2) <= 2; cloud_xl(45, 3) <= 2; cloud_xl(45, 4) <= 2; cloud_xl(45, 5) <= 2; cloud_xl(45, 6) <= 1; cloud_xl(45, 7) <= 1; cloud_xl(45, 8) <= 1; cloud_xl(45, 9) <= 1; cloud_xl(45, 10) <= 1; cloud_xl(45, 11) <= 1; cloud_xl(45, 12) <= 0; cloud_xl(45, 13) <= 0; cloud_xl(45, 14) <= 0; cloud_xl(45, 15) <= 0; cloud_xl(45, 16) <= 0; cloud_xl(45, 17) <= 0; cloud_xl(45, 18) <= 0; cloud_xl(45, 19) <= 0; cloud_xl(45, 20) <= 0; cloud_xl(45, 21) <= 0; cloud_xl(45, 22) <= 0; cloud_xl(45, 23) <= 0; cloud_xl(45, 24) <= 0; cloud_xl(45, 25) <= 0; cloud_xl(45, 26) <= 0; cloud_xl(45, 27) <= 0; cloud_xl(45, 28) <= 0; cloud_xl(45, 29) <= 0; cloud_xl(45, 30) <= 0; cloud_xl(45, 31) <= 0; cloud_xl(45, 32) <= 0; cloud_xl(45, 33) <= 0; cloud_xl(45, 34) <= 0; cloud_xl(45, 35) <= 0; cloud_xl(45, 36) <= 0; cloud_xl(45, 37) <= 0; cloud_xl(45, 38) <= 0; cloud_xl(45, 39) <= 0; cloud_xl(45, 40) <= 0; cloud_xl(45, 41) <= 0; cloud_xl(45, 42) <= 0; cloud_xl(45, 43) <= 0; cloud_xl(45, 44) <= 0; cloud_xl(45, 45) <= 0; cloud_xl(45, 46) <= 0; cloud_xl(45, 47) <= 0; cloud_xl(45, 48) <= 0; cloud_xl(45, 49) <= 0; cloud_xl(45, 50) <= 0; cloud_xl(45, 51) <= 0; cloud_xl(45, 52) <= 0; cloud_xl(45, 53) <= 0; cloud_xl(45, 54) <= 0; cloud_xl(45, 55) <= 0; cloud_xl(45, 56) <= 0; cloud_xl(45, 57) <= 0; cloud_xl(45, 58) <= 0; cloud_xl(45, 59) <= 0; cloud_xl(45, 60) <= 0; cloud_xl(45, 61) <= 0; cloud_xl(45, 62) <= 0; cloud_xl(45, 63) <= 0; cloud_xl(45, 64) <= 0; cloud_xl(45, 65) <= 0; cloud_xl(45, 66) <= 1; cloud_xl(45, 67) <= 1; cloud_xl(45, 68) <= 1; cloud_xl(45, 69) <= 1; cloud_xl(45, 70) <= 1; cloud_xl(45, 71) <= 1; cloud_xl(45, 72) <= 2; cloud_xl(45, 73) <= 2; cloud_xl(45, 74) <= 2; cloud_xl(45, 75) <= 2; cloud_xl(45, 76) <= 2; cloud_xl(45, 77) <= 2; 
cloud_xl(46, 0) <= 2; cloud_xl(46, 1) <= 2; cloud_xl(46, 2) <= 2; cloud_xl(46, 3) <= 2; cloud_xl(46, 4) <= 2; cloud_xl(46, 5) <= 2; cloud_xl(46, 6) <= 1; cloud_xl(46, 7) <= 1; cloud_xl(46, 8) <= 1; cloud_xl(46, 9) <= 1; cloud_xl(46, 10) <= 1; cloud_xl(46, 11) <= 1; cloud_xl(46, 12) <= 0; cloud_xl(46, 13) <= 0; cloud_xl(46, 14) <= 0; cloud_xl(46, 15) <= 0; cloud_xl(46, 16) <= 0; cloud_xl(46, 17) <= 0; cloud_xl(46, 18) <= 0; cloud_xl(46, 19) <= 0; cloud_xl(46, 20) <= 0; cloud_xl(46, 21) <= 0; cloud_xl(46, 22) <= 0; cloud_xl(46, 23) <= 0; cloud_xl(46, 24) <= 0; cloud_xl(46, 25) <= 0; cloud_xl(46, 26) <= 0; cloud_xl(46, 27) <= 0; cloud_xl(46, 28) <= 0; cloud_xl(46, 29) <= 0; cloud_xl(46, 30) <= 0; cloud_xl(46, 31) <= 0; cloud_xl(46, 32) <= 0; cloud_xl(46, 33) <= 0; cloud_xl(46, 34) <= 0; cloud_xl(46, 35) <= 0; cloud_xl(46, 36) <= 0; cloud_xl(46, 37) <= 0; cloud_xl(46, 38) <= 0; cloud_xl(46, 39) <= 0; cloud_xl(46, 40) <= 0; cloud_xl(46, 41) <= 0; cloud_xl(46, 42) <= 0; cloud_xl(46, 43) <= 0; cloud_xl(46, 44) <= 0; cloud_xl(46, 45) <= 0; cloud_xl(46, 46) <= 0; cloud_xl(46, 47) <= 0; cloud_xl(46, 48) <= 0; cloud_xl(46, 49) <= 0; cloud_xl(46, 50) <= 0; cloud_xl(46, 51) <= 0; cloud_xl(46, 52) <= 0; cloud_xl(46, 53) <= 0; cloud_xl(46, 54) <= 0; cloud_xl(46, 55) <= 0; cloud_xl(46, 56) <= 0; cloud_xl(46, 57) <= 0; cloud_xl(46, 58) <= 0; cloud_xl(46, 59) <= 0; cloud_xl(46, 60) <= 0; cloud_xl(46, 61) <= 0; cloud_xl(46, 62) <= 0; cloud_xl(46, 63) <= 0; cloud_xl(46, 64) <= 0; cloud_xl(46, 65) <= 0; cloud_xl(46, 66) <= 1; cloud_xl(46, 67) <= 1; cloud_xl(46, 68) <= 1; cloud_xl(46, 69) <= 1; cloud_xl(46, 70) <= 1; cloud_xl(46, 71) <= 1; cloud_xl(46, 72) <= 2; cloud_xl(46, 73) <= 2; cloud_xl(46, 74) <= 2; cloud_xl(46, 75) <= 2; cloud_xl(46, 76) <= 2; cloud_xl(46, 77) <= 2; 
cloud_xl(47, 0) <= 2; cloud_xl(47, 1) <= 2; cloud_xl(47, 2) <= 2; cloud_xl(47, 3) <= 2; cloud_xl(47, 4) <= 2; cloud_xl(47, 5) <= 2; cloud_xl(47, 6) <= 1; cloud_xl(47, 7) <= 1; cloud_xl(47, 8) <= 1; cloud_xl(47, 9) <= 1; cloud_xl(47, 10) <= 1; cloud_xl(47, 11) <= 1; cloud_xl(47, 12) <= 0; cloud_xl(47, 13) <= 0; cloud_xl(47, 14) <= 0; cloud_xl(47, 15) <= 0; cloud_xl(47, 16) <= 0; cloud_xl(47, 17) <= 0; cloud_xl(47, 18) <= 0; cloud_xl(47, 19) <= 0; cloud_xl(47, 20) <= 0; cloud_xl(47, 21) <= 0; cloud_xl(47, 22) <= 0; cloud_xl(47, 23) <= 0; cloud_xl(47, 24) <= 0; cloud_xl(47, 25) <= 0; cloud_xl(47, 26) <= 0; cloud_xl(47, 27) <= 0; cloud_xl(47, 28) <= 0; cloud_xl(47, 29) <= 0; cloud_xl(47, 30) <= 0; cloud_xl(47, 31) <= 0; cloud_xl(47, 32) <= 0; cloud_xl(47, 33) <= 0; cloud_xl(47, 34) <= 0; cloud_xl(47, 35) <= 0; cloud_xl(47, 36) <= 0; cloud_xl(47, 37) <= 0; cloud_xl(47, 38) <= 0; cloud_xl(47, 39) <= 0; cloud_xl(47, 40) <= 0; cloud_xl(47, 41) <= 0; cloud_xl(47, 42) <= 0; cloud_xl(47, 43) <= 0; cloud_xl(47, 44) <= 0; cloud_xl(47, 45) <= 0; cloud_xl(47, 46) <= 0; cloud_xl(47, 47) <= 0; cloud_xl(47, 48) <= 0; cloud_xl(47, 49) <= 0; cloud_xl(47, 50) <= 0; cloud_xl(47, 51) <= 0; cloud_xl(47, 52) <= 0; cloud_xl(47, 53) <= 0; cloud_xl(47, 54) <= 0; cloud_xl(47, 55) <= 0; cloud_xl(47, 56) <= 0; cloud_xl(47, 57) <= 0; cloud_xl(47, 58) <= 0; cloud_xl(47, 59) <= 0; cloud_xl(47, 60) <= 0; cloud_xl(47, 61) <= 0; cloud_xl(47, 62) <= 0; cloud_xl(47, 63) <= 0; cloud_xl(47, 64) <= 0; cloud_xl(47, 65) <= 0; cloud_xl(47, 66) <= 1; cloud_xl(47, 67) <= 1; cloud_xl(47, 68) <= 1; cloud_xl(47, 69) <= 1; cloud_xl(47, 70) <= 1; cloud_xl(47, 71) <= 1; cloud_xl(47, 72) <= 2; cloud_xl(47, 73) <= 2; cloud_xl(47, 74) <= 2; cloud_xl(47, 75) <= 2; cloud_xl(47, 76) <= 2; cloud_xl(47, 77) <= 2; 
cloud_xl(48, 0) <= 2; cloud_xl(48, 1) <= 2; cloud_xl(48, 2) <= 2; cloud_xl(48, 3) <= 2; cloud_xl(48, 4) <= 2; cloud_xl(48, 5) <= 2; cloud_xl(48, 6) <= 2; cloud_xl(48, 7) <= 2; cloud_xl(48, 8) <= 2; cloud_xl(48, 9) <= 2; cloud_xl(48, 10) <= 2; cloud_xl(48, 11) <= 2; cloud_xl(48, 12) <= 1; cloud_xl(48, 13) <= 1; cloud_xl(48, 14) <= 1; cloud_xl(48, 15) <= 1; cloud_xl(48, 16) <= 1; cloud_xl(48, 17) <= 1; cloud_xl(48, 18) <= 1; cloud_xl(48, 19) <= 1; cloud_xl(48, 20) <= 1; cloud_xl(48, 21) <= 1; cloud_xl(48, 22) <= 1; cloud_xl(48, 23) <= 1; cloud_xl(48, 24) <= 1; cloud_xl(48, 25) <= 1; cloud_xl(48, 26) <= 1; cloud_xl(48, 27) <= 1; cloud_xl(48, 28) <= 1; cloud_xl(48, 29) <= 1; cloud_xl(48, 30) <= 1; cloud_xl(48, 31) <= 1; cloud_xl(48, 32) <= 1; cloud_xl(48, 33) <= 1; cloud_xl(48, 34) <= 1; cloud_xl(48, 35) <= 1; cloud_xl(48, 36) <= 1; cloud_xl(48, 37) <= 1; cloud_xl(48, 38) <= 1; cloud_xl(48, 39) <= 1; cloud_xl(48, 40) <= 1; cloud_xl(48, 41) <= 1; cloud_xl(48, 42) <= 1; cloud_xl(48, 43) <= 1; cloud_xl(48, 44) <= 1; cloud_xl(48, 45) <= 1; cloud_xl(48, 46) <= 1; cloud_xl(48, 47) <= 1; cloud_xl(48, 48) <= 1; cloud_xl(48, 49) <= 1; cloud_xl(48, 50) <= 1; cloud_xl(48, 51) <= 1; cloud_xl(48, 52) <= 1; cloud_xl(48, 53) <= 1; cloud_xl(48, 54) <= 1; cloud_xl(48, 55) <= 1; cloud_xl(48, 56) <= 1; cloud_xl(48, 57) <= 1; cloud_xl(48, 58) <= 1; cloud_xl(48, 59) <= 1; cloud_xl(48, 60) <= 1; cloud_xl(48, 61) <= 1; cloud_xl(48, 62) <= 1; cloud_xl(48, 63) <= 1; cloud_xl(48, 64) <= 1; cloud_xl(48, 65) <= 1; cloud_xl(48, 66) <= 2; cloud_xl(48, 67) <= 2; cloud_xl(48, 68) <= 2; cloud_xl(48, 69) <= 2; cloud_xl(48, 70) <= 2; cloud_xl(48, 71) <= 2; cloud_xl(48, 72) <= 2; cloud_xl(48, 73) <= 2; cloud_xl(48, 74) <= 2; cloud_xl(48, 75) <= 2; cloud_xl(48, 76) <= 2; cloud_xl(48, 77) <= 2; 
cloud_xl(49, 0) <= 2; cloud_xl(49, 1) <= 2; cloud_xl(49, 2) <= 2; cloud_xl(49, 3) <= 2; cloud_xl(49, 4) <= 2; cloud_xl(49, 5) <= 2; cloud_xl(49, 6) <= 2; cloud_xl(49, 7) <= 2; cloud_xl(49, 8) <= 2; cloud_xl(49, 9) <= 2; cloud_xl(49, 10) <= 2; cloud_xl(49, 11) <= 2; cloud_xl(49, 12) <= 1; cloud_xl(49, 13) <= 1; cloud_xl(49, 14) <= 1; cloud_xl(49, 15) <= 1; cloud_xl(49, 16) <= 1; cloud_xl(49, 17) <= 1; cloud_xl(49, 18) <= 1; cloud_xl(49, 19) <= 1; cloud_xl(49, 20) <= 1; cloud_xl(49, 21) <= 1; cloud_xl(49, 22) <= 1; cloud_xl(49, 23) <= 1; cloud_xl(49, 24) <= 1; cloud_xl(49, 25) <= 1; cloud_xl(49, 26) <= 1; cloud_xl(49, 27) <= 1; cloud_xl(49, 28) <= 1; cloud_xl(49, 29) <= 1; cloud_xl(49, 30) <= 1; cloud_xl(49, 31) <= 1; cloud_xl(49, 32) <= 1; cloud_xl(49, 33) <= 1; cloud_xl(49, 34) <= 1; cloud_xl(49, 35) <= 1; cloud_xl(49, 36) <= 1; cloud_xl(49, 37) <= 1; cloud_xl(49, 38) <= 1; cloud_xl(49, 39) <= 1; cloud_xl(49, 40) <= 1; cloud_xl(49, 41) <= 1; cloud_xl(49, 42) <= 1; cloud_xl(49, 43) <= 1; cloud_xl(49, 44) <= 1; cloud_xl(49, 45) <= 1; cloud_xl(49, 46) <= 1; cloud_xl(49, 47) <= 1; cloud_xl(49, 48) <= 1; cloud_xl(49, 49) <= 1; cloud_xl(49, 50) <= 1; cloud_xl(49, 51) <= 1; cloud_xl(49, 52) <= 1; cloud_xl(49, 53) <= 1; cloud_xl(49, 54) <= 1; cloud_xl(49, 55) <= 1; cloud_xl(49, 56) <= 1; cloud_xl(49, 57) <= 1; cloud_xl(49, 58) <= 1; cloud_xl(49, 59) <= 1; cloud_xl(49, 60) <= 1; cloud_xl(49, 61) <= 1; cloud_xl(49, 62) <= 1; cloud_xl(49, 63) <= 1; cloud_xl(49, 64) <= 1; cloud_xl(49, 65) <= 1; cloud_xl(49, 66) <= 2; cloud_xl(49, 67) <= 2; cloud_xl(49, 68) <= 2; cloud_xl(49, 69) <= 2; cloud_xl(49, 70) <= 2; cloud_xl(49, 71) <= 2; cloud_xl(49, 72) <= 2; cloud_xl(49, 73) <= 2; cloud_xl(49, 74) <= 2; cloud_xl(49, 75) <= 2; cloud_xl(49, 76) <= 2; cloud_xl(49, 77) <= 2; 
cloud_xl(50, 0) <= 2; cloud_xl(50, 1) <= 2; cloud_xl(50, 2) <= 2; cloud_xl(50, 3) <= 2; cloud_xl(50, 4) <= 2; cloud_xl(50, 5) <= 2; cloud_xl(50, 6) <= 2; cloud_xl(50, 7) <= 2; cloud_xl(50, 8) <= 2; cloud_xl(50, 9) <= 2; cloud_xl(50, 10) <= 2; cloud_xl(50, 11) <= 2; cloud_xl(50, 12) <= 1; cloud_xl(50, 13) <= 1; cloud_xl(50, 14) <= 1; cloud_xl(50, 15) <= 1; cloud_xl(50, 16) <= 1; cloud_xl(50, 17) <= 1; cloud_xl(50, 18) <= 1; cloud_xl(50, 19) <= 1; cloud_xl(50, 20) <= 1; cloud_xl(50, 21) <= 1; cloud_xl(50, 22) <= 1; cloud_xl(50, 23) <= 1; cloud_xl(50, 24) <= 1; cloud_xl(50, 25) <= 1; cloud_xl(50, 26) <= 1; cloud_xl(50, 27) <= 1; cloud_xl(50, 28) <= 1; cloud_xl(50, 29) <= 1; cloud_xl(50, 30) <= 1; cloud_xl(50, 31) <= 1; cloud_xl(50, 32) <= 1; cloud_xl(50, 33) <= 1; cloud_xl(50, 34) <= 1; cloud_xl(50, 35) <= 1; cloud_xl(50, 36) <= 1; cloud_xl(50, 37) <= 1; cloud_xl(50, 38) <= 1; cloud_xl(50, 39) <= 1; cloud_xl(50, 40) <= 1; cloud_xl(50, 41) <= 1; cloud_xl(50, 42) <= 1; cloud_xl(50, 43) <= 1; cloud_xl(50, 44) <= 1; cloud_xl(50, 45) <= 1; cloud_xl(50, 46) <= 1; cloud_xl(50, 47) <= 1; cloud_xl(50, 48) <= 1; cloud_xl(50, 49) <= 1; cloud_xl(50, 50) <= 1; cloud_xl(50, 51) <= 1; cloud_xl(50, 52) <= 1; cloud_xl(50, 53) <= 1; cloud_xl(50, 54) <= 1; cloud_xl(50, 55) <= 1; cloud_xl(50, 56) <= 1; cloud_xl(50, 57) <= 1; cloud_xl(50, 58) <= 1; cloud_xl(50, 59) <= 1; cloud_xl(50, 60) <= 1; cloud_xl(50, 61) <= 1; cloud_xl(50, 62) <= 1; cloud_xl(50, 63) <= 1; cloud_xl(50, 64) <= 1; cloud_xl(50, 65) <= 1; cloud_xl(50, 66) <= 2; cloud_xl(50, 67) <= 2; cloud_xl(50, 68) <= 2; cloud_xl(50, 69) <= 2; cloud_xl(50, 70) <= 2; cloud_xl(50, 71) <= 2; cloud_xl(50, 72) <= 2; cloud_xl(50, 73) <= 2; cloud_xl(50, 74) <= 2; cloud_xl(50, 75) <= 2; cloud_xl(50, 76) <= 2; cloud_xl(50, 77) <= 2; 
cloud_xl(51, 0) <= 2; cloud_xl(51, 1) <= 2; cloud_xl(51, 2) <= 2; cloud_xl(51, 3) <= 2; cloud_xl(51, 4) <= 2; cloud_xl(51, 5) <= 2; cloud_xl(51, 6) <= 2; cloud_xl(51, 7) <= 2; cloud_xl(51, 8) <= 2; cloud_xl(51, 9) <= 2; cloud_xl(51, 10) <= 2; cloud_xl(51, 11) <= 2; cloud_xl(51, 12) <= 1; cloud_xl(51, 13) <= 1; cloud_xl(51, 14) <= 1; cloud_xl(51, 15) <= 1; cloud_xl(51, 16) <= 1; cloud_xl(51, 17) <= 1; cloud_xl(51, 18) <= 1; cloud_xl(51, 19) <= 1; cloud_xl(51, 20) <= 1; cloud_xl(51, 21) <= 1; cloud_xl(51, 22) <= 1; cloud_xl(51, 23) <= 1; cloud_xl(51, 24) <= 1; cloud_xl(51, 25) <= 1; cloud_xl(51, 26) <= 1; cloud_xl(51, 27) <= 1; cloud_xl(51, 28) <= 1; cloud_xl(51, 29) <= 1; cloud_xl(51, 30) <= 1; cloud_xl(51, 31) <= 1; cloud_xl(51, 32) <= 1; cloud_xl(51, 33) <= 1; cloud_xl(51, 34) <= 1; cloud_xl(51, 35) <= 1; cloud_xl(51, 36) <= 1; cloud_xl(51, 37) <= 1; cloud_xl(51, 38) <= 1; cloud_xl(51, 39) <= 1; cloud_xl(51, 40) <= 1; cloud_xl(51, 41) <= 1; cloud_xl(51, 42) <= 1; cloud_xl(51, 43) <= 1; cloud_xl(51, 44) <= 1; cloud_xl(51, 45) <= 1; cloud_xl(51, 46) <= 1; cloud_xl(51, 47) <= 1; cloud_xl(51, 48) <= 1; cloud_xl(51, 49) <= 1; cloud_xl(51, 50) <= 1; cloud_xl(51, 51) <= 1; cloud_xl(51, 52) <= 1; cloud_xl(51, 53) <= 1; cloud_xl(51, 54) <= 1; cloud_xl(51, 55) <= 1; cloud_xl(51, 56) <= 1; cloud_xl(51, 57) <= 1; cloud_xl(51, 58) <= 1; cloud_xl(51, 59) <= 1; cloud_xl(51, 60) <= 1; cloud_xl(51, 61) <= 1; cloud_xl(51, 62) <= 1; cloud_xl(51, 63) <= 1; cloud_xl(51, 64) <= 1; cloud_xl(51, 65) <= 1; cloud_xl(51, 66) <= 2; cloud_xl(51, 67) <= 2; cloud_xl(51, 68) <= 2; cloud_xl(51, 69) <= 2; cloud_xl(51, 70) <= 2; cloud_xl(51, 71) <= 2; cloud_xl(51, 72) <= 2; cloud_xl(51, 73) <= 2; cloud_xl(51, 74) <= 2; cloud_xl(51, 75) <= 2; cloud_xl(51, 76) <= 2; cloud_xl(51, 77) <= 2; 
cloud_xl(52, 0) <= 2; cloud_xl(52, 1) <= 2; cloud_xl(52, 2) <= 2; cloud_xl(52, 3) <= 2; cloud_xl(52, 4) <= 2; cloud_xl(52, 5) <= 2; cloud_xl(52, 6) <= 2; cloud_xl(52, 7) <= 2; cloud_xl(52, 8) <= 2; cloud_xl(52, 9) <= 2; cloud_xl(52, 10) <= 2; cloud_xl(52, 11) <= 2; cloud_xl(52, 12) <= 1; cloud_xl(52, 13) <= 1; cloud_xl(52, 14) <= 1; cloud_xl(52, 15) <= 1; cloud_xl(52, 16) <= 1; cloud_xl(52, 17) <= 1; cloud_xl(52, 18) <= 1; cloud_xl(52, 19) <= 1; cloud_xl(52, 20) <= 1; cloud_xl(52, 21) <= 1; cloud_xl(52, 22) <= 1; cloud_xl(52, 23) <= 1; cloud_xl(52, 24) <= 1; cloud_xl(52, 25) <= 1; cloud_xl(52, 26) <= 1; cloud_xl(52, 27) <= 1; cloud_xl(52, 28) <= 1; cloud_xl(52, 29) <= 1; cloud_xl(52, 30) <= 1; cloud_xl(52, 31) <= 1; cloud_xl(52, 32) <= 1; cloud_xl(52, 33) <= 1; cloud_xl(52, 34) <= 1; cloud_xl(52, 35) <= 1; cloud_xl(52, 36) <= 1; cloud_xl(52, 37) <= 1; cloud_xl(52, 38) <= 1; cloud_xl(52, 39) <= 1; cloud_xl(52, 40) <= 1; cloud_xl(52, 41) <= 1; cloud_xl(52, 42) <= 1; cloud_xl(52, 43) <= 1; cloud_xl(52, 44) <= 1; cloud_xl(52, 45) <= 1; cloud_xl(52, 46) <= 1; cloud_xl(52, 47) <= 1; cloud_xl(52, 48) <= 1; cloud_xl(52, 49) <= 1; cloud_xl(52, 50) <= 1; cloud_xl(52, 51) <= 1; cloud_xl(52, 52) <= 1; cloud_xl(52, 53) <= 1; cloud_xl(52, 54) <= 1; cloud_xl(52, 55) <= 1; cloud_xl(52, 56) <= 1; cloud_xl(52, 57) <= 1; cloud_xl(52, 58) <= 1; cloud_xl(52, 59) <= 1; cloud_xl(52, 60) <= 1; cloud_xl(52, 61) <= 1; cloud_xl(52, 62) <= 1; cloud_xl(52, 63) <= 1; cloud_xl(52, 64) <= 1; cloud_xl(52, 65) <= 1; cloud_xl(52, 66) <= 2; cloud_xl(52, 67) <= 2; cloud_xl(52, 68) <= 2; cloud_xl(52, 69) <= 2; cloud_xl(52, 70) <= 2; cloud_xl(52, 71) <= 2; cloud_xl(52, 72) <= 2; cloud_xl(52, 73) <= 2; cloud_xl(52, 74) <= 2; cloud_xl(52, 75) <= 2; cloud_xl(52, 76) <= 2; cloud_xl(52, 77) <= 2; 
cloud_xl(53, 0) <= 2; cloud_xl(53, 1) <= 2; cloud_xl(53, 2) <= 2; cloud_xl(53, 3) <= 2; cloud_xl(53, 4) <= 2; cloud_xl(53, 5) <= 2; cloud_xl(53, 6) <= 2; cloud_xl(53, 7) <= 2; cloud_xl(53, 8) <= 2; cloud_xl(53, 9) <= 2; cloud_xl(53, 10) <= 2; cloud_xl(53, 11) <= 2; cloud_xl(53, 12) <= 1; cloud_xl(53, 13) <= 1; cloud_xl(53, 14) <= 1; cloud_xl(53, 15) <= 1; cloud_xl(53, 16) <= 1; cloud_xl(53, 17) <= 1; cloud_xl(53, 18) <= 1; cloud_xl(53, 19) <= 1; cloud_xl(53, 20) <= 1; cloud_xl(53, 21) <= 1; cloud_xl(53, 22) <= 1; cloud_xl(53, 23) <= 1; cloud_xl(53, 24) <= 1; cloud_xl(53, 25) <= 1; cloud_xl(53, 26) <= 1; cloud_xl(53, 27) <= 1; cloud_xl(53, 28) <= 1; cloud_xl(53, 29) <= 1; cloud_xl(53, 30) <= 1; cloud_xl(53, 31) <= 1; cloud_xl(53, 32) <= 1; cloud_xl(53, 33) <= 1; cloud_xl(53, 34) <= 1; cloud_xl(53, 35) <= 1; cloud_xl(53, 36) <= 1; cloud_xl(53, 37) <= 1; cloud_xl(53, 38) <= 1; cloud_xl(53, 39) <= 1; cloud_xl(53, 40) <= 1; cloud_xl(53, 41) <= 1; cloud_xl(53, 42) <= 1; cloud_xl(53, 43) <= 1; cloud_xl(53, 44) <= 1; cloud_xl(53, 45) <= 1; cloud_xl(53, 46) <= 1; cloud_xl(53, 47) <= 1; cloud_xl(53, 48) <= 1; cloud_xl(53, 49) <= 1; cloud_xl(53, 50) <= 1; cloud_xl(53, 51) <= 1; cloud_xl(53, 52) <= 1; cloud_xl(53, 53) <= 1; cloud_xl(53, 54) <= 1; cloud_xl(53, 55) <= 1; cloud_xl(53, 56) <= 1; cloud_xl(53, 57) <= 1; cloud_xl(53, 58) <= 1; cloud_xl(53, 59) <= 1; cloud_xl(53, 60) <= 1; cloud_xl(53, 61) <= 1; cloud_xl(53, 62) <= 1; cloud_xl(53, 63) <= 1; cloud_xl(53, 64) <= 1; cloud_xl(53, 65) <= 1; cloud_xl(53, 66) <= 2; cloud_xl(53, 67) <= 2; cloud_xl(53, 68) <= 2; cloud_xl(53, 69) <= 2; cloud_xl(53, 70) <= 2; cloud_xl(53, 71) <= 2; cloud_xl(53, 72) <= 2; cloud_xl(53, 73) <= 2; cloud_xl(53, 74) <= 2; cloud_xl(53, 75) <= 2; cloud_xl(53, 76) <= 2; cloud_xl(53, 77) <= 2; 


end Behavioral;
