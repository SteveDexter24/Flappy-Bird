library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package vpkg is
    type largeAB is array(0 to 143, 0 to 149) of integer;
end package;

use work.vpkg.all;


entity largeAngryBird is
    Port (angryBirdLarge: out largeAB );
end largeAngryBird;

architecture Behavioral of largeAngryBird is

begin
angryBirdLarge(0, 0) <= 0; angryBirdLarge(0, 1) <= 0; angryBirdLarge(0, 2) <= 0; angryBirdLarge(0, 3) <= 0; angryBirdLarge(0, 4) <= 0; angryBirdLarge(0, 5) <= 0; angryBirdLarge(0, 6) <= 0; angryBirdLarge(0, 7) <= 0; angryBirdLarge(0, 8) <= 0; angryBirdLarge(0, 9) <= 0; angryBirdLarge(0, 10) <= 0; angryBirdLarge(0, 11) <= 0; angryBirdLarge(0, 12) <= 0; angryBirdLarge(0, 13) <= 0; angryBirdLarge(0, 14) <= 0; angryBirdLarge(0, 15) <= 0; angryBirdLarge(0, 16) <= 0; angryBirdLarge(0, 17) <= 0; angryBirdLarge(0, 18) <= 0; angryBirdLarge(0, 19) <= 0; angryBirdLarge(0, 20) <= 0; angryBirdLarge(0, 21) <= 0; angryBirdLarge(0, 22) <= 0; angryBirdLarge(0, 23) <= 0; angryBirdLarge(0, 24) <= 0; angryBirdLarge(0, 25) <= 0; angryBirdLarge(0, 26) <= 0; angryBirdLarge(0, 27) <= 0; angryBirdLarge(0, 28) <= 0; angryBirdLarge(0, 29) <= 0; angryBirdLarge(0, 30) <= 0; angryBirdLarge(0, 31) <= 0; angryBirdLarge(0, 32) <= 0; angryBirdLarge(0, 33) <= 0; angryBirdLarge(0, 34) <= 0; angryBirdLarge(0, 35) <= 0; angryBirdLarge(0, 36) <= 0; angryBirdLarge(0, 37) <= 0; angryBirdLarge(0, 38) <= 0; angryBirdLarge(0, 39) <= 0; angryBirdLarge(0, 40) <= 0; angryBirdLarge(0, 41) <= 0; angryBirdLarge(0, 42) <= 0; angryBirdLarge(0, 43) <= 0; angryBirdLarge(0, 44) <= 0; angryBirdLarge(0, 45) <= 0; angryBirdLarge(0, 46) <= 0; angryBirdLarge(0, 47) <= 0; angryBirdLarge(0, 48) <= 0; angryBirdLarge(0, 49) <= 0; angryBirdLarge(0, 50) <= 0; angryBirdLarge(0, 51) <= 0; angryBirdLarge(0, 52) <= 0; angryBirdLarge(0, 53) <= 0; angryBirdLarge(0, 54) <= 0; angryBirdLarge(0, 55) <= 0; angryBirdLarge(0, 56) <= 0; angryBirdLarge(0, 57) <= 0; angryBirdLarge(0, 58) <= 0; angryBirdLarge(0, 59) <= 0; angryBirdLarge(0, 60) <= 0; angryBirdLarge(0, 61) <= 0; angryBirdLarge(0, 62) <= 0; angryBirdLarge(0, 63) <= 0; angryBirdLarge(0, 64) <= 0; angryBirdLarge(0, 65) <= 0; angryBirdLarge(0, 66) <= 0; angryBirdLarge(0, 67) <= 0; angryBirdLarge(0, 68) <= 0; angryBirdLarge(0, 69) <= 0; angryBirdLarge(0, 70) <= 0; angryBirdLarge(0, 71) <= 0; angryBirdLarge(0, 72) <= 5; angryBirdLarge(0, 73) <= 5; angryBirdLarge(0, 74) <= 5; angryBirdLarge(0, 75) <= 5; angryBirdLarge(0, 76) <= 5; angryBirdLarge(0, 77) <= 5; angryBirdLarge(0, 78) <= 5; angryBirdLarge(0, 79) <= 5; angryBirdLarge(0, 80) <= 5; angryBirdLarge(0, 81) <= 5; angryBirdLarge(0, 82) <= 5; angryBirdLarge(0, 83) <= 5; angryBirdLarge(0, 84) <= 5; angryBirdLarge(0, 85) <= 5; angryBirdLarge(0, 86) <= 5; angryBirdLarge(0, 87) <= 5; angryBirdLarge(0, 88) <= 5; angryBirdLarge(0, 89) <= 5; angryBirdLarge(0, 90) <= 0; angryBirdLarge(0, 91) <= 0; angryBirdLarge(0, 92) <= 0; angryBirdLarge(0, 93) <= 0; angryBirdLarge(0, 94) <= 0; angryBirdLarge(0, 95) <= 0; angryBirdLarge(0, 96) <= 0; angryBirdLarge(0, 97) <= 0; angryBirdLarge(0, 98) <= 0; angryBirdLarge(0, 99) <= 0; angryBirdLarge(0, 100) <= 0; angryBirdLarge(0, 101) <= 0; angryBirdLarge(0, 102) <= 0; angryBirdLarge(0, 103) <= 0; angryBirdLarge(0, 104) <= 0; angryBirdLarge(0, 105) <= 0; angryBirdLarge(0, 106) <= 0; angryBirdLarge(0, 107) <= 0; angryBirdLarge(0, 108) <= 0; angryBirdLarge(0, 109) <= 0; angryBirdLarge(0, 110) <= 0; angryBirdLarge(0, 111) <= 0; angryBirdLarge(0, 112) <= 0; angryBirdLarge(0, 113) <= 0; angryBirdLarge(0, 114) <= 0; angryBirdLarge(0, 115) <= 0; angryBirdLarge(0, 116) <= 0; angryBirdLarge(0, 117) <= 0; angryBirdLarge(0, 118) <= 0; angryBirdLarge(0, 119) <= 0; angryBirdLarge(0, 120) <= 0; angryBirdLarge(0, 121) <= 0; angryBirdLarge(0, 122) <= 0; angryBirdLarge(0, 123) <= 0; angryBirdLarge(0, 124) <= 0; angryBirdLarge(0, 125) <= 0; angryBirdLarge(0, 126) <= 0; angryBirdLarge(0, 127) <= 0; angryBirdLarge(0, 128) <= 0; angryBirdLarge(0, 129) <= 0; angryBirdLarge(0, 130) <= 0; angryBirdLarge(0, 131) <= 0; angryBirdLarge(0, 132) <= 0; angryBirdLarge(0, 133) <= 0; angryBirdLarge(0, 134) <= 0; angryBirdLarge(0, 135) <= 0; angryBirdLarge(0, 136) <= 0; angryBirdLarge(0, 137) <= 0; angryBirdLarge(0, 138) <= 0; angryBirdLarge(0, 139) <= 0; angryBirdLarge(0, 140) <= 0; angryBirdLarge(0, 141) <= 0; angryBirdLarge(0, 142) <= 0; angryBirdLarge(0, 143) <= 0; angryBirdLarge(0, 144) <= 0; angryBirdLarge(0, 145) <= 0; angryBirdLarge(0, 146) <= 0; angryBirdLarge(0, 147) <= 0; angryBirdLarge(0, 148) <= 0; angryBirdLarge(0, 149) <= 0; 
angryBirdLarge(1, 0) <= 0; angryBirdLarge(1, 1) <= 0; angryBirdLarge(1, 2) <= 0; angryBirdLarge(1, 3) <= 0; angryBirdLarge(1, 4) <= 0; angryBirdLarge(1, 5) <= 0; angryBirdLarge(1, 6) <= 0; angryBirdLarge(1, 7) <= 0; angryBirdLarge(1, 8) <= 0; angryBirdLarge(1, 9) <= 0; angryBirdLarge(1, 10) <= 0; angryBirdLarge(1, 11) <= 0; angryBirdLarge(1, 12) <= 0; angryBirdLarge(1, 13) <= 0; angryBirdLarge(1, 14) <= 0; angryBirdLarge(1, 15) <= 0; angryBirdLarge(1, 16) <= 0; angryBirdLarge(1, 17) <= 0; angryBirdLarge(1, 18) <= 0; angryBirdLarge(1, 19) <= 0; angryBirdLarge(1, 20) <= 0; angryBirdLarge(1, 21) <= 0; angryBirdLarge(1, 22) <= 0; angryBirdLarge(1, 23) <= 0; angryBirdLarge(1, 24) <= 0; angryBirdLarge(1, 25) <= 0; angryBirdLarge(1, 26) <= 0; angryBirdLarge(1, 27) <= 0; angryBirdLarge(1, 28) <= 0; angryBirdLarge(1, 29) <= 0; angryBirdLarge(1, 30) <= 0; angryBirdLarge(1, 31) <= 0; angryBirdLarge(1, 32) <= 0; angryBirdLarge(1, 33) <= 0; angryBirdLarge(1, 34) <= 0; angryBirdLarge(1, 35) <= 0; angryBirdLarge(1, 36) <= 0; angryBirdLarge(1, 37) <= 0; angryBirdLarge(1, 38) <= 0; angryBirdLarge(1, 39) <= 0; angryBirdLarge(1, 40) <= 0; angryBirdLarge(1, 41) <= 0; angryBirdLarge(1, 42) <= 0; angryBirdLarge(1, 43) <= 0; angryBirdLarge(1, 44) <= 0; angryBirdLarge(1, 45) <= 0; angryBirdLarge(1, 46) <= 0; angryBirdLarge(1, 47) <= 0; angryBirdLarge(1, 48) <= 0; angryBirdLarge(1, 49) <= 0; angryBirdLarge(1, 50) <= 0; angryBirdLarge(1, 51) <= 0; angryBirdLarge(1, 52) <= 0; angryBirdLarge(1, 53) <= 0; angryBirdLarge(1, 54) <= 0; angryBirdLarge(1, 55) <= 0; angryBirdLarge(1, 56) <= 0; angryBirdLarge(1, 57) <= 0; angryBirdLarge(1, 58) <= 0; angryBirdLarge(1, 59) <= 0; angryBirdLarge(1, 60) <= 0; angryBirdLarge(1, 61) <= 0; angryBirdLarge(1, 62) <= 0; angryBirdLarge(1, 63) <= 0; angryBirdLarge(1, 64) <= 0; angryBirdLarge(1, 65) <= 0; angryBirdLarge(1, 66) <= 0; angryBirdLarge(1, 67) <= 0; angryBirdLarge(1, 68) <= 0; angryBirdLarge(1, 69) <= 0; angryBirdLarge(1, 70) <= 0; angryBirdLarge(1, 71) <= 0; angryBirdLarge(1, 72) <= 5; angryBirdLarge(1, 73) <= 5; angryBirdLarge(1, 74) <= 5; angryBirdLarge(1, 75) <= 5; angryBirdLarge(1, 76) <= 5; angryBirdLarge(1, 77) <= 5; angryBirdLarge(1, 78) <= 5; angryBirdLarge(1, 79) <= 5; angryBirdLarge(1, 80) <= 5; angryBirdLarge(1, 81) <= 5; angryBirdLarge(1, 82) <= 5; angryBirdLarge(1, 83) <= 5; angryBirdLarge(1, 84) <= 5; angryBirdLarge(1, 85) <= 5; angryBirdLarge(1, 86) <= 5; angryBirdLarge(1, 87) <= 5; angryBirdLarge(1, 88) <= 5; angryBirdLarge(1, 89) <= 5; angryBirdLarge(1, 90) <= 0; angryBirdLarge(1, 91) <= 0; angryBirdLarge(1, 92) <= 0; angryBirdLarge(1, 93) <= 0; angryBirdLarge(1, 94) <= 0; angryBirdLarge(1, 95) <= 0; angryBirdLarge(1, 96) <= 0; angryBirdLarge(1, 97) <= 0; angryBirdLarge(1, 98) <= 0; angryBirdLarge(1, 99) <= 0; angryBirdLarge(1, 100) <= 0; angryBirdLarge(1, 101) <= 0; angryBirdLarge(1, 102) <= 0; angryBirdLarge(1, 103) <= 0; angryBirdLarge(1, 104) <= 0; angryBirdLarge(1, 105) <= 0; angryBirdLarge(1, 106) <= 0; angryBirdLarge(1, 107) <= 0; angryBirdLarge(1, 108) <= 0; angryBirdLarge(1, 109) <= 0; angryBirdLarge(1, 110) <= 0; angryBirdLarge(1, 111) <= 0; angryBirdLarge(1, 112) <= 0; angryBirdLarge(1, 113) <= 0; angryBirdLarge(1, 114) <= 0; angryBirdLarge(1, 115) <= 0; angryBirdLarge(1, 116) <= 0; angryBirdLarge(1, 117) <= 0; angryBirdLarge(1, 118) <= 0; angryBirdLarge(1, 119) <= 0; angryBirdLarge(1, 120) <= 0; angryBirdLarge(1, 121) <= 0; angryBirdLarge(1, 122) <= 0; angryBirdLarge(1, 123) <= 0; angryBirdLarge(1, 124) <= 0; angryBirdLarge(1, 125) <= 0; angryBirdLarge(1, 126) <= 0; angryBirdLarge(1, 127) <= 0; angryBirdLarge(1, 128) <= 0; angryBirdLarge(1, 129) <= 0; angryBirdLarge(1, 130) <= 0; angryBirdLarge(1, 131) <= 0; angryBirdLarge(1, 132) <= 0; angryBirdLarge(1, 133) <= 0; angryBirdLarge(1, 134) <= 0; angryBirdLarge(1, 135) <= 0; angryBirdLarge(1, 136) <= 0; angryBirdLarge(1, 137) <= 0; angryBirdLarge(1, 138) <= 0; angryBirdLarge(1, 139) <= 0; angryBirdLarge(1, 140) <= 0; angryBirdLarge(1, 141) <= 0; angryBirdLarge(1, 142) <= 0; angryBirdLarge(1, 143) <= 0; angryBirdLarge(1, 144) <= 0; angryBirdLarge(1, 145) <= 0; angryBirdLarge(1, 146) <= 0; angryBirdLarge(1, 147) <= 0; angryBirdLarge(1, 148) <= 0; angryBirdLarge(1, 149) <= 0; 
angryBirdLarge(2, 0) <= 0; angryBirdLarge(2, 1) <= 0; angryBirdLarge(2, 2) <= 0; angryBirdLarge(2, 3) <= 0; angryBirdLarge(2, 4) <= 0; angryBirdLarge(2, 5) <= 0; angryBirdLarge(2, 6) <= 0; angryBirdLarge(2, 7) <= 0; angryBirdLarge(2, 8) <= 0; angryBirdLarge(2, 9) <= 0; angryBirdLarge(2, 10) <= 0; angryBirdLarge(2, 11) <= 0; angryBirdLarge(2, 12) <= 0; angryBirdLarge(2, 13) <= 0; angryBirdLarge(2, 14) <= 0; angryBirdLarge(2, 15) <= 0; angryBirdLarge(2, 16) <= 0; angryBirdLarge(2, 17) <= 0; angryBirdLarge(2, 18) <= 0; angryBirdLarge(2, 19) <= 0; angryBirdLarge(2, 20) <= 0; angryBirdLarge(2, 21) <= 0; angryBirdLarge(2, 22) <= 0; angryBirdLarge(2, 23) <= 0; angryBirdLarge(2, 24) <= 0; angryBirdLarge(2, 25) <= 0; angryBirdLarge(2, 26) <= 0; angryBirdLarge(2, 27) <= 0; angryBirdLarge(2, 28) <= 0; angryBirdLarge(2, 29) <= 0; angryBirdLarge(2, 30) <= 0; angryBirdLarge(2, 31) <= 0; angryBirdLarge(2, 32) <= 0; angryBirdLarge(2, 33) <= 0; angryBirdLarge(2, 34) <= 0; angryBirdLarge(2, 35) <= 0; angryBirdLarge(2, 36) <= 0; angryBirdLarge(2, 37) <= 0; angryBirdLarge(2, 38) <= 0; angryBirdLarge(2, 39) <= 0; angryBirdLarge(2, 40) <= 0; angryBirdLarge(2, 41) <= 0; angryBirdLarge(2, 42) <= 0; angryBirdLarge(2, 43) <= 0; angryBirdLarge(2, 44) <= 0; angryBirdLarge(2, 45) <= 0; angryBirdLarge(2, 46) <= 0; angryBirdLarge(2, 47) <= 0; angryBirdLarge(2, 48) <= 0; angryBirdLarge(2, 49) <= 0; angryBirdLarge(2, 50) <= 0; angryBirdLarge(2, 51) <= 0; angryBirdLarge(2, 52) <= 0; angryBirdLarge(2, 53) <= 0; angryBirdLarge(2, 54) <= 0; angryBirdLarge(2, 55) <= 0; angryBirdLarge(2, 56) <= 0; angryBirdLarge(2, 57) <= 0; angryBirdLarge(2, 58) <= 0; angryBirdLarge(2, 59) <= 0; angryBirdLarge(2, 60) <= 0; angryBirdLarge(2, 61) <= 0; angryBirdLarge(2, 62) <= 0; angryBirdLarge(2, 63) <= 0; angryBirdLarge(2, 64) <= 0; angryBirdLarge(2, 65) <= 0; angryBirdLarge(2, 66) <= 0; angryBirdLarge(2, 67) <= 0; angryBirdLarge(2, 68) <= 0; angryBirdLarge(2, 69) <= 0; angryBirdLarge(2, 70) <= 0; angryBirdLarge(2, 71) <= 0; angryBirdLarge(2, 72) <= 5; angryBirdLarge(2, 73) <= 5; angryBirdLarge(2, 74) <= 5; angryBirdLarge(2, 75) <= 5; angryBirdLarge(2, 76) <= 5; angryBirdLarge(2, 77) <= 5; angryBirdLarge(2, 78) <= 5; angryBirdLarge(2, 79) <= 5; angryBirdLarge(2, 80) <= 5; angryBirdLarge(2, 81) <= 5; angryBirdLarge(2, 82) <= 5; angryBirdLarge(2, 83) <= 5; angryBirdLarge(2, 84) <= 5; angryBirdLarge(2, 85) <= 5; angryBirdLarge(2, 86) <= 5; angryBirdLarge(2, 87) <= 5; angryBirdLarge(2, 88) <= 5; angryBirdLarge(2, 89) <= 5; angryBirdLarge(2, 90) <= 0; angryBirdLarge(2, 91) <= 0; angryBirdLarge(2, 92) <= 0; angryBirdLarge(2, 93) <= 0; angryBirdLarge(2, 94) <= 0; angryBirdLarge(2, 95) <= 0; angryBirdLarge(2, 96) <= 0; angryBirdLarge(2, 97) <= 0; angryBirdLarge(2, 98) <= 0; angryBirdLarge(2, 99) <= 0; angryBirdLarge(2, 100) <= 0; angryBirdLarge(2, 101) <= 0; angryBirdLarge(2, 102) <= 0; angryBirdLarge(2, 103) <= 0; angryBirdLarge(2, 104) <= 0; angryBirdLarge(2, 105) <= 0; angryBirdLarge(2, 106) <= 0; angryBirdLarge(2, 107) <= 0; angryBirdLarge(2, 108) <= 0; angryBirdLarge(2, 109) <= 0; angryBirdLarge(2, 110) <= 0; angryBirdLarge(2, 111) <= 0; angryBirdLarge(2, 112) <= 0; angryBirdLarge(2, 113) <= 0; angryBirdLarge(2, 114) <= 0; angryBirdLarge(2, 115) <= 0; angryBirdLarge(2, 116) <= 0; angryBirdLarge(2, 117) <= 0; angryBirdLarge(2, 118) <= 0; angryBirdLarge(2, 119) <= 0; angryBirdLarge(2, 120) <= 0; angryBirdLarge(2, 121) <= 0; angryBirdLarge(2, 122) <= 0; angryBirdLarge(2, 123) <= 0; angryBirdLarge(2, 124) <= 0; angryBirdLarge(2, 125) <= 0; angryBirdLarge(2, 126) <= 0; angryBirdLarge(2, 127) <= 0; angryBirdLarge(2, 128) <= 0; angryBirdLarge(2, 129) <= 0; angryBirdLarge(2, 130) <= 0; angryBirdLarge(2, 131) <= 0; angryBirdLarge(2, 132) <= 0; angryBirdLarge(2, 133) <= 0; angryBirdLarge(2, 134) <= 0; angryBirdLarge(2, 135) <= 0; angryBirdLarge(2, 136) <= 0; angryBirdLarge(2, 137) <= 0; angryBirdLarge(2, 138) <= 0; angryBirdLarge(2, 139) <= 0; angryBirdLarge(2, 140) <= 0; angryBirdLarge(2, 141) <= 0; angryBirdLarge(2, 142) <= 0; angryBirdLarge(2, 143) <= 0; angryBirdLarge(2, 144) <= 0; angryBirdLarge(2, 145) <= 0; angryBirdLarge(2, 146) <= 0; angryBirdLarge(2, 147) <= 0; angryBirdLarge(2, 148) <= 0; angryBirdLarge(2, 149) <= 0; 
angryBirdLarge(3, 0) <= 0; angryBirdLarge(3, 1) <= 0; angryBirdLarge(3, 2) <= 0; angryBirdLarge(3, 3) <= 0; angryBirdLarge(3, 4) <= 0; angryBirdLarge(3, 5) <= 0; angryBirdLarge(3, 6) <= 0; angryBirdLarge(3, 7) <= 0; angryBirdLarge(3, 8) <= 0; angryBirdLarge(3, 9) <= 0; angryBirdLarge(3, 10) <= 0; angryBirdLarge(3, 11) <= 0; angryBirdLarge(3, 12) <= 0; angryBirdLarge(3, 13) <= 0; angryBirdLarge(3, 14) <= 0; angryBirdLarge(3, 15) <= 0; angryBirdLarge(3, 16) <= 0; angryBirdLarge(3, 17) <= 0; angryBirdLarge(3, 18) <= 0; angryBirdLarge(3, 19) <= 0; angryBirdLarge(3, 20) <= 0; angryBirdLarge(3, 21) <= 0; angryBirdLarge(3, 22) <= 0; angryBirdLarge(3, 23) <= 0; angryBirdLarge(3, 24) <= 0; angryBirdLarge(3, 25) <= 0; angryBirdLarge(3, 26) <= 0; angryBirdLarge(3, 27) <= 0; angryBirdLarge(3, 28) <= 0; angryBirdLarge(3, 29) <= 0; angryBirdLarge(3, 30) <= 0; angryBirdLarge(3, 31) <= 0; angryBirdLarge(3, 32) <= 0; angryBirdLarge(3, 33) <= 0; angryBirdLarge(3, 34) <= 0; angryBirdLarge(3, 35) <= 0; angryBirdLarge(3, 36) <= 0; angryBirdLarge(3, 37) <= 0; angryBirdLarge(3, 38) <= 0; angryBirdLarge(3, 39) <= 0; angryBirdLarge(3, 40) <= 0; angryBirdLarge(3, 41) <= 0; angryBirdLarge(3, 42) <= 0; angryBirdLarge(3, 43) <= 0; angryBirdLarge(3, 44) <= 0; angryBirdLarge(3, 45) <= 0; angryBirdLarge(3, 46) <= 0; angryBirdLarge(3, 47) <= 0; angryBirdLarge(3, 48) <= 0; angryBirdLarge(3, 49) <= 0; angryBirdLarge(3, 50) <= 0; angryBirdLarge(3, 51) <= 0; angryBirdLarge(3, 52) <= 0; angryBirdLarge(3, 53) <= 0; angryBirdLarge(3, 54) <= 0; angryBirdLarge(3, 55) <= 0; angryBirdLarge(3, 56) <= 0; angryBirdLarge(3, 57) <= 0; angryBirdLarge(3, 58) <= 0; angryBirdLarge(3, 59) <= 0; angryBirdLarge(3, 60) <= 0; angryBirdLarge(3, 61) <= 0; angryBirdLarge(3, 62) <= 0; angryBirdLarge(3, 63) <= 0; angryBirdLarge(3, 64) <= 0; angryBirdLarge(3, 65) <= 0; angryBirdLarge(3, 66) <= 0; angryBirdLarge(3, 67) <= 0; angryBirdLarge(3, 68) <= 0; angryBirdLarge(3, 69) <= 0; angryBirdLarge(3, 70) <= 0; angryBirdLarge(3, 71) <= 0; angryBirdLarge(3, 72) <= 5; angryBirdLarge(3, 73) <= 5; angryBirdLarge(3, 74) <= 5; angryBirdLarge(3, 75) <= 5; angryBirdLarge(3, 76) <= 5; angryBirdLarge(3, 77) <= 5; angryBirdLarge(3, 78) <= 5; angryBirdLarge(3, 79) <= 5; angryBirdLarge(3, 80) <= 5; angryBirdLarge(3, 81) <= 5; angryBirdLarge(3, 82) <= 5; angryBirdLarge(3, 83) <= 5; angryBirdLarge(3, 84) <= 5; angryBirdLarge(3, 85) <= 5; angryBirdLarge(3, 86) <= 5; angryBirdLarge(3, 87) <= 5; angryBirdLarge(3, 88) <= 5; angryBirdLarge(3, 89) <= 5; angryBirdLarge(3, 90) <= 0; angryBirdLarge(3, 91) <= 0; angryBirdLarge(3, 92) <= 0; angryBirdLarge(3, 93) <= 0; angryBirdLarge(3, 94) <= 0; angryBirdLarge(3, 95) <= 0; angryBirdLarge(3, 96) <= 0; angryBirdLarge(3, 97) <= 0; angryBirdLarge(3, 98) <= 0; angryBirdLarge(3, 99) <= 0; angryBirdLarge(3, 100) <= 0; angryBirdLarge(3, 101) <= 0; angryBirdLarge(3, 102) <= 0; angryBirdLarge(3, 103) <= 0; angryBirdLarge(3, 104) <= 0; angryBirdLarge(3, 105) <= 0; angryBirdLarge(3, 106) <= 0; angryBirdLarge(3, 107) <= 0; angryBirdLarge(3, 108) <= 0; angryBirdLarge(3, 109) <= 0; angryBirdLarge(3, 110) <= 0; angryBirdLarge(3, 111) <= 0; angryBirdLarge(3, 112) <= 0; angryBirdLarge(3, 113) <= 0; angryBirdLarge(3, 114) <= 0; angryBirdLarge(3, 115) <= 0; angryBirdLarge(3, 116) <= 0; angryBirdLarge(3, 117) <= 0; angryBirdLarge(3, 118) <= 0; angryBirdLarge(3, 119) <= 0; angryBirdLarge(3, 120) <= 0; angryBirdLarge(3, 121) <= 0; angryBirdLarge(3, 122) <= 0; angryBirdLarge(3, 123) <= 0; angryBirdLarge(3, 124) <= 0; angryBirdLarge(3, 125) <= 0; angryBirdLarge(3, 126) <= 0; angryBirdLarge(3, 127) <= 0; angryBirdLarge(3, 128) <= 0; angryBirdLarge(3, 129) <= 0; angryBirdLarge(3, 130) <= 0; angryBirdLarge(3, 131) <= 0; angryBirdLarge(3, 132) <= 0; angryBirdLarge(3, 133) <= 0; angryBirdLarge(3, 134) <= 0; angryBirdLarge(3, 135) <= 0; angryBirdLarge(3, 136) <= 0; angryBirdLarge(3, 137) <= 0; angryBirdLarge(3, 138) <= 0; angryBirdLarge(3, 139) <= 0; angryBirdLarge(3, 140) <= 0; angryBirdLarge(3, 141) <= 0; angryBirdLarge(3, 142) <= 0; angryBirdLarge(3, 143) <= 0; angryBirdLarge(3, 144) <= 0; angryBirdLarge(3, 145) <= 0; angryBirdLarge(3, 146) <= 0; angryBirdLarge(3, 147) <= 0; angryBirdLarge(3, 148) <= 0; angryBirdLarge(3, 149) <= 0; 
angryBirdLarge(4, 0) <= 0; angryBirdLarge(4, 1) <= 0; angryBirdLarge(4, 2) <= 0; angryBirdLarge(4, 3) <= 0; angryBirdLarge(4, 4) <= 0; angryBirdLarge(4, 5) <= 0; angryBirdLarge(4, 6) <= 0; angryBirdLarge(4, 7) <= 0; angryBirdLarge(4, 8) <= 0; angryBirdLarge(4, 9) <= 0; angryBirdLarge(4, 10) <= 0; angryBirdLarge(4, 11) <= 0; angryBirdLarge(4, 12) <= 0; angryBirdLarge(4, 13) <= 0; angryBirdLarge(4, 14) <= 0; angryBirdLarge(4, 15) <= 0; angryBirdLarge(4, 16) <= 0; angryBirdLarge(4, 17) <= 0; angryBirdLarge(4, 18) <= 0; angryBirdLarge(4, 19) <= 0; angryBirdLarge(4, 20) <= 0; angryBirdLarge(4, 21) <= 0; angryBirdLarge(4, 22) <= 0; angryBirdLarge(4, 23) <= 0; angryBirdLarge(4, 24) <= 0; angryBirdLarge(4, 25) <= 0; angryBirdLarge(4, 26) <= 0; angryBirdLarge(4, 27) <= 0; angryBirdLarge(4, 28) <= 0; angryBirdLarge(4, 29) <= 0; angryBirdLarge(4, 30) <= 0; angryBirdLarge(4, 31) <= 0; angryBirdLarge(4, 32) <= 0; angryBirdLarge(4, 33) <= 0; angryBirdLarge(4, 34) <= 0; angryBirdLarge(4, 35) <= 0; angryBirdLarge(4, 36) <= 0; angryBirdLarge(4, 37) <= 0; angryBirdLarge(4, 38) <= 0; angryBirdLarge(4, 39) <= 0; angryBirdLarge(4, 40) <= 0; angryBirdLarge(4, 41) <= 0; angryBirdLarge(4, 42) <= 0; angryBirdLarge(4, 43) <= 0; angryBirdLarge(4, 44) <= 0; angryBirdLarge(4, 45) <= 0; angryBirdLarge(4, 46) <= 0; angryBirdLarge(4, 47) <= 0; angryBirdLarge(4, 48) <= 0; angryBirdLarge(4, 49) <= 0; angryBirdLarge(4, 50) <= 0; angryBirdLarge(4, 51) <= 0; angryBirdLarge(4, 52) <= 0; angryBirdLarge(4, 53) <= 0; angryBirdLarge(4, 54) <= 0; angryBirdLarge(4, 55) <= 0; angryBirdLarge(4, 56) <= 0; angryBirdLarge(4, 57) <= 0; angryBirdLarge(4, 58) <= 0; angryBirdLarge(4, 59) <= 0; angryBirdLarge(4, 60) <= 0; angryBirdLarge(4, 61) <= 0; angryBirdLarge(4, 62) <= 0; angryBirdLarge(4, 63) <= 0; angryBirdLarge(4, 64) <= 0; angryBirdLarge(4, 65) <= 0; angryBirdLarge(4, 66) <= 0; angryBirdLarge(4, 67) <= 0; angryBirdLarge(4, 68) <= 0; angryBirdLarge(4, 69) <= 0; angryBirdLarge(4, 70) <= 0; angryBirdLarge(4, 71) <= 0; angryBirdLarge(4, 72) <= 5; angryBirdLarge(4, 73) <= 5; angryBirdLarge(4, 74) <= 5; angryBirdLarge(4, 75) <= 5; angryBirdLarge(4, 76) <= 5; angryBirdLarge(4, 77) <= 5; angryBirdLarge(4, 78) <= 5; angryBirdLarge(4, 79) <= 5; angryBirdLarge(4, 80) <= 5; angryBirdLarge(4, 81) <= 5; angryBirdLarge(4, 82) <= 5; angryBirdLarge(4, 83) <= 5; angryBirdLarge(4, 84) <= 5; angryBirdLarge(4, 85) <= 5; angryBirdLarge(4, 86) <= 5; angryBirdLarge(4, 87) <= 5; angryBirdLarge(4, 88) <= 5; angryBirdLarge(4, 89) <= 5; angryBirdLarge(4, 90) <= 0; angryBirdLarge(4, 91) <= 0; angryBirdLarge(4, 92) <= 0; angryBirdLarge(4, 93) <= 0; angryBirdLarge(4, 94) <= 0; angryBirdLarge(4, 95) <= 0; angryBirdLarge(4, 96) <= 0; angryBirdLarge(4, 97) <= 0; angryBirdLarge(4, 98) <= 0; angryBirdLarge(4, 99) <= 0; angryBirdLarge(4, 100) <= 0; angryBirdLarge(4, 101) <= 0; angryBirdLarge(4, 102) <= 0; angryBirdLarge(4, 103) <= 0; angryBirdLarge(4, 104) <= 0; angryBirdLarge(4, 105) <= 0; angryBirdLarge(4, 106) <= 0; angryBirdLarge(4, 107) <= 0; angryBirdLarge(4, 108) <= 0; angryBirdLarge(4, 109) <= 0; angryBirdLarge(4, 110) <= 0; angryBirdLarge(4, 111) <= 0; angryBirdLarge(4, 112) <= 0; angryBirdLarge(4, 113) <= 0; angryBirdLarge(4, 114) <= 0; angryBirdLarge(4, 115) <= 0; angryBirdLarge(4, 116) <= 0; angryBirdLarge(4, 117) <= 0; angryBirdLarge(4, 118) <= 0; angryBirdLarge(4, 119) <= 0; angryBirdLarge(4, 120) <= 0; angryBirdLarge(4, 121) <= 0; angryBirdLarge(4, 122) <= 0; angryBirdLarge(4, 123) <= 0; angryBirdLarge(4, 124) <= 0; angryBirdLarge(4, 125) <= 0; angryBirdLarge(4, 126) <= 0; angryBirdLarge(4, 127) <= 0; angryBirdLarge(4, 128) <= 0; angryBirdLarge(4, 129) <= 0; angryBirdLarge(4, 130) <= 0; angryBirdLarge(4, 131) <= 0; angryBirdLarge(4, 132) <= 0; angryBirdLarge(4, 133) <= 0; angryBirdLarge(4, 134) <= 0; angryBirdLarge(4, 135) <= 0; angryBirdLarge(4, 136) <= 0; angryBirdLarge(4, 137) <= 0; angryBirdLarge(4, 138) <= 0; angryBirdLarge(4, 139) <= 0; angryBirdLarge(4, 140) <= 0; angryBirdLarge(4, 141) <= 0; angryBirdLarge(4, 142) <= 0; angryBirdLarge(4, 143) <= 0; angryBirdLarge(4, 144) <= 0; angryBirdLarge(4, 145) <= 0; angryBirdLarge(4, 146) <= 0; angryBirdLarge(4, 147) <= 0; angryBirdLarge(4, 148) <= 0; angryBirdLarge(4, 149) <= 0; 
angryBirdLarge(5, 0) <= 0; angryBirdLarge(5, 1) <= 0; angryBirdLarge(5, 2) <= 0; angryBirdLarge(5, 3) <= 0; angryBirdLarge(5, 4) <= 0; angryBirdLarge(5, 5) <= 0; angryBirdLarge(5, 6) <= 0; angryBirdLarge(5, 7) <= 0; angryBirdLarge(5, 8) <= 0; angryBirdLarge(5, 9) <= 0; angryBirdLarge(5, 10) <= 0; angryBirdLarge(5, 11) <= 0; angryBirdLarge(5, 12) <= 0; angryBirdLarge(5, 13) <= 0; angryBirdLarge(5, 14) <= 0; angryBirdLarge(5, 15) <= 0; angryBirdLarge(5, 16) <= 0; angryBirdLarge(5, 17) <= 0; angryBirdLarge(5, 18) <= 0; angryBirdLarge(5, 19) <= 0; angryBirdLarge(5, 20) <= 0; angryBirdLarge(5, 21) <= 0; angryBirdLarge(5, 22) <= 0; angryBirdLarge(5, 23) <= 0; angryBirdLarge(5, 24) <= 0; angryBirdLarge(5, 25) <= 0; angryBirdLarge(5, 26) <= 0; angryBirdLarge(5, 27) <= 0; angryBirdLarge(5, 28) <= 0; angryBirdLarge(5, 29) <= 0; angryBirdLarge(5, 30) <= 0; angryBirdLarge(5, 31) <= 0; angryBirdLarge(5, 32) <= 0; angryBirdLarge(5, 33) <= 0; angryBirdLarge(5, 34) <= 0; angryBirdLarge(5, 35) <= 0; angryBirdLarge(5, 36) <= 0; angryBirdLarge(5, 37) <= 0; angryBirdLarge(5, 38) <= 0; angryBirdLarge(5, 39) <= 0; angryBirdLarge(5, 40) <= 0; angryBirdLarge(5, 41) <= 0; angryBirdLarge(5, 42) <= 0; angryBirdLarge(5, 43) <= 0; angryBirdLarge(5, 44) <= 0; angryBirdLarge(5, 45) <= 0; angryBirdLarge(5, 46) <= 0; angryBirdLarge(5, 47) <= 0; angryBirdLarge(5, 48) <= 0; angryBirdLarge(5, 49) <= 0; angryBirdLarge(5, 50) <= 0; angryBirdLarge(5, 51) <= 0; angryBirdLarge(5, 52) <= 0; angryBirdLarge(5, 53) <= 0; angryBirdLarge(5, 54) <= 0; angryBirdLarge(5, 55) <= 0; angryBirdLarge(5, 56) <= 0; angryBirdLarge(5, 57) <= 0; angryBirdLarge(5, 58) <= 0; angryBirdLarge(5, 59) <= 0; angryBirdLarge(5, 60) <= 0; angryBirdLarge(5, 61) <= 0; angryBirdLarge(5, 62) <= 0; angryBirdLarge(5, 63) <= 0; angryBirdLarge(5, 64) <= 0; angryBirdLarge(5, 65) <= 0; angryBirdLarge(5, 66) <= 0; angryBirdLarge(5, 67) <= 0; angryBirdLarge(5, 68) <= 0; angryBirdLarge(5, 69) <= 0; angryBirdLarge(5, 70) <= 0; angryBirdLarge(5, 71) <= 0; angryBirdLarge(5, 72) <= 5; angryBirdLarge(5, 73) <= 5; angryBirdLarge(5, 74) <= 5; angryBirdLarge(5, 75) <= 5; angryBirdLarge(5, 76) <= 5; angryBirdLarge(5, 77) <= 5; angryBirdLarge(5, 78) <= 5; angryBirdLarge(5, 79) <= 5; angryBirdLarge(5, 80) <= 5; angryBirdLarge(5, 81) <= 5; angryBirdLarge(5, 82) <= 5; angryBirdLarge(5, 83) <= 5; angryBirdLarge(5, 84) <= 5; angryBirdLarge(5, 85) <= 5; angryBirdLarge(5, 86) <= 5; angryBirdLarge(5, 87) <= 5; angryBirdLarge(5, 88) <= 5; angryBirdLarge(5, 89) <= 5; angryBirdLarge(5, 90) <= 0; angryBirdLarge(5, 91) <= 0; angryBirdLarge(5, 92) <= 0; angryBirdLarge(5, 93) <= 0; angryBirdLarge(5, 94) <= 0; angryBirdLarge(5, 95) <= 0; angryBirdLarge(5, 96) <= 0; angryBirdLarge(5, 97) <= 0; angryBirdLarge(5, 98) <= 0; angryBirdLarge(5, 99) <= 0; angryBirdLarge(5, 100) <= 0; angryBirdLarge(5, 101) <= 0; angryBirdLarge(5, 102) <= 0; angryBirdLarge(5, 103) <= 0; angryBirdLarge(5, 104) <= 0; angryBirdLarge(5, 105) <= 0; angryBirdLarge(5, 106) <= 0; angryBirdLarge(5, 107) <= 0; angryBirdLarge(5, 108) <= 0; angryBirdLarge(5, 109) <= 0; angryBirdLarge(5, 110) <= 0; angryBirdLarge(5, 111) <= 0; angryBirdLarge(5, 112) <= 0; angryBirdLarge(5, 113) <= 0; angryBirdLarge(5, 114) <= 0; angryBirdLarge(5, 115) <= 0; angryBirdLarge(5, 116) <= 0; angryBirdLarge(5, 117) <= 0; angryBirdLarge(5, 118) <= 0; angryBirdLarge(5, 119) <= 0; angryBirdLarge(5, 120) <= 0; angryBirdLarge(5, 121) <= 0; angryBirdLarge(5, 122) <= 0; angryBirdLarge(5, 123) <= 0; angryBirdLarge(5, 124) <= 0; angryBirdLarge(5, 125) <= 0; angryBirdLarge(5, 126) <= 0; angryBirdLarge(5, 127) <= 0; angryBirdLarge(5, 128) <= 0; angryBirdLarge(5, 129) <= 0; angryBirdLarge(5, 130) <= 0; angryBirdLarge(5, 131) <= 0; angryBirdLarge(5, 132) <= 0; angryBirdLarge(5, 133) <= 0; angryBirdLarge(5, 134) <= 0; angryBirdLarge(5, 135) <= 0; angryBirdLarge(5, 136) <= 0; angryBirdLarge(5, 137) <= 0; angryBirdLarge(5, 138) <= 0; angryBirdLarge(5, 139) <= 0; angryBirdLarge(5, 140) <= 0; angryBirdLarge(5, 141) <= 0; angryBirdLarge(5, 142) <= 0; angryBirdLarge(5, 143) <= 0; angryBirdLarge(5, 144) <= 0; angryBirdLarge(5, 145) <= 0; angryBirdLarge(5, 146) <= 0; angryBirdLarge(5, 147) <= 0; angryBirdLarge(5, 148) <= 0; angryBirdLarge(5, 149) <= 0; 
angryBirdLarge(6, 0) <= 0; angryBirdLarge(6, 1) <= 0; angryBirdLarge(6, 2) <= 0; angryBirdLarge(6, 3) <= 0; angryBirdLarge(6, 4) <= 0; angryBirdLarge(6, 5) <= 0; angryBirdLarge(6, 6) <= 0; angryBirdLarge(6, 7) <= 0; angryBirdLarge(6, 8) <= 0; angryBirdLarge(6, 9) <= 0; angryBirdLarge(6, 10) <= 0; angryBirdLarge(6, 11) <= 0; angryBirdLarge(6, 12) <= 0; angryBirdLarge(6, 13) <= 0; angryBirdLarge(6, 14) <= 0; angryBirdLarge(6, 15) <= 0; angryBirdLarge(6, 16) <= 0; angryBirdLarge(6, 17) <= 0; angryBirdLarge(6, 18) <= 0; angryBirdLarge(6, 19) <= 0; angryBirdLarge(6, 20) <= 0; angryBirdLarge(6, 21) <= 0; angryBirdLarge(6, 22) <= 0; angryBirdLarge(6, 23) <= 0; angryBirdLarge(6, 24) <= 0; angryBirdLarge(6, 25) <= 0; angryBirdLarge(6, 26) <= 0; angryBirdLarge(6, 27) <= 0; angryBirdLarge(6, 28) <= 0; angryBirdLarge(6, 29) <= 0; angryBirdLarge(6, 30) <= 0; angryBirdLarge(6, 31) <= 0; angryBirdLarge(6, 32) <= 0; angryBirdLarge(6, 33) <= 0; angryBirdLarge(6, 34) <= 0; angryBirdLarge(6, 35) <= 0; angryBirdLarge(6, 36) <= 0; angryBirdLarge(6, 37) <= 0; angryBirdLarge(6, 38) <= 0; angryBirdLarge(6, 39) <= 0; angryBirdLarge(6, 40) <= 0; angryBirdLarge(6, 41) <= 0; angryBirdLarge(6, 42) <= 0; angryBirdLarge(6, 43) <= 0; angryBirdLarge(6, 44) <= 0; angryBirdLarge(6, 45) <= 0; angryBirdLarge(6, 46) <= 0; angryBirdLarge(6, 47) <= 0; angryBirdLarge(6, 48) <= 0; angryBirdLarge(6, 49) <= 0; angryBirdLarge(6, 50) <= 0; angryBirdLarge(6, 51) <= 0; angryBirdLarge(6, 52) <= 0; angryBirdLarge(6, 53) <= 0; angryBirdLarge(6, 54) <= 0; angryBirdLarge(6, 55) <= 0; angryBirdLarge(6, 56) <= 0; angryBirdLarge(6, 57) <= 0; angryBirdLarge(6, 58) <= 0; angryBirdLarge(6, 59) <= 0; angryBirdLarge(6, 60) <= 0; angryBirdLarge(6, 61) <= 0; angryBirdLarge(6, 62) <= 0; angryBirdLarge(6, 63) <= 0; angryBirdLarge(6, 64) <= 0; angryBirdLarge(6, 65) <= 0; angryBirdLarge(6, 66) <= 5; angryBirdLarge(6, 67) <= 5; angryBirdLarge(6, 68) <= 5; angryBirdLarge(6, 69) <= 5; angryBirdLarge(6, 70) <= 5; angryBirdLarge(6, 71) <= 5; angryBirdLarge(6, 72) <= 4; angryBirdLarge(6, 73) <= 4; angryBirdLarge(6, 74) <= 4; angryBirdLarge(6, 75) <= 4; angryBirdLarge(6, 76) <= 4; angryBirdLarge(6, 77) <= 4; angryBirdLarge(6, 78) <= 4; angryBirdLarge(6, 79) <= 4; angryBirdLarge(6, 80) <= 4; angryBirdLarge(6, 81) <= 4; angryBirdLarge(6, 82) <= 4; angryBirdLarge(6, 83) <= 4; angryBirdLarge(6, 84) <= 4; angryBirdLarge(6, 85) <= 4; angryBirdLarge(6, 86) <= 4; angryBirdLarge(6, 87) <= 4; angryBirdLarge(6, 88) <= 4; angryBirdLarge(6, 89) <= 4; angryBirdLarge(6, 90) <= 5; angryBirdLarge(6, 91) <= 5; angryBirdLarge(6, 92) <= 5; angryBirdLarge(6, 93) <= 5; angryBirdLarge(6, 94) <= 5; angryBirdLarge(6, 95) <= 5; angryBirdLarge(6, 96) <= 0; angryBirdLarge(6, 97) <= 0; angryBirdLarge(6, 98) <= 0; angryBirdLarge(6, 99) <= 0; angryBirdLarge(6, 100) <= 0; angryBirdLarge(6, 101) <= 0; angryBirdLarge(6, 102) <= 0; angryBirdLarge(6, 103) <= 0; angryBirdLarge(6, 104) <= 0; angryBirdLarge(6, 105) <= 0; angryBirdLarge(6, 106) <= 0; angryBirdLarge(6, 107) <= 0; angryBirdLarge(6, 108) <= 0; angryBirdLarge(6, 109) <= 0; angryBirdLarge(6, 110) <= 0; angryBirdLarge(6, 111) <= 0; angryBirdLarge(6, 112) <= 0; angryBirdLarge(6, 113) <= 0; angryBirdLarge(6, 114) <= 0; angryBirdLarge(6, 115) <= 0; angryBirdLarge(6, 116) <= 0; angryBirdLarge(6, 117) <= 0; angryBirdLarge(6, 118) <= 0; angryBirdLarge(6, 119) <= 0; angryBirdLarge(6, 120) <= 0; angryBirdLarge(6, 121) <= 0; angryBirdLarge(6, 122) <= 0; angryBirdLarge(6, 123) <= 0; angryBirdLarge(6, 124) <= 0; angryBirdLarge(6, 125) <= 0; angryBirdLarge(6, 126) <= 0; angryBirdLarge(6, 127) <= 0; angryBirdLarge(6, 128) <= 0; angryBirdLarge(6, 129) <= 0; angryBirdLarge(6, 130) <= 0; angryBirdLarge(6, 131) <= 0; angryBirdLarge(6, 132) <= 0; angryBirdLarge(6, 133) <= 0; angryBirdLarge(6, 134) <= 0; angryBirdLarge(6, 135) <= 0; angryBirdLarge(6, 136) <= 0; angryBirdLarge(6, 137) <= 0; angryBirdLarge(6, 138) <= 0; angryBirdLarge(6, 139) <= 0; angryBirdLarge(6, 140) <= 0; angryBirdLarge(6, 141) <= 0; angryBirdLarge(6, 142) <= 0; angryBirdLarge(6, 143) <= 0; angryBirdLarge(6, 144) <= 0; angryBirdLarge(6, 145) <= 0; angryBirdLarge(6, 146) <= 0; angryBirdLarge(6, 147) <= 0; angryBirdLarge(6, 148) <= 0; angryBirdLarge(6, 149) <= 0; 
angryBirdLarge(7, 0) <= 0; angryBirdLarge(7, 1) <= 0; angryBirdLarge(7, 2) <= 0; angryBirdLarge(7, 3) <= 0; angryBirdLarge(7, 4) <= 0; angryBirdLarge(7, 5) <= 0; angryBirdLarge(7, 6) <= 0; angryBirdLarge(7, 7) <= 0; angryBirdLarge(7, 8) <= 0; angryBirdLarge(7, 9) <= 0; angryBirdLarge(7, 10) <= 0; angryBirdLarge(7, 11) <= 0; angryBirdLarge(7, 12) <= 0; angryBirdLarge(7, 13) <= 0; angryBirdLarge(7, 14) <= 0; angryBirdLarge(7, 15) <= 0; angryBirdLarge(7, 16) <= 0; angryBirdLarge(7, 17) <= 0; angryBirdLarge(7, 18) <= 0; angryBirdLarge(7, 19) <= 0; angryBirdLarge(7, 20) <= 0; angryBirdLarge(7, 21) <= 0; angryBirdLarge(7, 22) <= 0; angryBirdLarge(7, 23) <= 0; angryBirdLarge(7, 24) <= 0; angryBirdLarge(7, 25) <= 0; angryBirdLarge(7, 26) <= 0; angryBirdLarge(7, 27) <= 0; angryBirdLarge(7, 28) <= 0; angryBirdLarge(7, 29) <= 0; angryBirdLarge(7, 30) <= 0; angryBirdLarge(7, 31) <= 0; angryBirdLarge(7, 32) <= 0; angryBirdLarge(7, 33) <= 0; angryBirdLarge(7, 34) <= 0; angryBirdLarge(7, 35) <= 0; angryBirdLarge(7, 36) <= 0; angryBirdLarge(7, 37) <= 0; angryBirdLarge(7, 38) <= 0; angryBirdLarge(7, 39) <= 0; angryBirdLarge(7, 40) <= 0; angryBirdLarge(7, 41) <= 0; angryBirdLarge(7, 42) <= 0; angryBirdLarge(7, 43) <= 0; angryBirdLarge(7, 44) <= 0; angryBirdLarge(7, 45) <= 0; angryBirdLarge(7, 46) <= 0; angryBirdLarge(7, 47) <= 0; angryBirdLarge(7, 48) <= 0; angryBirdLarge(7, 49) <= 0; angryBirdLarge(7, 50) <= 0; angryBirdLarge(7, 51) <= 0; angryBirdLarge(7, 52) <= 0; angryBirdLarge(7, 53) <= 0; angryBirdLarge(7, 54) <= 0; angryBirdLarge(7, 55) <= 0; angryBirdLarge(7, 56) <= 0; angryBirdLarge(7, 57) <= 0; angryBirdLarge(7, 58) <= 0; angryBirdLarge(7, 59) <= 0; angryBirdLarge(7, 60) <= 0; angryBirdLarge(7, 61) <= 0; angryBirdLarge(7, 62) <= 0; angryBirdLarge(7, 63) <= 0; angryBirdLarge(7, 64) <= 0; angryBirdLarge(7, 65) <= 0; angryBirdLarge(7, 66) <= 5; angryBirdLarge(7, 67) <= 5; angryBirdLarge(7, 68) <= 5; angryBirdLarge(7, 69) <= 5; angryBirdLarge(7, 70) <= 5; angryBirdLarge(7, 71) <= 5; angryBirdLarge(7, 72) <= 4; angryBirdLarge(7, 73) <= 4; angryBirdLarge(7, 74) <= 4; angryBirdLarge(7, 75) <= 4; angryBirdLarge(7, 76) <= 4; angryBirdLarge(7, 77) <= 4; angryBirdLarge(7, 78) <= 4; angryBirdLarge(7, 79) <= 4; angryBirdLarge(7, 80) <= 4; angryBirdLarge(7, 81) <= 4; angryBirdLarge(7, 82) <= 4; angryBirdLarge(7, 83) <= 4; angryBirdLarge(7, 84) <= 4; angryBirdLarge(7, 85) <= 4; angryBirdLarge(7, 86) <= 4; angryBirdLarge(7, 87) <= 4; angryBirdLarge(7, 88) <= 4; angryBirdLarge(7, 89) <= 4; angryBirdLarge(7, 90) <= 5; angryBirdLarge(7, 91) <= 5; angryBirdLarge(7, 92) <= 5; angryBirdLarge(7, 93) <= 5; angryBirdLarge(7, 94) <= 5; angryBirdLarge(7, 95) <= 5; angryBirdLarge(7, 96) <= 0; angryBirdLarge(7, 97) <= 0; angryBirdLarge(7, 98) <= 0; angryBirdLarge(7, 99) <= 0; angryBirdLarge(7, 100) <= 0; angryBirdLarge(7, 101) <= 0; angryBirdLarge(7, 102) <= 0; angryBirdLarge(7, 103) <= 0; angryBirdLarge(7, 104) <= 0; angryBirdLarge(7, 105) <= 0; angryBirdLarge(7, 106) <= 0; angryBirdLarge(7, 107) <= 0; angryBirdLarge(7, 108) <= 0; angryBirdLarge(7, 109) <= 0; angryBirdLarge(7, 110) <= 0; angryBirdLarge(7, 111) <= 0; angryBirdLarge(7, 112) <= 0; angryBirdLarge(7, 113) <= 0; angryBirdLarge(7, 114) <= 0; angryBirdLarge(7, 115) <= 0; angryBirdLarge(7, 116) <= 0; angryBirdLarge(7, 117) <= 0; angryBirdLarge(7, 118) <= 0; angryBirdLarge(7, 119) <= 0; angryBirdLarge(7, 120) <= 0; angryBirdLarge(7, 121) <= 0; angryBirdLarge(7, 122) <= 0; angryBirdLarge(7, 123) <= 0; angryBirdLarge(7, 124) <= 0; angryBirdLarge(7, 125) <= 0; angryBirdLarge(7, 126) <= 0; angryBirdLarge(7, 127) <= 0; angryBirdLarge(7, 128) <= 0; angryBirdLarge(7, 129) <= 0; angryBirdLarge(7, 130) <= 0; angryBirdLarge(7, 131) <= 0; angryBirdLarge(7, 132) <= 0; angryBirdLarge(7, 133) <= 0; angryBirdLarge(7, 134) <= 0; angryBirdLarge(7, 135) <= 0; angryBirdLarge(7, 136) <= 0; angryBirdLarge(7, 137) <= 0; angryBirdLarge(7, 138) <= 0; angryBirdLarge(7, 139) <= 0; angryBirdLarge(7, 140) <= 0; angryBirdLarge(7, 141) <= 0; angryBirdLarge(7, 142) <= 0; angryBirdLarge(7, 143) <= 0; angryBirdLarge(7, 144) <= 0; angryBirdLarge(7, 145) <= 0; angryBirdLarge(7, 146) <= 0; angryBirdLarge(7, 147) <= 0; angryBirdLarge(7, 148) <= 0; angryBirdLarge(7, 149) <= 0; 
angryBirdLarge(8, 0) <= 0; angryBirdLarge(8, 1) <= 0; angryBirdLarge(8, 2) <= 0; angryBirdLarge(8, 3) <= 0; angryBirdLarge(8, 4) <= 0; angryBirdLarge(8, 5) <= 0; angryBirdLarge(8, 6) <= 0; angryBirdLarge(8, 7) <= 0; angryBirdLarge(8, 8) <= 0; angryBirdLarge(8, 9) <= 0; angryBirdLarge(8, 10) <= 0; angryBirdLarge(8, 11) <= 0; angryBirdLarge(8, 12) <= 0; angryBirdLarge(8, 13) <= 0; angryBirdLarge(8, 14) <= 0; angryBirdLarge(8, 15) <= 0; angryBirdLarge(8, 16) <= 0; angryBirdLarge(8, 17) <= 0; angryBirdLarge(8, 18) <= 0; angryBirdLarge(8, 19) <= 0; angryBirdLarge(8, 20) <= 0; angryBirdLarge(8, 21) <= 0; angryBirdLarge(8, 22) <= 0; angryBirdLarge(8, 23) <= 0; angryBirdLarge(8, 24) <= 0; angryBirdLarge(8, 25) <= 0; angryBirdLarge(8, 26) <= 0; angryBirdLarge(8, 27) <= 0; angryBirdLarge(8, 28) <= 0; angryBirdLarge(8, 29) <= 0; angryBirdLarge(8, 30) <= 0; angryBirdLarge(8, 31) <= 0; angryBirdLarge(8, 32) <= 0; angryBirdLarge(8, 33) <= 0; angryBirdLarge(8, 34) <= 0; angryBirdLarge(8, 35) <= 0; angryBirdLarge(8, 36) <= 0; angryBirdLarge(8, 37) <= 0; angryBirdLarge(8, 38) <= 0; angryBirdLarge(8, 39) <= 0; angryBirdLarge(8, 40) <= 0; angryBirdLarge(8, 41) <= 0; angryBirdLarge(8, 42) <= 0; angryBirdLarge(8, 43) <= 0; angryBirdLarge(8, 44) <= 0; angryBirdLarge(8, 45) <= 0; angryBirdLarge(8, 46) <= 0; angryBirdLarge(8, 47) <= 0; angryBirdLarge(8, 48) <= 0; angryBirdLarge(8, 49) <= 0; angryBirdLarge(8, 50) <= 0; angryBirdLarge(8, 51) <= 0; angryBirdLarge(8, 52) <= 0; angryBirdLarge(8, 53) <= 0; angryBirdLarge(8, 54) <= 0; angryBirdLarge(8, 55) <= 0; angryBirdLarge(8, 56) <= 0; angryBirdLarge(8, 57) <= 0; angryBirdLarge(8, 58) <= 0; angryBirdLarge(8, 59) <= 0; angryBirdLarge(8, 60) <= 0; angryBirdLarge(8, 61) <= 0; angryBirdLarge(8, 62) <= 0; angryBirdLarge(8, 63) <= 0; angryBirdLarge(8, 64) <= 0; angryBirdLarge(8, 65) <= 0; angryBirdLarge(8, 66) <= 5; angryBirdLarge(8, 67) <= 5; angryBirdLarge(8, 68) <= 5; angryBirdLarge(8, 69) <= 5; angryBirdLarge(8, 70) <= 5; angryBirdLarge(8, 71) <= 5; angryBirdLarge(8, 72) <= 4; angryBirdLarge(8, 73) <= 4; angryBirdLarge(8, 74) <= 4; angryBirdLarge(8, 75) <= 4; angryBirdLarge(8, 76) <= 4; angryBirdLarge(8, 77) <= 4; angryBirdLarge(8, 78) <= 4; angryBirdLarge(8, 79) <= 4; angryBirdLarge(8, 80) <= 4; angryBirdLarge(8, 81) <= 4; angryBirdLarge(8, 82) <= 4; angryBirdLarge(8, 83) <= 4; angryBirdLarge(8, 84) <= 4; angryBirdLarge(8, 85) <= 4; angryBirdLarge(8, 86) <= 4; angryBirdLarge(8, 87) <= 4; angryBirdLarge(8, 88) <= 4; angryBirdLarge(8, 89) <= 4; angryBirdLarge(8, 90) <= 5; angryBirdLarge(8, 91) <= 5; angryBirdLarge(8, 92) <= 5; angryBirdLarge(8, 93) <= 5; angryBirdLarge(8, 94) <= 5; angryBirdLarge(8, 95) <= 5; angryBirdLarge(8, 96) <= 0; angryBirdLarge(8, 97) <= 0; angryBirdLarge(8, 98) <= 0; angryBirdLarge(8, 99) <= 0; angryBirdLarge(8, 100) <= 0; angryBirdLarge(8, 101) <= 0; angryBirdLarge(8, 102) <= 0; angryBirdLarge(8, 103) <= 0; angryBirdLarge(8, 104) <= 0; angryBirdLarge(8, 105) <= 0; angryBirdLarge(8, 106) <= 0; angryBirdLarge(8, 107) <= 0; angryBirdLarge(8, 108) <= 0; angryBirdLarge(8, 109) <= 0; angryBirdLarge(8, 110) <= 0; angryBirdLarge(8, 111) <= 0; angryBirdLarge(8, 112) <= 0; angryBirdLarge(8, 113) <= 0; angryBirdLarge(8, 114) <= 0; angryBirdLarge(8, 115) <= 0; angryBirdLarge(8, 116) <= 0; angryBirdLarge(8, 117) <= 0; angryBirdLarge(8, 118) <= 0; angryBirdLarge(8, 119) <= 0; angryBirdLarge(8, 120) <= 0; angryBirdLarge(8, 121) <= 0; angryBirdLarge(8, 122) <= 0; angryBirdLarge(8, 123) <= 0; angryBirdLarge(8, 124) <= 0; angryBirdLarge(8, 125) <= 0; angryBirdLarge(8, 126) <= 0; angryBirdLarge(8, 127) <= 0; angryBirdLarge(8, 128) <= 0; angryBirdLarge(8, 129) <= 0; angryBirdLarge(8, 130) <= 0; angryBirdLarge(8, 131) <= 0; angryBirdLarge(8, 132) <= 0; angryBirdLarge(8, 133) <= 0; angryBirdLarge(8, 134) <= 0; angryBirdLarge(8, 135) <= 0; angryBirdLarge(8, 136) <= 0; angryBirdLarge(8, 137) <= 0; angryBirdLarge(8, 138) <= 0; angryBirdLarge(8, 139) <= 0; angryBirdLarge(8, 140) <= 0; angryBirdLarge(8, 141) <= 0; angryBirdLarge(8, 142) <= 0; angryBirdLarge(8, 143) <= 0; angryBirdLarge(8, 144) <= 0; angryBirdLarge(8, 145) <= 0; angryBirdLarge(8, 146) <= 0; angryBirdLarge(8, 147) <= 0; angryBirdLarge(8, 148) <= 0; angryBirdLarge(8, 149) <= 0; 
angryBirdLarge(9, 0) <= 0; angryBirdLarge(9, 1) <= 0; angryBirdLarge(9, 2) <= 0; angryBirdLarge(9, 3) <= 0; angryBirdLarge(9, 4) <= 0; angryBirdLarge(9, 5) <= 0; angryBirdLarge(9, 6) <= 0; angryBirdLarge(9, 7) <= 0; angryBirdLarge(9, 8) <= 0; angryBirdLarge(9, 9) <= 0; angryBirdLarge(9, 10) <= 0; angryBirdLarge(9, 11) <= 0; angryBirdLarge(9, 12) <= 0; angryBirdLarge(9, 13) <= 0; angryBirdLarge(9, 14) <= 0; angryBirdLarge(9, 15) <= 0; angryBirdLarge(9, 16) <= 0; angryBirdLarge(9, 17) <= 0; angryBirdLarge(9, 18) <= 0; angryBirdLarge(9, 19) <= 0; angryBirdLarge(9, 20) <= 0; angryBirdLarge(9, 21) <= 0; angryBirdLarge(9, 22) <= 0; angryBirdLarge(9, 23) <= 0; angryBirdLarge(9, 24) <= 0; angryBirdLarge(9, 25) <= 0; angryBirdLarge(9, 26) <= 0; angryBirdLarge(9, 27) <= 0; angryBirdLarge(9, 28) <= 0; angryBirdLarge(9, 29) <= 0; angryBirdLarge(9, 30) <= 0; angryBirdLarge(9, 31) <= 0; angryBirdLarge(9, 32) <= 0; angryBirdLarge(9, 33) <= 0; angryBirdLarge(9, 34) <= 0; angryBirdLarge(9, 35) <= 0; angryBirdLarge(9, 36) <= 0; angryBirdLarge(9, 37) <= 0; angryBirdLarge(9, 38) <= 0; angryBirdLarge(9, 39) <= 0; angryBirdLarge(9, 40) <= 0; angryBirdLarge(9, 41) <= 0; angryBirdLarge(9, 42) <= 0; angryBirdLarge(9, 43) <= 0; angryBirdLarge(9, 44) <= 0; angryBirdLarge(9, 45) <= 0; angryBirdLarge(9, 46) <= 0; angryBirdLarge(9, 47) <= 0; angryBirdLarge(9, 48) <= 0; angryBirdLarge(9, 49) <= 0; angryBirdLarge(9, 50) <= 0; angryBirdLarge(9, 51) <= 0; angryBirdLarge(9, 52) <= 0; angryBirdLarge(9, 53) <= 0; angryBirdLarge(9, 54) <= 0; angryBirdLarge(9, 55) <= 0; angryBirdLarge(9, 56) <= 0; angryBirdLarge(9, 57) <= 0; angryBirdLarge(9, 58) <= 0; angryBirdLarge(9, 59) <= 0; angryBirdLarge(9, 60) <= 0; angryBirdLarge(9, 61) <= 0; angryBirdLarge(9, 62) <= 0; angryBirdLarge(9, 63) <= 0; angryBirdLarge(9, 64) <= 0; angryBirdLarge(9, 65) <= 0; angryBirdLarge(9, 66) <= 5; angryBirdLarge(9, 67) <= 5; angryBirdLarge(9, 68) <= 5; angryBirdLarge(9, 69) <= 5; angryBirdLarge(9, 70) <= 5; angryBirdLarge(9, 71) <= 5; angryBirdLarge(9, 72) <= 4; angryBirdLarge(9, 73) <= 4; angryBirdLarge(9, 74) <= 4; angryBirdLarge(9, 75) <= 4; angryBirdLarge(9, 76) <= 4; angryBirdLarge(9, 77) <= 4; angryBirdLarge(9, 78) <= 4; angryBirdLarge(9, 79) <= 4; angryBirdLarge(9, 80) <= 4; angryBirdLarge(9, 81) <= 4; angryBirdLarge(9, 82) <= 4; angryBirdLarge(9, 83) <= 4; angryBirdLarge(9, 84) <= 4; angryBirdLarge(9, 85) <= 4; angryBirdLarge(9, 86) <= 4; angryBirdLarge(9, 87) <= 4; angryBirdLarge(9, 88) <= 4; angryBirdLarge(9, 89) <= 4; angryBirdLarge(9, 90) <= 5; angryBirdLarge(9, 91) <= 5; angryBirdLarge(9, 92) <= 5; angryBirdLarge(9, 93) <= 5; angryBirdLarge(9, 94) <= 5; angryBirdLarge(9, 95) <= 5; angryBirdLarge(9, 96) <= 0; angryBirdLarge(9, 97) <= 0; angryBirdLarge(9, 98) <= 0; angryBirdLarge(9, 99) <= 0; angryBirdLarge(9, 100) <= 0; angryBirdLarge(9, 101) <= 0; angryBirdLarge(9, 102) <= 0; angryBirdLarge(9, 103) <= 0; angryBirdLarge(9, 104) <= 0; angryBirdLarge(9, 105) <= 0; angryBirdLarge(9, 106) <= 0; angryBirdLarge(9, 107) <= 0; angryBirdLarge(9, 108) <= 0; angryBirdLarge(9, 109) <= 0; angryBirdLarge(9, 110) <= 0; angryBirdLarge(9, 111) <= 0; angryBirdLarge(9, 112) <= 0; angryBirdLarge(9, 113) <= 0; angryBirdLarge(9, 114) <= 0; angryBirdLarge(9, 115) <= 0; angryBirdLarge(9, 116) <= 0; angryBirdLarge(9, 117) <= 0; angryBirdLarge(9, 118) <= 0; angryBirdLarge(9, 119) <= 0; angryBirdLarge(9, 120) <= 0; angryBirdLarge(9, 121) <= 0; angryBirdLarge(9, 122) <= 0; angryBirdLarge(9, 123) <= 0; angryBirdLarge(9, 124) <= 0; angryBirdLarge(9, 125) <= 0; angryBirdLarge(9, 126) <= 0; angryBirdLarge(9, 127) <= 0; angryBirdLarge(9, 128) <= 0; angryBirdLarge(9, 129) <= 0; angryBirdLarge(9, 130) <= 0; angryBirdLarge(9, 131) <= 0; angryBirdLarge(9, 132) <= 0; angryBirdLarge(9, 133) <= 0; angryBirdLarge(9, 134) <= 0; angryBirdLarge(9, 135) <= 0; angryBirdLarge(9, 136) <= 0; angryBirdLarge(9, 137) <= 0; angryBirdLarge(9, 138) <= 0; angryBirdLarge(9, 139) <= 0; angryBirdLarge(9, 140) <= 0; angryBirdLarge(9, 141) <= 0; angryBirdLarge(9, 142) <= 0; angryBirdLarge(9, 143) <= 0; angryBirdLarge(9, 144) <= 0; angryBirdLarge(9, 145) <= 0; angryBirdLarge(9, 146) <= 0; angryBirdLarge(9, 147) <= 0; angryBirdLarge(9, 148) <= 0; angryBirdLarge(9, 149) <= 0; 
angryBirdLarge(10, 0) <= 0; angryBirdLarge(10, 1) <= 0; angryBirdLarge(10, 2) <= 0; angryBirdLarge(10, 3) <= 0; angryBirdLarge(10, 4) <= 0; angryBirdLarge(10, 5) <= 0; angryBirdLarge(10, 6) <= 0; angryBirdLarge(10, 7) <= 0; angryBirdLarge(10, 8) <= 0; angryBirdLarge(10, 9) <= 0; angryBirdLarge(10, 10) <= 0; angryBirdLarge(10, 11) <= 0; angryBirdLarge(10, 12) <= 0; angryBirdLarge(10, 13) <= 0; angryBirdLarge(10, 14) <= 0; angryBirdLarge(10, 15) <= 0; angryBirdLarge(10, 16) <= 0; angryBirdLarge(10, 17) <= 0; angryBirdLarge(10, 18) <= 0; angryBirdLarge(10, 19) <= 0; angryBirdLarge(10, 20) <= 0; angryBirdLarge(10, 21) <= 0; angryBirdLarge(10, 22) <= 0; angryBirdLarge(10, 23) <= 0; angryBirdLarge(10, 24) <= 0; angryBirdLarge(10, 25) <= 0; angryBirdLarge(10, 26) <= 0; angryBirdLarge(10, 27) <= 0; angryBirdLarge(10, 28) <= 0; angryBirdLarge(10, 29) <= 0; angryBirdLarge(10, 30) <= 0; angryBirdLarge(10, 31) <= 0; angryBirdLarge(10, 32) <= 0; angryBirdLarge(10, 33) <= 0; angryBirdLarge(10, 34) <= 0; angryBirdLarge(10, 35) <= 0; angryBirdLarge(10, 36) <= 0; angryBirdLarge(10, 37) <= 0; angryBirdLarge(10, 38) <= 0; angryBirdLarge(10, 39) <= 0; angryBirdLarge(10, 40) <= 0; angryBirdLarge(10, 41) <= 0; angryBirdLarge(10, 42) <= 0; angryBirdLarge(10, 43) <= 0; angryBirdLarge(10, 44) <= 0; angryBirdLarge(10, 45) <= 0; angryBirdLarge(10, 46) <= 0; angryBirdLarge(10, 47) <= 0; angryBirdLarge(10, 48) <= 0; angryBirdLarge(10, 49) <= 0; angryBirdLarge(10, 50) <= 0; angryBirdLarge(10, 51) <= 0; angryBirdLarge(10, 52) <= 0; angryBirdLarge(10, 53) <= 0; angryBirdLarge(10, 54) <= 0; angryBirdLarge(10, 55) <= 0; angryBirdLarge(10, 56) <= 0; angryBirdLarge(10, 57) <= 0; angryBirdLarge(10, 58) <= 0; angryBirdLarge(10, 59) <= 0; angryBirdLarge(10, 60) <= 0; angryBirdLarge(10, 61) <= 0; angryBirdLarge(10, 62) <= 0; angryBirdLarge(10, 63) <= 0; angryBirdLarge(10, 64) <= 0; angryBirdLarge(10, 65) <= 0; angryBirdLarge(10, 66) <= 5; angryBirdLarge(10, 67) <= 5; angryBirdLarge(10, 68) <= 5; angryBirdLarge(10, 69) <= 5; angryBirdLarge(10, 70) <= 5; angryBirdLarge(10, 71) <= 5; angryBirdLarge(10, 72) <= 4; angryBirdLarge(10, 73) <= 4; angryBirdLarge(10, 74) <= 4; angryBirdLarge(10, 75) <= 4; angryBirdLarge(10, 76) <= 4; angryBirdLarge(10, 77) <= 4; angryBirdLarge(10, 78) <= 4; angryBirdLarge(10, 79) <= 4; angryBirdLarge(10, 80) <= 4; angryBirdLarge(10, 81) <= 4; angryBirdLarge(10, 82) <= 4; angryBirdLarge(10, 83) <= 4; angryBirdLarge(10, 84) <= 4; angryBirdLarge(10, 85) <= 4; angryBirdLarge(10, 86) <= 4; angryBirdLarge(10, 87) <= 4; angryBirdLarge(10, 88) <= 4; angryBirdLarge(10, 89) <= 4; angryBirdLarge(10, 90) <= 5; angryBirdLarge(10, 91) <= 5; angryBirdLarge(10, 92) <= 5; angryBirdLarge(10, 93) <= 5; angryBirdLarge(10, 94) <= 5; angryBirdLarge(10, 95) <= 5; angryBirdLarge(10, 96) <= 0; angryBirdLarge(10, 97) <= 0; angryBirdLarge(10, 98) <= 0; angryBirdLarge(10, 99) <= 0; angryBirdLarge(10, 100) <= 0; angryBirdLarge(10, 101) <= 0; angryBirdLarge(10, 102) <= 0; angryBirdLarge(10, 103) <= 0; angryBirdLarge(10, 104) <= 0; angryBirdLarge(10, 105) <= 0; angryBirdLarge(10, 106) <= 0; angryBirdLarge(10, 107) <= 0; angryBirdLarge(10, 108) <= 0; angryBirdLarge(10, 109) <= 0; angryBirdLarge(10, 110) <= 0; angryBirdLarge(10, 111) <= 0; angryBirdLarge(10, 112) <= 0; angryBirdLarge(10, 113) <= 0; angryBirdLarge(10, 114) <= 0; angryBirdLarge(10, 115) <= 0; angryBirdLarge(10, 116) <= 0; angryBirdLarge(10, 117) <= 0; angryBirdLarge(10, 118) <= 0; angryBirdLarge(10, 119) <= 0; angryBirdLarge(10, 120) <= 0; angryBirdLarge(10, 121) <= 0; angryBirdLarge(10, 122) <= 0; angryBirdLarge(10, 123) <= 0; angryBirdLarge(10, 124) <= 0; angryBirdLarge(10, 125) <= 0; angryBirdLarge(10, 126) <= 0; angryBirdLarge(10, 127) <= 0; angryBirdLarge(10, 128) <= 0; angryBirdLarge(10, 129) <= 0; angryBirdLarge(10, 130) <= 0; angryBirdLarge(10, 131) <= 0; angryBirdLarge(10, 132) <= 0; angryBirdLarge(10, 133) <= 0; angryBirdLarge(10, 134) <= 0; angryBirdLarge(10, 135) <= 0; angryBirdLarge(10, 136) <= 0; angryBirdLarge(10, 137) <= 0; angryBirdLarge(10, 138) <= 0; angryBirdLarge(10, 139) <= 0; angryBirdLarge(10, 140) <= 0; angryBirdLarge(10, 141) <= 0; angryBirdLarge(10, 142) <= 0; angryBirdLarge(10, 143) <= 0; angryBirdLarge(10, 144) <= 0; angryBirdLarge(10, 145) <= 0; angryBirdLarge(10, 146) <= 0; angryBirdLarge(10, 147) <= 0; angryBirdLarge(10, 148) <= 0; angryBirdLarge(10, 149) <= 0; 
angryBirdLarge(11, 0) <= 0; angryBirdLarge(11, 1) <= 0; angryBirdLarge(11, 2) <= 0; angryBirdLarge(11, 3) <= 0; angryBirdLarge(11, 4) <= 0; angryBirdLarge(11, 5) <= 0; angryBirdLarge(11, 6) <= 0; angryBirdLarge(11, 7) <= 0; angryBirdLarge(11, 8) <= 0; angryBirdLarge(11, 9) <= 0; angryBirdLarge(11, 10) <= 0; angryBirdLarge(11, 11) <= 0; angryBirdLarge(11, 12) <= 0; angryBirdLarge(11, 13) <= 0; angryBirdLarge(11, 14) <= 0; angryBirdLarge(11, 15) <= 0; angryBirdLarge(11, 16) <= 0; angryBirdLarge(11, 17) <= 0; angryBirdLarge(11, 18) <= 0; angryBirdLarge(11, 19) <= 0; angryBirdLarge(11, 20) <= 0; angryBirdLarge(11, 21) <= 0; angryBirdLarge(11, 22) <= 0; angryBirdLarge(11, 23) <= 0; angryBirdLarge(11, 24) <= 0; angryBirdLarge(11, 25) <= 0; angryBirdLarge(11, 26) <= 0; angryBirdLarge(11, 27) <= 0; angryBirdLarge(11, 28) <= 0; angryBirdLarge(11, 29) <= 0; angryBirdLarge(11, 30) <= 0; angryBirdLarge(11, 31) <= 0; angryBirdLarge(11, 32) <= 0; angryBirdLarge(11, 33) <= 0; angryBirdLarge(11, 34) <= 0; angryBirdLarge(11, 35) <= 0; angryBirdLarge(11, 36) <= 0; angryBirdLarge(11, 37) <= 0; angryBirdLarge(11, 38) <= 0; angryBirdLarge(11, 39) <= 0; angryBirdLarge(11, 40) <= 0; angryBirdLarge(11, 41) <= 0; angryBirdLarge(11, 42) <= 0; angryBirdLarge(11, 43) <= 0; angryBirdLarge(11, 44) <= 0; angryBirdLarge(11, 45) <= 0; angryBirdLarge(11, 46) <= 0; angryBirdLarge(11, 47) <= 0; angryBirdLarge(11, 48) <= 0; angryBirdLarge(11, 49) <= 0; angryBirdLarge(11, 50) <= 0; angryBirdLarge(11, 51) <= 0; angryBirdLarge(11, 52) <= 0; angryBirdLarge(11, 53) <= 0; angryBirdLarge(11, 54) <= 0; angryBirdLarge(11, 55) <= 0; angryBirdLarge(11, 56) <= 0; angryBirdLarge(11, 57) <= 0; angryBirdLarge(11, 58) <= 0; angryBirdLarge(11, 59) <= 0; angryBirdLarge(11, 60) <= 0; angryBirdLarge(11, 61) <= 0; angryBirdLarge(11, 62) <= 0; angryBirdLarge(11, 63) <= 0; angryBirdLarge(11, 64) <= 0; angryBirdLarge(11, 65) <= 0; angryBirdLarge(11, 66) <= 5; angryBirdLarge(11, 67) <= 5; angryBirdLarge(11, 68) <= 5; angryBirdLarge(11, 69) <= 5; angryBirdLarge(11, 70) <= 5; angryBirdLarge(11, 71) <= 5; angryBirdLarge(11, 72) <= 4; angryBirdLarge(11, 73) <= 4; angryBirdLarge(11, 74) <= 4; angryBirdLarge(11, 75) <= 4; angryBirdLarge(11, 76) <= 4; angryBirdLarge(11, 77) <= 4; angryBirdLarge(11, 78) <= 4; angryBirdLarge(11, 79) <= 4; angryBirdLarge(11, 80) <= 4; angryBirdLarge(11, 81) <= 4; angryBirdLarge(11, 82) <= 4; angryBirdLarge(11, 83) <= 4; angryBirdLarge(11, 84) <= 4; angryBirdLarge(11, 85) <= 4; angryBirdLarge(11, 86) <= 4; angryBirdLarge(11, 87) <= 4; angryBirdLarge(11, 88) <= 4; angryBirdLarge(11, 89) <= 4; angryBirdLarge(11, 90) <= 5; angryBirdLarge(11, 91) <= 5; angryBirdLarge(11, 92) <= 5; angryBirdLarge(11, 93) <= 5; angryBirdLarge(11, 94) <= 5; angryBirdLarge(11, 95) <= 5; angryBirdLarge(11, 96) <= 0; angryBirdLarge(11, 97) <= 0; angryBirdLarge(11, 98) <= 0; angryBirdLarge(11, 99) <= 0; angryBirdLarge(11, 100) <= 0; angryBirdLarge(11, 101) <= 0; angryBirdLarge(11, 102) <= 0; angryBirdLarge(11, 103) <= 0; angryBirdLarge(11, 104) <= 0; angryBirdLarge(11, 105) <= 0; angryBirdLarge(11, 106) <= 0; angryBirdLarge(11, 107) <= 0; angryBirdLarge(11, 108) <= 0; angryBirdLarge(11, 109) <= 0; angryBirdLarge(11, 110) <= 0; angryBirdLarge(11, 111) <= 0; angryBirdLarge(11, 112) <= 0; angryBirdLarge(11, 113) <= 0; angryBirdLarge(11, 114) <= 0; angryBirdLarge(11, 115) <= 0; angryBirdLarge(11, 116) <= 0; angryBirdLarge(11, 117) <= 0; angryBirdLarge(11, 118) <= 0; angryBirdLarge(11, 119) <= 0; angryBirdLarge(11, 120) <= 0; angryBirdLarge(11, 121) <= 0; angryBirdLarge(11, 122) <= 0; angryBirdLarge(11, 123) <= 0; angryBirdLarge(11, 124) <= 0; angryBirdLarge(11, 125) <= 0; angryBirdLarge(11, 126) <= 0; angryBirdLarge(11, 127) <= 0; angryBirdLarge(11, 128) <= 0; angryBirdLarge(11, 129) <= 0; angryBirdLarge(11, 130) <= 0; angryBirdLarge(11, 131) <= 0; angryBirdLarge(11, 132) <= 0; angryBirdLarge(11, 133) <= 0; angryBirdLarge(11, 134) <= 0; angryBirdLarge(11, 135) <= 0; angryBirdLarge(11, 136) <= 0; angryBirdLarge(11, 137) <= 0; angryBirdLarge(11, 138) <= 0; angryBirdLarge(11, 139) <= 0; angryBirdLarge(11, 140) <= 0; angryBirdLarge(11, 141) <= 0; angryBirdLarge(11, 142) <= 0; angryBirdLarge(11, 143) <= 0; angryBirdLarge(11, 144) <= 0; angryBirdLarge(11, 145) <= 0; angryBirdLarge(11, 146) <= 0; angryBirdLarge(11, 147) <= 0; angryBirdLarge(11, 148) <= 0; angryBirdLarge(11, 149) <= 0; 
angryBirdLarge(12, 0) <= 0; angryBirdLarge(12, 1) <= 0; angryBirdLarge(12, 2) <= 0; angryBirdLarge(12, 3) <= 0; angryBirdLarge(12, 4) <= 0; angryBirdLarge(12, 5) <= 0; angryBirdLarge(12, 6) <= 0; angryBirdLarge(12, 7) <= 0; angryBirdLarge(12, 8) <= 0; angryBirdLarge(12, 9) <= 0; angryBirdLarge(12, 10) <= 0; angryBirdLarge(12, 11) <= 0; angryBirdLarge(12, 12) <= 0; angryBirdLarge(12, 13) <= 0; angryBirdLarge(12, 14) <= 0; angryBirdLarge(12, 15) <= 0; angryBirdLarge(12, 16) <= 0; angryBirdLarge(12, 17) <= 0; angryBirdLarge(12, 18) <= 0; angryBirdLarge(12, 19) <= 0; angryBirdLarge(12, 20) <= 0; angryBirdLarge(12, 21) <= 0; angryBirdLarge(12, 22) <= 0; angryBirdLarge(12, 23) <= 0; angryBirdLarge(12, 24) <= 0; angryBirdLarge(12, 25) <= 0; angryBirdLarge(12, 26) <= 0; angryBirdLarge(12, 27) <= 0; angryBirdLarge(12, 28) <= 0; angryBirdLarge(12, 29) <= 0; angryBirdLarge(12, 30) <= 0; angryBirdLarge(12, 31) <= 0; angryBirdLarge(12, 32) <= 0; angryBirdLarge(12, 33) <= 0; angryBirdLarge(12, 34) <= 0; angryBirdLarge(12, 35) <= 0; angryBirdLarge(12, 36) <= 0; angryBirdLarge(12, 37) <= 0; angryBirdLarge(12, 38) <= 0; angryBirdLarge(12, 39) <= 0; angryBirdLarge(12, 40) <= 0; angryBirdLarge(12, 41) <= 0; angryBirdLarge(12, 42) <= 0; angryBirdLarge(12, 43) <= 0; angryBirdLarge(12, 44) <= 0; angryBirdLarge(12, 45) <= 0; angryBirdLarge(12, 46) <= 0; angryBirdLarge(12, 47) <= 0; angryBirdLarge(12, 48) <= 5; angryBirdLarge(12, 49) <= 5; angryBirdLarge(12, 50) <= 5; angryBirdLarge(12, 51) <= 5; angryBirdLarge(12, 52) <= 5; angryBirdLarge(12, 53) <= 5; angryBirdLarge(12, 54) <= 5; angryBirdLarge(12, 55) <= 5; angryBirdLarge(12, 56) <= 5; angryBirdLarge(12, 57) <= 5; angryBirdLarge(12, 58) <= 5; angryBirdLarge(12, 59) <= 5; angryBirdLarge(12, 60) <= 5; angryBirdLarge(12, 61) <= 5; angryBirdLarge(12, 62) <= 5; angryBirdLarge(12, 63) <= 5; angryBirdLarge(12, 64) <= 5; angryBirdLarge(12, 65) <= 5; angryBirdLarge(12, 66) <= 5; angryBirdLarge(12, 67) <= 5; angryBirdLarge(12, 68) <= 5; angryBirdLarge(12, 69) <= 5; angryBirdLarge(12, 70) <= 5; angryBirdLarge(12, 71) <= 5; angryBirdLarge(12, 72) <= 4; angryBirdLarge(12, 73) <= 4; angryBirdLarge(12, 74) <= 4; angryBirdLarge(12, 75) <= 4; angryBirdLarge(12, 76) <= 4; angryBirdLarge(12, 77) <= 4; angryBirdLarge(12, 78) <= 4; angryBirdLarge(12, 79) <= 4; angryBirdLarge(12, 80) <= 4; angryBirdLarge(12, 81) <= 4; angryBirdLarge(12, 82) <= 4; angryBirdLarge(12, 83) <= 4; angryBirdLarge(12, 84) <= 4; angryBirdLarge(12, 85) <= 4; angryBirdLarge(12, 86) <= 4; angryBirdLarge(12, 87) <= 4; angryBirdLarge(12, 88) <= 4; angryBirdLarge(12, 89) <= 4; angryBirdLarge(12, 90) <= 4; angryBirdLarge(12, 91) <= 4; angryBirdLarge(12, 92) <= 4; angryBirdLarge(12, 93) <= 4; angryBirdLarge(12, 94) <= 4; angryBirdLarge(12, 95) <= 4; angryBirdLarge(12, 96) <= 5; angryBirdLarge(12, 97) <= 5; angryBirdLarge(12, 98) <= 5; angryBirdLarge(12, 99) <= 5; angryBirdLarge(12, 100) <= 5; angryBirdLarge(12, 101) <= 5; angryBirdLarge(12, 102) <= 0; angryBirdLarge(12, 103) <= 0; angryBirdLarge(12, 104) <= 0; angryBirdLarge(12, 105) <= 0; angryBirdLarge(12, 106) <= 0; angryBirdLarge(12, 107) <= 0; angryBirdLarge(12, 108) <= 0; angryBirdLarge(12, 109) <= 0; angryBirdLarge(12, 110) <= 0; angryBirdLarge(12, 111) <= 0; angryBirdLarge(12, 112) <= 0; angryBirdLarge(12, 113) <= 0; angryBirdLarge(12, 114) <= 0; angryBirdLarge(12, 115) <= 0; angryBirdLarge(12, 116) <= 0; angryBirdLarge(12, 117) <= 0; angryBirdLarge(12, 118) <= 0; angryBirdLarge(12, 119) <= 0; angryBirdLarge(12, 120) <= 0; angryBirdLarge(12, 121) <= 0; angryBirdLarge(12, 122) <= 0; angryBirdLarge(12, 123) <= 0; angryBirdLarge(12, 124) <= 0; angryBirdLarge(12, 125) <= 0; angryBirdLarge(12, 126) <= 0; angryBirdLarge(12, 127) <= 0; angryBirdLarge(12, 128) <= 0; angryBirdLarge(12, 129) <= 0; angryBirdLarge(12, 130) <= 0; angryBirdLarge(12, 131) <= 0; angryBirdLarge(12, 132) <= 0; angryBirdLarge(12, 133) <= 0; angryBirdLarge(12, 134) <= 0; angryBirdLarge(12, 135) <= 0; angryBirdLarge(12, 136) <= 0; angryBirdLarge(12, 137) <= 0; angryBirdLarge(12, 138) <= 0; angryBirdLarge(12, 139) <= 0; angryBirdLarge(12, 140) <= 0; angryBirdLarge(12, 141) <= 0; angryBirdLarge(12, 142) <= 0; angryBirdLarge(12, 143) <= 0; angryBirdLarge(12, 144) <= 0; angryBirdLarge(12, 145) <= 0; angryBirdLarge(12, 146) <= 0; angryBirdLarge(12, 147) <= 0; angryBirdLarge(12, 148) <= 0; angryBirdLarge(12, 149) <= 0; 
angryBirdLarge(13, 0) <= 0; angryBirdLarge(13, 1) <= 0; angryBirdLarge(13, 2) <= 0; angryBirdLarge(13, 3) <= 0; angryBirdLarge(13, 4) <= 0; angryBirdLarge(13, 5) <= 0; angryBirdLarge(13, 6) <= 0; angryBirdLarge(13, 7) <= 0; angryBirdLarge(13, 8) <= 0; angryBirdLarge(13, 9) <= 0; angryBirdLarge(13, 10) <= 0; angryBirdLarge(13, 11) <= 0; angryBirdLarge(13, 12) <= 0; angryBirdLarge(13, 13) <= 0; angryBirdLarge(13, 14) <= 0; angryBirdLarge(13, 15) <= 0; angryBirdLarge(13, 16) <= 0; angryBirdLarge(13, 17) <= 0; angryBirdLarge(13, 18) <= 0; angryBirdLarge(13, 19) <= 0; angryBirdLarge(13, 20) <= 0; angryBirdLarge(13, 21) <= 0; angryBirdLarge(13, 22) <= 0; angryBirdLarge(13, 23) <= 0; angryBirdLarge(13, 24) <= 0; angryBirdLarge(13, 25) <= 0; angryBirdLarge(13, 26) <= 0; angryBirdLarge(13, 27) <= 0; angryBirdLarge(13, 28) <= 0; angryBirdLarge(13, 29) <= 0; angryBirdLarge(13, 30) <= 0; angryBirdLarge(13, 31) <= 0; angryBirdLarge(13, 32) <= 0; angryBirdLarge(13, 33) <= 0; angryBirdLarge(13, 34) <= 0; angryBirdLarge(13, 35) <= 0; angryBirdLarge(13, 36) <= 0; angryBirdLarge(13, 37) <= 0; angryBirdLarge(13, 38) <= 0; angryBirdLarge(13, 39) <= 0; angryBirdLarge(13, 40) <= 0; angryBirdLarge(13, 41) <= 0; angryBirdLarge(13, 42) <= 0; angryBirdLarge(13, 43) <= 0; angryBirdLarge(13, 44) <= 0; angryBirdLarge(13, 45) <= 0; angryBirdLarge(13, 46) <= 0; angryBirdLarge(13, 47) <= 0; angryBirdLarge(13, 48) <= 5; angryBirdLarge(13, 49) <= 5; angryBirdLarge(13, 50) <= 5; angryBirdLarge(13, 51) <= 5; angryBirdLarge(13, 52) <= 5; angryBirdLarge(13, 53) <= 5; angryBirdLarge(13, 54) <= 5; angryBirdLarge(13, 55) <= 5; angryBirdLarge(13, 56) <= 5; angryBirdLarge(13, 57) <= 5; angryBirdLarge(13, 58) <= 5; angryBirdLarge(13, 59) <= 5; angryBirdLarge(13, 60) <= 5; angryBirdLarge(13, 61) <= 5; angryBirdLarge(13, 62) <= 5; angryBirdLarge(13, 63) <= 5; angryBirdLarge(13, 64) <= 5; angryBirdLarge(13, 65) <= 5; angryBirdLarge(13, 66) <= 5; angryBirdLarge(13, 67) <= 5; angryBirdLarge(13, 68) <= 5; angryBirdLarge(13, 69) <= 5; angryBirdLarge(13, 70) <= 5; angryBirdLarge(13, 71) <= 5; angryBirdLarge(13, 72) <= 4; angryBirdLarge(13, 73) <= 4; angryBirdLarge(13, 74) <= 4; angryBirdLarge(13, 75) <= 4; angryBirdLarge(13, 76) <= 4; angryBirdLarge(13, 77) <= 4; angryBirdLarge(13, 78) <= 4; angryBirdLarge(13, 79) <= 4; angryBirdLarge(13, 80) <= 4; angryBirdLarge(13, 81) <= 4; angryBirdLarge(13, 82) <= 4; angryBirdLarge(13, 83) <= 4; angryBirdLarge(13, 84) <= 4; angryBirdLarge(13, 85) <= 4; angryBirdLarge(13, 86) <= 4; angryBirdLarge(13, 87) <= 4; angryBirdLarge(13, 88) <= 4; angryBirdLarge(13, 89) <= 4; angryBirdLarge(13, 90) <= 4; angryBirdLarge(13, 91) <= 4; angryBirdLarge(13, 92) <= 4; angryBirdLarge(13, 93) <= 4; angryBirdLarge(13, 94) <= 4; angryBirdLarge(13, 95) <= 4; angryBirdLarge(13, 96) <= 5; angryBirdLarge(13, 97) <= 5; angryBirdLarge(13, 98) <= 5; angryBirdLarge(13, 99) <= 5; angryBirdLarge(13, 100) <= 5; angryBirdLarge(13, 101) <= 5; angryBirdLarge(13, 102) <= 0; angryBirdLarge(13, 103) <= 0; angryBirdLarge(13, 104) <= 0; angryBirdLarge(13, 105) <= 0; angryBirdLarge(13, 106) <= 0; angryBirdLarge(13, 107) <= 0; angryBirdLarge(13, 108) <= 0; angryBirdLarge(13, 109) <= 0; angryBirdLarge(13, 110) <= 0; angryBirdLarge(13, 111) <= 0; angryBirdLarge(13, 112) <= 0; angryBirdLarge(13, 113) <= 0; angryBirdLarge(13, 114) <= 0; angryBirdLarge(13, 115) <= 0; angryBirdLarge(13, 116) <= 0; angryBirdLarge(13, 117) <= 0; angryBirdLarge(13, 118) <= 0; angryBirdLarge(13, 119) <= 0; angryBirdLarge(13, 120) <= 0; angryBirdLarge(13, 121) <= 0; angryBirdLarge(13, 122) <= 0; angryBirdLarge(13, 123) <= 0; angryBirdLarge(13, 124) <= 0; angryBirdLarge(13, 125) <= 0; angryBirdLarge(13, 126) <= 0; angryBirdLarge(13, 127) <= 0; angryBirdLarge(13, 128) <= 0; angryBirdLarge(13, 129) <= 0; angryBirdLarge(13, 130) <= 0; angryBirdLarge(13, 131) <= 0; angryBirdLarge(13, 132) <= 0; angryBirdLarge(13, 133) <= 0; angryBirdLarge(13, 134) <= 0; angryBirdLarge(13, 135) <= 0; angryBirdLarge(13, 136) <= 0; angryBirdLarge(13, 137) <= 0; angryBirdLarge(13, 138) <= 0; angryBirdLarge(13, 139) <= 0; angryBirdLarge(13, 140) <= 0; angryBirdLarge(13, 141) <= 0; angryBirdLarge(13, 142) <= 0; angryBirdLarge(13, 143) <= 0; angryBirdLarge(13, 144) <= 0; angryBirdLarge(13, 145) <= 0; angryBirdLarge(13, 146) <= 0; angryBirdLarge(13, 147) <= 0; angryBirdLarge(13, 148) <= 0; angryBirdLarge(13, 149) <= 0; 
angryBirdLarge(14, 0) <= 0; angryBirdLarge(14, 1) <= 0; angryBirdLarge(14, 2) <= 0; angryBirdLarge(14, 3) <= 0; angryBirdLarge(14, 4) <= 0; angryBirdLarge(14, 5) <= 0; angryBirdLarge(14, 6) <= 0; angryBirdLarge(14, 7) <= 0; angryBirdLarge(14, 8) <= 0; angryBirdLarge(14, 9) <= 0; angryBirdLarge(14, 10) <= 0; angryBirdLarge(14, 11) <= 0; angryBirdLarge(14, 12) <= 0; angryBirdLarge(14, 13) <= 0; angryBirdLarge(14, 14) <= 0; angryBirdLarge(14, 15) <= 0; angryBirdLarge(14, 16) <= 0; angryBirdLarge(14, 17) <= 0; angryBirdLarge(14, 18) <= 0; angryBirdLarge(14, 19) <= 0; angryBirdLarge(14, 20) <= 0; angryBirdLarge(14, 21) <= 0; angryBirdLarge(14, 22) <= 0; angryBirdLarge(14, 23) <= 0; angryBirdLarge(14, 24) <= 0; angryBirdLarge(14, 25) <= 0; angryBirdLarge(14, 26) <= 0; angryBirdLarge(14, 27) <= 0; angryBirdLarge(14, 28) <= 0; angryBirdLarge(14, 29) <= 0; angryBirdLarge(14, 30) <= 0; angryBirdLarge(14, 31) <= 0; angryBirdLarge(14, 32) <= 0; angryBirdLarge(14, 33) <= 0; angryBirdLarge(14, 34) <= 0; angryBirdLarge(14, 35) <= 0; angryBirdLarge(14, 36) <= 0; angryBirdLarge(14, 37) <= 0; angryBirdLarge(14, 38) <= 0; angryBirdLarge(14, 39) <= 0; angryBirdLarge(14, 40) <= 0; angryBirdLarge(14, 41) <= 0; angryBirdLarge(14, 42) <= 0; angryBirdLarge(14, 43) <= 0; angryBirdLarge(14, 44) <= 0; angryBirdLarge(14, 45) <= 0; angryBirdLarge(14, 46) <= 0; angryBirdLarge(14, 47) <= 0; angryBirdLarge(14, 48) <= 5; angryBirdLarge(14, 49) <= 5; angryBirdLarge(14, 50) <= 5; angryBirdLarge(14, 51) <= 5; angryBirdLarge(14, 52) <= 5; angryBirdLarge(14, 53) <= 5; angryBirdLarge(14, 54) <= 5; angryBirdLarge(14, 55) <= 5; angryBirdLarge(14, 56) <= 5; angryBirdLarge(14, 57) <= 5; angryBirdLarge(14, 58) <= 5; angryBirdLarge(14, 59) <= 5; angryBirdLarge(14, 60) <= 5; angryBirdLarge(14, 61) <= 5; angryBirdLarge(14, 62) <= 5; angryBirdLarge(14, 63) <= 5; angryBirdLarge(14, 64) <= 5; angryBirdLarge(14, 65) <= 5; angryBirdLarge(14, 66) <= 5; angryBirdLarge(14, 67) <= 5; angryBirdLarge(14, 68) <= 5; angryBirdLarge(14, 69) <= 5; angryBirdLarge(14, 70) <= 5; angryBirdLarge(14, 71) <= 5; angryBirdLarge(14, 72) <= 4; angryBirdLarge(14, 73) <= 4; angryBirdLarge(14, 74) <= 4; angryBirdLarge(14, 75) <= 4; angryBirdLarge(14, 76) <= 4; angryBirdLarge(14, 77) <= 4; angryBirdLarge(14, 78) <= 4; angryBirdLarge(14, 79) <= 4; angryBirdLarge(14, 80) <= 4; angryBirdLarge(14, 81) <= 4; angryBirdLarge(14, 82) <= 4; angryBirdLarge(14, 83) <= 4; angryBirdLarge(14, 84) <= 4; angryBirdLarge(14, 85) <= 4; angryBirdLarge(14, 86) <= 4; angryBirdLarge(14, 87) <= 4; angryBirdLarge(14, 88) <= 4; angryBirdLarge(14, 89) <= 4; angryBirdLarge(14, 90) <= 4; angryBirdLarge(14, 91) <= 4; angryBirdLarge(14, 92) <= 4; angryBirdLarge(14, 93) <= 4; angryBirdLarge(14, 94) <= 4; angryBirdLarge(14, 95) <= 4; angryBirdLarge(14, 96) <= 5; angryBirdLarge(14, 97) <= 5; angryBirdLarge(14, 98) <= 5; angryBirdLarge(14, 99) <= 5; angryBirdLarge(14, 100) <= 5; angryBirdLarge(14, 101) <= 5; angryBirdLarge(14, 102) <= 0; angryBirdLarge(14, 103) <= 0; angryBirdLarge(14, 104) <= 0; angryBirdLarge(14, 105) <= 0; angryBirdLarge(14, 106) <= 0; angryBirdLarge(14, 107) <= 0; angryBirdLarge(14, 108) <= 0; angryBirdLarge(14, 109) <= 0; angryBirdLarge(14, 110) <= 0; angryBirdLarge(14, 111) <= 0; angryBirdLarge(14, 112) <= 0; angryBirdLarge(14, 113) <= 0; angryBirdLarge(14, 114) <= 0; angryBirdLarge(14, 115) <= 0; angryBirdLarge(14, 116) <= 0; angryBirdLarge(14, 117) <= 0; angryBirdLarge(14, 118) <= 0; angryBirdLarge(14, 119) <= 0; angryBirdLarge(14, 120) <= 0; angryBirdLarge(14, 121) <= 0; angryBirdLarge(14, 122) <= 0; angryBirdLarge(14, 123) <= 0; angryBirdLarge(14, 124) <= 0; angryBirdLarge(14, 125) <= 0; angryBirdLarge(14, 126) <= 0; angryBirdLarge(14, 127) <= 0; angryBirdLarge(14, 128) <= 0; angryBirdLarge(14, 129) <= 0; angryBirdLarge(14, 130) <= 0; angryBirdLarge(14, 131) <= 0; angryBirdLarge(14, 132) <= 0; angryBirdLarge(14, 133) <= 0; angryBirdLarge(14, 134) <= 0; angryBirdLarge(14, 135) <= 0; angryBirdLarge(14, 136) <= 0; angryBirdLarge(14, 137) <= 0; angryBirdLarge(14, 138) <= 0; angryBirdLarge(14, 139) <= 0; angryBirdLarge(14, 140) <= 0; angryBirdLarge(14, 141) <= 0; angryBirdLarge(14, 142) <= 0; angryBirdLarge(14, 143) <= 0; angryBirdLarge(14, 144) <= 0; angryBirdLarge(14, 145) <= 0; angryBirdLarge(14, 146) <= 0; angryBirdLarge(14, 147) <= 0; angryBirdLarge(14, 148) <= 0; angryBirdLarge(14, 149) <= 0; 
angryBirdLarge(15, 0) <= 0; angryBirdLarge(15, 1) <= 0; angryBirdLarge(15, 2) <= 0; angryBirdLarge(15, 3) <= 0; angryBirdLarge(15, 4) <= 0; angryBirdLarge(15, 5) <= 0; angryBirdLarge(15, 6) <= 0; angryBirdLarge(15, 7) <= 0; angryBirdLarge(15, 8) <= 0; angryBirdLarge(15, 9) <= 0; angryBirdLarge(15, 10) <= 0; angryBirdLarge(15, 11) <= 0; angryBirdLarge(15, 12) <= 0; angryBirdLarge(15, 13) <= 0; angryBirdLarge(15, 14) <= 0; angryBirdLarge(15, 15) <= 0; angryBirdLarge(15, 16) <= 0; angryBirdLarge(15, 17) <= 0; angryBirdLarge(15, 18) <= 0; angryBirdLarge(15, 19) <= 0; angryBirdLarge(15, 20) <= 0; angryBirdLarge(15, 21) <= 0; angryBirdLarge(15, 22) <= 0; angryBirdLarge(15, 23) <= 0; angryBirdLarge(15, 24) <= 0; angryBirdLarge(15, 25) <= 0; angryBirdLarge(15, 26) <= 0; angryBirdLarge(15, 27) <= 0; angryBirdLarge(15, 28) <= 0; angryBirdLarge(15, 29) <= 0; angryBirdLarge(15, 30) <= 0; angryBirdLarge(15, 31) <= 0; angryBirdLarge(15, 32) <= 0; angryBirdLarge(15, 33) <= 0; angryBirdLarge(15, 34) <= 0; angryBirdLarge(15, 35) <= 0; angryBirdLarge(15, 36) <= 0; angryBirdLarge(15, 37) <= 0; angryBirdLarge(15, 38) <= 0; angryBirdLarge(15, 39) <= 0; angryBirdLarge(15, 40) <= 0; angryBirdLarge(15, 41) <= 0; angryBirdLarge(15, 42) <= 0; angryBirdLarge(15, 43) <= 0; angryBirdLarge(15, 44) <= 0; angryBirdLarge(15, 45) <= 0; angryBirdLarge(15, 46) <= 0; angryBirdLarge(15, 47) <= 0; angryBirdLarge(15, 48) <= 5; angryBirdLarge(15, 49) <= 5; angryBirdLarge(15, 50) <= 5; angryBirdLarge(15, 51) <= 5; angryBirdLarge(15, 52) <= 5; angryBirdLarge(15, 53) <= 5; angryBirdLarge(15, 54) <= 5; angryBirdLarge(15, 55) <= 5; angryBirdLarge(15, 56) <= 5; angryBirdLarge(15, 57) <= 5; angryBirdLarge(15, 58) <= 5; angryBirdLarge(15, 59) <= 5; angryBirdLarge(15, 60) <= 5; angryBirdLarge(15, 61) <= 5; angryBirdLarge(15, 62) <= 5; angryBirdLarge(15, 63) <= 5; angryBirdLarge(15, 64) <= 5; angryBirdLarge(15, 65) <= 5; angryBirdLarge(15, 66) <= 5; angryBirdLarge(15, 67) <= 5; angryBirdLarge(15, 68) <= 5; angryBirdLarge(15, 69) <= 5; angryBirdLarge(15, 70) <= 5; angryBirdLarge(15, 71) <= 5; angryBirdLarge(15, 72) <= 4; angryBirdLarge(15, 73) <= 4; angryBirdLarge(15, 74) <= 4; angryBirdLarge(15, 75) <= 4; angryBirdLarge(15, 76) <= 4; angryBirdLarge(15, 77) <= 4; angryBirdLarge(15, 78) <= 4; angryBirdLarge(15, 79) <= 4; angryBirdLarge(15, 80) <= 4; angryBirdLarge(15, 81) <= 4; angryBirdLarge(15, 82) <= 4; angryBirdLarge(15, 83) <= 4; angryBirdLarge(15, 84) <= 4; angryBirdLarge(15, 85) <= 4; angryBirdLarge(15, 86) <= 4; angryBirdLarge(15, 87) <= 4; angryBirdLarge(15, 88) <= 4; angryBirdLarge(15, 89) <= 4; angryBirdLarge(15, 90) <= 4; angryBirdLarge(15, 91) <= 4; angryBirdLarge(15, 92) <= 4; angryBirdLarge(15, 93) <= 4; angryBirdLarge(15, 94) <= 4; angryBirdLarge(15, 95) <= 4; angryBirdLarge(15, 96) <= 5; angryBirdLarge(15, 97) <= 5; angryBirdLarge(15, 98) <= 5; angryBirdLarge(15, 99) <= 5; angryBirdLarge(15, 100) <= 5; angryBirdLarge(15, 101) <= 5; angryBirdLarge(15, 102) <= 0; angryBirdLarge(15, 103) <= 0; angryBirdLarge(15, 104) <= 0; angryBirdLarge(15, 105) <= 0; angryBirdLarge(15, 106) <= 0; angryBirdLarge(15, 107) <= 0; angryBirdLarge(15, 108) <= 0; angryBirdLarge(15, 109) <= 0; angryBirdLarge(15, 110) <= 0; angryBirdLarge(15, 111) <= 0; angryBirdLarge(15, 112) <= 0; angryBirdLarge(15, 113) <= 0; angryBirdLarge(15, 114) <= 0; angryBirdLarge(15, 115) <= 0; angryBirdLarge(15, 116) <= 0; angryBirdLarge(15, 117) <= 0; angryBirdLarge(15, 118) <= 0; angryBirdLarge(15, 119) <= 0; angryBirdLarge(15, 120) <= 0; angryBirdLarge(15, 121) <= 0; angryBirdLarge(15, 122) <= 0; angryBirdLarge(15, 123) <= 0; angryBirdLarge(15, 124) <= 0; angryBirdLarge(15, 125) <= 0; angryBirdLarge(15, 126) <= 0; angryBirdLarge(15, 127) <= 0; angryBirdLarge(15, 128) <= 0; angryBirdLarge(15, 129) <= 0; angryBirdLarge(15, 130) <= 0; angryBirdLarge(15, 131) <= 0; angryBirdLarge(15, 132) <= 0; angryBirdLarge(15, 133) <= 0; angryBirdLarge(15, 134) <= 0; angryBirdLarge(15, 135) <= 0; angryBirdLarge(15, 136) <= 0; angryBirdLarge(15, 137) <= 0; angryBirdLarge(15, 138) <= 0; angryBirdLarge(15, 139) <= 0; angryBirdLarge(15, 140) <= 0; angryBirdLarge(15, 141) <= 0; angryBirdLarge(15, 142) <= 0; angryBirdLarge(15, 143) <= 0; angryBirdLarge(15, 144) <= 0; angryBirdLarge(15, 145) <= 0; angryBirdLarge(15, 146) <= 0; angryBirdLarge(15, 147) <= 0; angryBirdLarge(15, 148) <= 0; angryBirdLarge(15, 149) <= 0; 
angryBirdLarge(16, 0) <= 0; angryBirdLarge(16, 1) <= 0; angryBirdLarge(16, 2) <= 0; angryBirdLarge(16, 3) <= 0; angryBirdLarge(16, 4) <= 0; angryBirdLarge(16, 5) <= 0; angryBirdLarge(16, 6) <= 0; angryBirdLarge(16, 7) <= 0; angryBirdLarge(16, 8) <= 0; angryBirdLarge(16, 9) <= 0; angryBirdLarge(16, 10) <= 0; angryBirdLarge(16, 11) <= 0; angryBirdLarge(16, 12) <= 0; angryBirdLarge(16, 13) <= 0; angryBirdLarge(16, 14) <= 0; angryBirdLarge(16, 15) <= 0; angryBirdLarge(16, 16) <= 0; angryBirdLarge(16, 17) <= 0; angryBirdLarge(16, 18) <= 0; angryBirdLarge(16, 19) <= 0; angryBirdLarge(16, 20) <= 0; angryBirdLarge(16, 21) <= 0; angryBirdLarge(16, 22) <= 0; angryBirdLarge(16, 23) <= 0; angryBirdLarge(16, 24) <= 0; angryBirdLarge(16, 25) <= 0; angryBirdLarge(16, 26) <= 0; angryBirdLarge(16, 27) <= 0; angryBirdLarge(16, 28) <= 0; angryBirdLarge(16, 29) <= 0; angryBirdLarge(16, 30) <= 0; angryBirdLarge(16, 31) <= 0; angryBirdLarge(16, 32) <= 0; angryBirdLarge(16, 33) <= 0; angryBirdLarge(16, 34) <= 0; angryBirdLarge(16, 35) <= 0; angryBirdLarge(16, 36) <= 0; angryBirdLarge(16, 37) <= 0; angryBirdLarge(16, 38) <= 0; angryBirdLarge(16, 39) <= 0; angryBirdLarge(16, 40) <= 0; angryBirdLarge(16, 41) <= 0; angryBirdLarge(16, 42) <= 0; angryBirdLarge(16, 43) <= 0; angryBirdLarge(16, 44) <= 0; angryBirdLarge(16, 45) <= 0; angryBirdLarge(16, 46) <= 0; angryBirdLarge(16, 47) <= 0; angryBirdLarge(16, 48) <= 5; angryBirdLarge(16, 49) <= 5; angryBirdLarge(16, 50) <= 5; angryBirdLarge(16, 51) <= 5; angryBirdLarge(16, 52) <= 5; angryBirdLarge(16, 53) <= 5; angryBirdLarge(16, 54) <= 5; angryBirdLarge(16, 55) <= 5; angryBirdLarge(16, 56) <= 5; angryBirdLarge(16, 57) <= 5; angryBirdLarge(16, 58) <= 5; angryBirdLarge(16, 59) <= 5; angryBirdLarge(16, 60) <= 5; angryBirdLarge(16, 61) <= 5; angryBirdLarge(16, 62) <= 5; angryBirdLarge(16, 63) <= 5; angryBirdLarge(16, 64) <= 5; angryBirdLarge(16, 65) <= 5; angryBirdLarge(16, 66) <= 5; angryBirdLarge(16, 67) <= 5; angryBirdLarge(16, 68) <= 5; angryBirdLarge(16, 69) <= 5; angryBirdLarge(16, 70) <= 5; angryBirdLarge(16, 71) <= 5; angryBirdLarge(16, 72) <= 4; angryBirdLarge(16, 73) <= 4; angryBirdLarge(16, 74) <= 4; angryBirdLarge(16, 75) <= 4; angryBirdLarge(16, 76) <= 4; angryBirdLarge(16, 77) <= 4; angryBirdLarge(16, 78) <= 4; angryBirdLarge(16, 79) <= 4; angryBirdLarge(16, 80) <= 4; angryBirdLarge(16, 81) <= 4; angryBirdLarge(16, 82) <= 4; angryBirdLarge(16, 83) <= 4; angryBirdLarge(16, 84) <= 4; angryBirdLarge(16, 85) <= 4; angryBirdLarge(16, 86) <= 4; angryBirdLarge(16, 87) <= 4; angryBirdLarge(16, 88) <= 4; angryBirdLarge(16, 89) <= 4; angryBirdLarge(16, 90) <= 4; angryBirdLarge(16, 91) <= 4; angryBirdLarge(16, 92) <= 4; angryBirdLarge(16, 93) <= 4; angryBirdLarge(16, 94) <= 4; angryBirdLarge(16, 95) <= 4; angryBirdLarge(16, 96) <= 5; angryBirdLarge(16, 97) <= 5; angryBirdLarge(16, 98) <= 5; angryBirdLarge(16, 99) <= 5; angryBirdLarge(16, 100) <= 5; angryBirdLarge(16, 101) <= 5; angryBirdLarge(16, 102) <= 0; angryBirdLarge(16, 103) <= 0; angryBirdLarge(16, 104) <= 0; angryBirdLarge(16, 105) <= 0; angryBirdLarge(16, 106) <= 0; angryBirdLarge(16, 107) <= 0; angryBirdLarge(16, 108) <= 0; angryBirdLarge(16, 109) <= 0; angryBirdLarge(16, 110) <= 0; angryBirdLarge(16, 111) <= 0; angryBirdLarge(16, 112) <= 0; angryBirdLarge(16, 113) <= 0; angryBirdLarge(16, 114) <= 0; angryBirdLarge(16, 115) <= 0; angryBirdLarge(16, 116) <= 0; angryBirdLarge(16, 117) <= 0; angryBirdLarge(16, 118) <= 0; angryBirdLarge(16, 119) <= 0; angryBirdLarge(16, 120) <= 0; angryBirdLarge(16, 121) <= 0; angryBirdLarge(16, 122) <= 0; angryBirdLarge(16, 123) <= 0; angryBirdLarge(16, 124) <= 0; angryBirdLarge(16, 125) <= 0; angryBirdLarge(16, 126) <= 0; angryBirdLarge(16, 127) <= 0; angryBirdLarge(16, 128) <= 0; angryBirdLarge(16, 129) <= 0; angryBirdLarge(16, 130) <= 0; angryBirdLarge(16, 131) <= 0; angryBirdLarge(16, 132) <= 0; angryBirdLarge(16, 133) <= 0; angryBirdLarge(16, 134) <= 0; angryBirdLarge(16, 135) <= 0; angryBirdLarge(16, 136) <= 0; angryBirdLarge(16, 137) <= 0; angryBirdLarge(16, 138) <= 0; angryBirdLarge(16, 139) <= 0; angryBirdLarge(16, 140) <= 0; angryBirdLarge(16, 141) <= 0; angryBirdLarge(16, 142) <= 0; angryBirdLarge(16, 143) <= 0; angryBirdLarge(16, 144) <= 0; angryBirdLarge(16, 145) <= 0; angryBirdLarge(16, 146) <= 0; angryBirdLarge(16, 147) <= 0; angryBirdLarge(16, 148) <= 0; angryBirdLarge(16, 149) <= 0; 
angryBirdLarge(17, 0) <= 0; angryBirdLarge(17, 1) <= 0; angryBirdLarge(17, 2) <= 0; angryBirdLarge(17, 3) <= 0; angryBirdLarge(17, 4) <= 0; angryBirdLarge(17, 5) <= 0; angryBirdLarge(17, 6) <= 0; angryBirdLarge(17, 7) <= 0; angryBirdLarge(17, 8) <= 0; angryBirdLarge(17, 9) <= 0; angryBirdLarge(17, 10) <= 0; angryBirdLarge(17, 11) <= 0; angryBirdLarge(17, 12) <= 0; angryBirdLarge(17, 13) <= 0; angryBirdLarge(17, 14) <= 0; angryBirdLarge(17, 15) <= 0; angryBirdLarge(17, 16) <= 0; angryBirdLarge(17, 17) <= 0; angryBirdLarge(17, 18) <= 0; angryBirdLarge(17, 19) <= 0; angryBirdLarge(17, 20) <= 0; angryBirdLarge(17, 21) <= 0; angryBirdLarge(17, 22) <= 0; angryBirdLarge(17, 23) <= 0; angryBirdLarge(17, 24) <= 0; angryBirdLarge(17, 25) <= 0; angryBirdLarge(17, 26) <= 0; angryBirdLarge(17, 27) <= 0; angryBirdLarge(17, 28) <= 0; angryBirdLarge(17, 29) <= 0; angryBirdLarge(17, 30) <= 0; angryBirdLarge(17, 31) <= 0; angryBirdLarge(17, 32) <= 0; angryBirdLarge(17, 33) <= 0; angryBirdLarge(17, 34) <= 0; angryBirdLarge(17, 35) <= 0; angryBirdLarge(17, 36) <= 0; angryBirdLarge(17, 37) <= 0; angryBirdLarge(17, 38) <= 0; angryBirdLarge(17, 39) <= 0; angryBirdLarge(17, 40) <= 0; angryBirdLarge(17, 41) <= 0; angryBirdLarge(17, 42) <= 0; angryBirdLarge(17, 43) <= 0; angryBirdLarge(17, 44) <= 0; angryBirdLarge(17, 45) <= 0; angryBirdLarge(17, 46) <= 0; angryBirdLarge(17, 47) <= 0; angryBirdLarge(17, 48) <= 5; angryBirdLarge(17, 49) <= 5; angryBirdLarge(17, 50) <= 5; angryBirdLarge(17, 51) <= 5; angryBirdLarge(17, 52) <= 5; angryBirdLarge(17, 53) <= 5; angryBirdLarge(17, 54) <= 5; angryBirdLarge(17, 55) <= 5; angryBirdLarge(17, 56) <= 5; angryBirdLarge(17, 57) <= 5; angryBirdLarge(17, 58) <= 5; angryBirdLarge(17, 59) <= 5; angryBirdLarge(17, 60) <= 5; angryBirdLarge(17, 61) <= 5; angryBirdLarge(17, 62) <= 5; angryBirdLarge(17, 63) <= 5; angryBirdLarge(17, 64) <= 5; angryBirdLarge(17, 65) <= 5; angryBirdLarge(17, 66) <= 5; angryBirdLarge(17, 67) <= 5; angryBirdLarge(17, 68) <= 5; angryBirdLarge(17, 69) <= 5; angryBirdLarge(17, 70) <= 5; angryBirdLarge(17, 71) <= 5; angryBirdLarge(17, 72) <= 4; angryBirdLarge(17, 73) <= 4; angryBirdLarge(17, 74) <= 4; angryBirdLarge(17, 75) <= 4; angryBirdLarge(17, 76) <= 4; angryBirdLarge(17, 77) <= 4; angryBirdLarge(17, 78) <= 4; angryBirdLarge(17, 79) <= 4; angryBirdLarge(17, 80) <= 4; angryBirdLarge(17, 81) <= 4; angryBirdLarge(17, 82) <= 4; angryBirdLarge(17, 83) <= 4; angryBirdLarge(17, 84) <= 4; angryBirdLarge(17, 85) <= 4; angryBirdLarge(17, 86) <= 4; angryBirdLarge(17, 87) <= 4; angryBirdLarge(17, 88) <= 4; angryBirdLarge(17, 89) <= 4; angryBirdLarge(17, 90) <= 4; angryBirdLarge(17, 91) <= 4; angryBirdLarge(17, 92) <= 4; angryBirdLarge(17, 93) <= 4; angryBirdLarge(17, 94) <= 4; angryBirdLarge(17, 95) <= 4; angryBirdLarge(17, 96) <= 5; angryBirdLarge(17, 97) <= 5; angryBirdLarge(17, 98) <= 5; angryBirdLarge(17, 99) <= 5; angryBirdLarge(17, 100) <= 5; angryBirdLarge(17, 101) <= 5; angryBirdLarge(17, 102) <= 0; angryBirdLarge(17, 103) <= 0; angryBirdLarge(17, 104) <= 0; angryBirdLarge(17, 105) <= 0; angryBirdLarge(17, 106) <= 0; angryBirdLarge(17, 107) <= 0; angryBirdLarge(17, 108) <= 0; angryBirdLarge(17, 109) <= 0; angryBirdLarge(17, 110) <= 0; angryBirdLarge(17, 111) <= 0; angryBirdLarge(17, 112) <= 0; angryBirdLarge(17, 113) <= 0; angryBirdLarge(17, 114) <= 0; angryBirdLarge(17, 115) <= 0; angryBirdLarge(17, 116) <= 0; angryBirdLarge(17, 117) <= 0; angryBirdLarge(17, 118) <= 0; angryBirdLarge(17, 119) <= 0; angryBirdLarge(17, 120) <= 0; angryBirdLarge(17, 121) <= 0; angryBirdLarge(17, 122) <= 0; angryBirdLarge(17, 123) <= 0; angryBirdLarge(17, 124) <= 0; angryBirdLarge(17, 125) <= 0; angryBirdLarge(17, 126) <= 0; angryBirdLarge(17, 127) <= 0; angryBirdLarge(17, 128) <= 0; angryBirdLarge(17, 129) <= 0; angryBirdLarge(17, 130) <= 0; angryBirdLarge(17, 131) <= 0; angryBirdLarge(17, 132) <= 0; angryBirdLarge(17, 133) <= 0; angryBirdLarge(17, 134) <= 0; angryBirdLarge(17, 135) <= 0; angryBirdLarge(17, 136) <= 0; angryBirdLarge(17, 137) <= 0; angryBirdLarge(17, 138) <= 0; angryBirdLarge(17, 139) <= 0; angryBirdLarge(17, 140) <= 0; angryBirdLarge(17, 141) <= 0; angryBirdLarge(17, 142) <= 0; angryBirdLarge(17, 143) <= 0; angryBirdLarge(17, 144) <= 0; angryBirdLarge(17, 145) <= 0; angryBirdLarge(17, 146) <= 0; angryBirdLarge(17, 147) <= 0; angryBirdLarge(17, 148) <= 0; angryBirdLarge(17, 149) <= 0; 
angryBirdLarge(18, 0) <= 0; angryBirdLarge(18, 1) <= 0; angryBirdLarge(18, 2) <= 0; angryBirdLarge(18, 3) <= 0; angryBirdLarge(18, 4) <= 0; angryBirdLarge(18, 5) <= 0; angryBirdLarge(18, 6) <= 0; angryBirdLarge(18, 7) <= 0; angryBirdLarge(18, 8) <= 0; angryBirdLarge(18, 9) <= 0; angryBirdLarge(18, 10) <= 0; angryBirdLarge(18, 11) <= 0; angryBirdLarge(18, 12) <= 0; angryBirdLarge(18, 13) <= 0; angryBirdLarge(18, 14) <= 0; angryBirdLarge(18, 15) <= 0; angryBirdLarge(18, 16) <= 0; angryBirdLarge(18, 17) <= 0; angryBirdLarge(18, 18) <= 0; angryBirdLarge(18, 19) <= 0; angryBirdLarge(18, 20) <= 0; angryBirdLarge(18, 21) <= 0; angryBirdLarge(18, 22) <= 0; angryBirdLarge(18, 23) <= 0; angryBirdLarge(18, 24) <= 0; angryBirdLarge(18, 25) <= 0; angryBirdLarge(18, 26) <= 0; angryBirdLarge(18, 27) <= 0; angryBirdLarge(18, 28) <= 0; angryBirdLarge(18, 29) <= 0; angryBirdLarge(18, 30) <= 0; angryBirdLarge(18, 31) <= 0; angryBirdLarge(18, 32) <= 0; angryBirdLarge(18, 33) <= 0; angryBirdLarge(18, 34) <= 0; angryBirdLarge(18, 35) <= 0; angryBirdLarge(18, 36) <= 0; angryBirdLarge(18, 37) <= 0; angryBirdLarge(18, 38) <= 0; angryBirdLarge(18, 39) <= 0; angryBirdLarge(18, 40) <= 0; angryBirdLarge(18, 41) <= 0; angryBirdLarge(18, 42) <= 5; angryBirdLarge(18, 43) <= 5; angryBirdLarge(18, 44) <= 5; angryBirdLarge(18, 45) <= 5; angryBirdLarge(18, 46) <= 5; angryBirdLarge(18, 47) <= 5; angryBirdLarge(18, 48) <= 4; angryBirdLarge(18, 49) <= 4; angryBirdLarge(18, 50) <= 4; angryBirdLarge(18, 51) <= 4; angryBirdLarge(18, 52) <= 4; angryBirdLarge(18, 53) <= 4; angryBirdLarge(18, 54) <= 4; angryBirdLarge(18, 55) <= 4; angryBirdLarge(18, 56) <= 4; angryBirdLarge(18, 57) <= 4; angryBirdLarge(18, 58) <= 4; angryBirdLarge(18, 59) <= 4; angryBirdLarge(18, 60) <= 4; angryBirdLarge(18, 61) <= 4; angryBirdLarge(18, 62) <= 4; angryBirdLarge(18, 63) <= 4; angryBirdLarge(18, 64) <= 4; angryBirdLarge(18, 65) <= 4; angryBirdLarge(18, 66) <= 4; angryBirdLarge(18, 67) <= 4; angryBirdLarge(18, 68) <= 4; angryBirdLarge(18, 69) <= 4; angryBirdLarge(18, 70) <= 4; angryBirdLarge(18, 71) <= 4; angryBirdLarge(18, 72) <= 4; angryBirdLarge(18, 73) <= 4; angryBirdLarge(18, 74) <= 4; angryBirdLarge(18, 75) <= 4; angryBirdLarge(18, 76) <= 4; angryBirdLarge(18, 77) <= 4; angryBirdLarge(18, 78) <= 4; angryBirdLarge(18, 79) <= 4; angryBirdLarge(18, 80) <= 4; angryBirdLarge(18, 81) <= 4; angryBirdLarge(18, 82) <= 4; angryBirdLarge(18, 83) <= 4; angryBirdLarge(18, 84) <= 4; angryBirdLarge(18, 85) <= 4; angryBirdLarge(18, 86) <= 4; angryBirdLarge(18, 87) <= 4; angryBirdLarge(18, 88) <= 4; angryBirdLarge(18, 89) <= 4; angryBirdLarge(18, 90) <= 4; angryBirdLarge(18, 91) <= 4; angryBirdLarge(18, 92) <= 4; angryBirdLarge(18, 93) <= 4; angryBirdLarge(18, 94) <= 4; angryBirdLarge(18, 95) <= 4; angryBirdLarge(18, 96) <= 4; angryBirdLarge(18, 97) <= 4; angryBirdLarge(18, 98) <= 4; angryBirdLarge(18, 99) <= 4; angryBirdLarge(18, 100) <= 4; angryBirdLarge(18, 101) <= 4; angryBirdLarge(18, 102) <= 5; angryBirdLarge(18, 103) <= 5; angryBirdLarge(18, 104) <= 5; angryBirdLarge(18, 105) <= 5; angryBirdLarge(18, 106) <= 5; angryBirdLarge(18, 107) <= 5; angryBirdLarge(18, 108) <= 0; angryBirdLarge(18, 109) <= 0; angryBirdLarge(18, 110) <= 0; angryBirdLarge(18, 111) <= 0; angryBirdLarge(18, 112) <= 0; angryBirdLarge(18, 113) <= 0; angryBirdLarge(18, 114) <= 0; angryBirdLarge(18, 115) <= 0; angryBirdLarge(18, 116) <= 0; angryBirdLarge(18, 117) <= 0; angryBirdLarge(18, 118) <= 0; angryBirdLarge(18, 119) <= 0; angryBirdLarge(18, 120) <= 0; angryBirdLarge(18, 121) <= 0; angryBirdLarge(18, 122) <= 0; angryBirdLarge(18, 123) <= 0; angryBirdLarge(18, 124) <= 0; angryBirdLarge(18, 125) <= 0; angryBirdLarge(18, 126) <= 0; angryBirdLarge(18, 127) <= 0; angryBirdLarge(18, 128) <= 0; angryBirdLarge(18, 129) <= 0; angryBirdLarge(18, 130) <= 0; angryBirdLarge(18, 131) <= 0; angryBirdLarge(18, 132) <= 0; angryBirdLarge(18, 133) <= 0; angryBirdLarge(18, 134) <= 0; angryBirdLarge(18, 135) <= 0; angryBirdLarge(18, 136) <= 0; angryBirdLarge(18, 137) <= 0; angryBirdLarge(18, 138) <= 0; angryBirdLarge(18, 139) <= 0; angryBirdLarge(18, 140) <= 0; angryBirdLarge(18, 141) <= 0; angryBirdLarge(18, 142) <= 0; angryBirdLarge(18, 143) <= 0; angryBirdLarge(18, 144) <= 0; angryBirdLarge(18, 145) <= 0; angryBirdLarge(18, 146) <= 0; angryBirdLarge(18, 147) <= 0; angryBirdLarge(18, 148) <= 0; angryBirdLarge(18, 149) <= 0; 
angryBirdLarge(19, 0) <= 0; angryBirdLarge(19, 1) <= 0; angryBirdLarge(19, 2) <= 0; angryBirdLarge(19, 3) <= 0; angryBirdLarge(19, 4) <= 0; angryBirdLarge(19, 5) <= 0; angryBirdLarge(19, 6) <= 0; angryBirdLarge(19, 7) <= 0; angryBirdLarge(19, 8) <= 0; angryBirdLarge(19, 9) <= 0; angryBirdLarge(19, 10) <= 0; angryBirdLarge(19, 11) <= 0; angryBirdLarge(19, 12) <= 0; angryBirdLarge(19, 13) <= 0; angryBirdLarge(19, 14) <= 0; angryBirdLarge(19, 15) <= 0; angryBirdLarge(19, 16) <= 0; angryBirdLarge(19, 17) <= 0; angryBirdLarge(19, 18) <= 0; angryBirdLarge(19, 19) <= 0; angryBirdLarge(19, 20) <= 0; angryBirdLarge(19, 21) <= 0; angryBirdLarge(19, 22) <= 0; angryBirdLarge(19, 23) <= 0; angryBirdLarge(19, 24) <= 0; angryBirdLarge(19, 25) <= 0; angryBirdLarge(19, 26) <= 0; angryBirdLarge(19, 27) <= 0; angryBirdLarge(19, 28) <= 0; angryBirdLarge(19, 29) <= 0; angryBirdLarge(19, 30) <= 0; angryBirdLarge(19, 31) <= 0; angryBirdLarge(19, 32) <= 0; angryBirdLarge(19, 33) <= 0; angryBirdLarge(19, 34) <= 0; angryBirdLarge(19, 35) <= 0; angryBirdLarge(19, 36) <= 0; angryBirdLarge(19, 37) <= 0; angryBirdLarge(19, 38) <= 0; angryBirdLarge(19, 39) <= 0; angryBirdLarge(19, 40) <= 0; angryBirdLarge(19, 41) <= 0; angryBirdLarge(19, 42) <= 5; angryBirdLarge(19, 43) <= 5; angryBirdLarge(19, 44) <= 5; angryBirdLarge(19, 45) <= 5; angryBirdLarge(19, 46) <= 5; angryBirdLarge(19, 47) <= 5; angryBirdLarge(19, 48) <= 4; angryBirdLarge(19, 49) <= 4; angryBirdLarge(19, 50) <= 4; angryBirdLarge(19, 51) <= 4; angryBirdLarge(19, 52) <= 4; angryBirdLarge(19, 53) <= 4; angryBirdLarge(19, 54) <= 4; angryBirdLarge(19, 55) <= 4; angryBirdLarge(19, 56) <= 4; angryBirdLarge(19, 57) <= 4; angryBirdLarge(19, 58) <= 4; angryBirdLarge(19, 59) <= 4; angryBirdLarge(19, 60) <= 4; angryBirdLarge(19, 61) <= 4; angryBirdLarge(19, 62) <= 4; angryBirdLarge(19, 63) <= 4; angryBirdLarge(19, 64) <= 4; angryBirdLarge(19, 65) <= 4; angryBirdLarge(19, 66) <= 4; angryBirdLarge(19, 67) <= 4; angryBirdLarge(19, 68) <= 4; angryBirdLarge(19, 69) <= 4; angryBirdLarge(19, 70) <= 4; angryBirdLarge(19, 71) <= 4; angryBirdLarge(19, 72) <= 4; angryBirdLarge(19, 73) <= 4; angryBirdLarge(19, 74) <= 4; angryBirdLarge(19, 75) <= 4; angryBirdLarge(19, 76) <= 4; angryBirdLarge(19, 77) <= 4; angryBirdLarge(19, 78) <= 4; angryBirdLarge(19, 79) <= 4; angryBirdLarge(19, 80) <= 4; angryBirdLarge(19, 81) <= 4; angryBirdLarge(19, 82) <= 4; angryBirdLarge(19, 83) <= 4; angryBirdLarge(19, 84) <= 4; angryBirdLarge(19, 85) <= 4; angryBirdLarge(19, 86) <= 4; angryBirdLarge(19, 87) <= 4; angryBirdLarge(19, 88) <= 4; angryBirdLarge(19, 89) <= 4; angryBirdLarge(19, 90) <= 4; angryBirdLarge(19, 91) <= 4; angryBirdLarge(19, 92) <= 4; angryBirdLarge(19, 93) <= 4; angryBirdLarge(19, 94) <= 4; angryBirdLarge(19, 95) <= 4; angryBirdLarge(19, 96) <= 4; angryBirdLarge(19, 97) <= 4; angryBirdLarge(19, 98) <= 4; angryBirdLarge(19, 99) <= 4; angryBirdLarge(19, 100) <= 4; angryBirdLarge(19, 101) <= 4; angryBirdLarge(19, 102) <= 5; angryBirdLarge(19, 103) <= 5; angryBirdLarge(19, 104) <= 5; angryBirdLarge(19, 105) <= 5; angryBirdLarge(19, 106) <= 5; angryBirdLarge(19, 107) <= 5; angryBirdLarge(19, 108) <= 0; angryBirdLarge(19, 109) <= 0; angryBirdLarge(19, 110) <= 0; angryBirdLarge(19, 111) <= 0; angryBirdLarge(19, 112) <= 0; angryBirdLarge(19, 113) <= 0; angryBirdLarge(19, 114) <= 0; angryBirdLarge(19, 115) <= 0; angryBirdLarge(19, 116) <= 0; angryBirdLarge(19, 117) <= 0; angryBirdLarge(19, 118) <= 0; angryBirdLarge(19, 119) <= 0; angryBirdLarge(19, 120) <= 0; angryBirdLarge(19, 121) <= 0; angryBirdLarge(19, 122) <= 0; angryBirdLarge(19, 123) <= 0; angryBirdLarge(19, 124) <= 0; angryBirdLarge(19, 125) <= 0; angryBirdLarge(19, 126) <= 0; angryBirdLarge(19, 127) <= 0; angryBirdLarge(19, 128) <= 0; angryBirdLarge(19, 129) <= 0; angryBirdLarge(19, 130) <= 0; angryBirdLarge(19, 131) <= 0; angryBirdLarge(19, 132) <= 0; angryBirdLarge(19, 133) <= 0; angryBirdLarge(19, 134) <= 0; angryBirdLarge(19, 135) <= 0; angryBirdLarge(19, 136) <= 0; angryBirdLarge(19, 137) <= 0; angryBirdLarge(19, 138) <= 0; angryBirdLarge(19, 139) <= 0; angryBirdLarge(19, 140) <= 0; angryBirdLarge(19, 141) <= 0; angryBirdLarge(19, 142) <= 0; angryBirdLarge(19, 143) <= 0; angryBirdLarge(19, 144) <= 0; angryBirdLarge(19, 145) <= 0; angryBirdLarge(19, 146) <= 0; angryBirdLarge(19, 147) <= 0; angryBirdLarge(19, 148) <= 0; angryBirdLarge(19, 149) <= 0; 
angryBirdLarge(20, 0) <= 0; angryBirdLarge(20, 1) <= 0; angryBirdLarge(20, 2) <= 0; angryBirdLarge(20, 3) <= 0; angryBirdLarge(20, 4) <= 0; angryBirdLarge(20, 5) <= 0; angryBirdLarge(20, 6) <= 0; angryBirdLarge(20, 7) <= 0; angryBirdLarge(20, 8) <= 0; angryBirdLarge(20, 9) <= 0; angryBirdLarge(20, 10) <= 0; angryBirdLarge(20, 11) <= 0; angryBirdLarge(20, 12) <= 0; angryBirdLarge(20, 13) <= 0; angryBirdLarge(20, 14) <= 0; angryBirdLarge(20, 15) <= 0; angryBirdLarge(20, 16) <= 0; angryBirdLarge(20, 17) <= 0; angryBirdLarge(20, 18) <= 0; angryBirdLarge(20, 19) <= 0; angryBirdLarge(20, 20) <= 0; angryBirdLarge(20, 21) <= 0; angryBirdLarge(20, 22) <= 0; angryBirdLarge(20, 23) <= 0; angryBirdLarge(20, 24) <= 0; angryBirdLarge(20, 25) <= 0; angryBirdLarge(20, 26) <= 0; angryBirdLarge(20, 27) <= 0; angryBirdLarge(20, 28) <= 0; angryBirdLarge(20, 29) <= 0; angryBirdLarge(20, 30) <= 0; angryBirdLarge(20, 31) <= 0; angryBirdLarge(20, 32) <= 0; angryBirdLarge(20, 33) <= 0; angryBirdLarge(20, 34) <= 0; angryBirdLarge(20, 35) <= 0; angryBirdLarge(20, 36) <= 0; angryBirdLarge(20, 37) <= 0; angryBirdLarge(20, 38) <= 0; angryBirdLarge(20, 39) <= 0; angryBirdLarge(20, 40) <= 0; angryBirdLarge(20, 41) <= 0; angryBirdLarge(20, 42) <= 5; angryBirdLarge(20, 43) <= 5; angryBirdLarge(20, 44) <= 5; angryBirdLarge(20, 45) <= 5; angryBirdLarge(20, 46) <= 5; angryBirdLarge(20, 47) <= 5; angryBirdLarge(20, 48) <= 4; angryBirdLarge(20, 49) <= 4; angryBirdLarge(20, 50) <= 4; angryBirdLarge(20, 51) <= 4; angryBirdLarge(20, 52) <= 4; angryBirdLarge(20, 53) <= 4; angryBirdLarge(20, 54) <= 4; angryBirdLarge(20, 55) <= 4; angryBirdLarge(20, 56) <= 4; angryBirdLarge(20, 57) <= 4; angryBirdLarge(20, 58) <= 4; angryBirdLarge(20, 59) <= 4; angryBirdLarge(20, 60) <= 4; angryBirdLarge(20, 61) <= 4; angryBirdLarge(20, 62) <= 4; angryBirdLarge(20, 63) <= 4; angryBirdLarge(20, 64) <= 4; angryBirdLarge(20, 65) <= 4; angryBirdLarge(20, 66) <= 4; angryBirdLarge(20, 67) <= 4; angryBirdLarge(20, 68) <= 4; angryBirdLarge(20, 69) <= 4; angryBirdLarge(20, 70) <= 4; angryBirdLarge(20, 71) <= 4; angryBirdLarge(20, 72) <= 4; angryBirdLarge(20, 73) <= 4; angryBirdLarge(20, 74) <= 4; angryBirdLarge(20, 75) <= 4; angryBirdLarge(20, 76) <= 4; angryBirdLarge(20, 77) <= 4; angryBirdLarge(20, 78) <= 4; angryBirdLarge(20, 79) <= 4; angryBirdLarge(20, 80) <= 4; angryBirdLarge(20, 81) <= 4; angryBirdLarge(20, 82) <= 4; angryBirdLarge(20, 83) <= 4; angryBirdLarge(20, 84) <= 4; angryBirdLarge(20, 85) <= 4; angryBirdLarge(20, 86) <= 4; angryBirdLarge(20, 87) <= 4; angryBirdLarge(20, 88) <= 4; angryBirdLarge(20, 89) <= 4; angryBirdLarge(20, 90) <= 4; angryBirdLarge(20, 91) <= 4; angryBirdLarge(20, 92) <= 4; angryBirdLarge(20, 93) <= 4; angryBirdLarge(20, 94) <= 4; angryBirdLarge(20, 95) <= 4; angryBirdLarge(20, 96) <= 4; angryBirdLarge(20, 97) <= 4; angryBirdLarge(20, 98) <= 4; angryBirdLarge(20, 99) <= 4; angryBirdLarge(20, 100) <= 4; angryBirdLarge(20, 101) <= 4; angryBirdLarge(20, 102) <= 5; angryBirdLarge(20, 103) <= 5; angryBirdLarge(20, 104) <= 5; angryBirdLarge(20, 105) <= 5; angryBirdLarge(20, 106) <= 5; angryBirdLarge(20, 107) <= 5; angryBirdLarge(20, 108) <= 0; angryBirdLarge(20, 109) <= 0; angryBirdLarge(20, 110) <= 0; angryBirdLarge(20, 111) <= 0; angryBirdLarge(20, 112) <= 0; angryBirdLarge(20, 113) <= 0; angryBirdLarge(20, 114) <= 0; angryBirdLarge(20, 115) <= 0; angryBirdLarge(20, 116) <= 0; angryBirdLarge(20, 117) <= 0; angryBirdLarge(20, 118) <= 0; angryBirdLarge(20, 119) <= 0; angryBirdLarge(20, 120) <= 0; angryBirdLarge(20, 121) <= 0; angryBirdLarge(20, 122) <= 0; angryBirdLarge(20, 123) <= 0; angryBirdLarge(20, 124) <= 0; angryBirdLarge(20, 125) <= 0; angryBirdLarge(20, 126) <= 0; angryBirdLarge(20, 127) <= 0; angryBirdLarge(20, 128) <= 0; angryBirdLarge(20, 129) <= 0; angryBirdLarge(20, 130) <= 0; angryBirdLarge(20, 131) <= 0; angryBirdLarge(20, 132) <= 0; angryBirdLarge(20, 133) <= 0; angryBirdLarge(20, 134) <= 0; angryBirdLarge(20, 135) <= 0; angryBirdLarge(20, 136) <= 0; angryBirdLarge(20, 137) <= 0; angryBirdLarge(20, 138) <= 0; angryBirdLarge(20, 139) <= 0; angryBirdLarge(20, 140) <= 0; angryBirdLarge(20, 141) <= 0; angryBirdLarge(20, 142) <= 0; angryBirdLarge(20, 143) <= 0; angryBirdLarge(20, 144) <= 0; angryBirdLarge(20, 145) <= 0; angryBirdLarge(20, 146) <= 0; angryBirdLarge(20, 147) <= 0; angryBirdLarge(20, 148) <= 0; angryBirdLarge(20, 149) <= 0; 
angryBirdLarge(21, 0) <= 0; angryBirdLarge(21, 1) <= 0; angryBirdLarge(21, 2) <= 0; angryBirdLarge(21, 3) <= 0; angryBirdLarge(21, 4) <= 0; angryBirdLarge(21, 5) <= 0; angryBirdLarge(21, 6) <= 0; angryBirdLarge(21, 7) <= 0; angryBirdLarge(21, 8) <= 0; angryBirdLarge(21, 9) <= 0; angryBirdLarge(21, 10) <= 0; angryBirdLarge(21, 11) <= 0; angryBirdLarge(21, 12) <= 0; angryBirdLarge(21, 13) <= 0; angryBirdLarge(21, 14) <= 0; angryBirdLarge(21, 15) <= 0; angryBirdLarge(21, 16) <= 0; angryBirdLarge(21, 17) <= 0; angryBirdLarge(21, 18) <= 0; angryBirdLarge(21, 19) <= 0; angryBirdLarge(21, 20) <= 0; angryBirdLarge(21, 21) <= 0; angryBirdLarge(21, 22) <= 0; angryBirdLarge(21, 23) <= 0; angryBirdLarge(21, 24) <= 0; angryBirdLarge(21, 25) <= 0; angryBirdLarge(21, 26) <= 0; angryBirdLarge(21, 27) <= 0; angryBirdLarge(21, 28) <= 0; angryBirdLarge(21, 29) <= 0; angryBirdLarge(21, 30) <= 0; angryBirdLarge(21, 31) <= 0; angryBirdLarge(21, 32) <= 0; angryBirdLarge(21, 33) <= 0; angryBirdLarge(21, 34) <= 0; angryBirdLarge(21, 35) <= 0; angryBirdLarge(21, 36) <= 0; angryBirdLarge(21, 37) <= 0; angryBirdLarge(21, 38) <= 0; angryBirdLarge(21, 39) <= 0; angryBirdLarge(21, 40) <= 0; angryBirdLarge(21, 41) <= 0; angryBirdLarge(21, 42) <= 5; angryBirdLarge(21, 43) <= 5; angryBirdLarge(21, 44) <= 5; angryBirdLarge(21, 45) <= 5; angryBirdLarge(21, 46) <= 5; angryBirdLarge(21, 47) <= 5; angryBirdLarge(21, 48) <= 4; angryBirdLarge(21, 49) <= 4; angryBirdLarge(21, 50) <= 4; angryBirdLarge(21, 51) <= 4; angryBirdLarge(21, 52) <= 4; angryBirdLarge(21, 53) <= 4; angryBirdLarge(21, 54) <= 4; angryBirdLarge(21, 55) <= 4; angryBirdLarge(21, 56) <= 4; angryBirdLarge(21, 57) <= 4; angryBirdLarge(21, 58) <= 4; angryBirdLarge(21, 59) <= 4; angryBirdLarge(21, 60) <= 4; angryBirdLarge(21, 61) <= 4; angryBirdLarge(21, 62) <= 4; angryBirdLarge(21, 63) <= 4; angryBirdLarge(21, 64) <= 4; angryBirdLarge(21, 65) <= 4; angryBirdLarge(21, 66) <= 4; angryBirdLarge(21, 67) <= 4; angryBirdLarge(21, 68) <= 4; angryBirdLarge(21, 69) <= 4; angryBirdLarge(21, 70) <= 4; angryBirdLarge(21, 71) <= 4; angryBirdLarge(21, 72) <= 4; angryBirdLarge(21, 73) <= 4; angryBirdLarge(21, 74) <= 4; angryBirdLarge(21, 75) <= 4; angryBirdLarge(21, 76) <= 4; angryBirdLarge(21, 77) <= 4; angryBirdLarge(21, 78) <= 4; angryBirdLarge(21, 79) <= 4; angryBirdLarge(21, 80) <= 4; angryBirdLarge(21, 81) <= 4; angryBirdLarge(21, 82) <= 4; angryBirdLarge(21, 83) <= 4; angryBirdLarge(21, 84) <= 4; angryBirdLarge(21, 85) <= 4; angryBirdLarge(21, 86) <= 4; angryBirdLarge(21, 87) <= 4; angryBirdLarge(21, 88) <= 4; angryBirdLarge(21, 89) <= 4; angryBirdLarge(21, 90) <= 4; angryBirdLarge(21, 91) <= 4; angryBirdLarge(21, 92) <= 4; angryBirdLarge(21, 93) <= 4; angryBirdLarge(21, 94) <= 4; angryBirdLarge(21, 95) <= 4; angryBirdLarge(21, 96) <= 4; angryBirdLarge(21, 97) <= 4; angryBirdLarge(21, 98) <= 4; angryBirdLarge(21, 99) <= 4; angryBirdLarge(21, 100) <= 4; angryBirdLarge(21, 101) <= 4; angryBirdLarge(21, 102) <= 5; angryBirdLarge(21, 103) <= 5; angryBirdLarge(21, 104) <= 5; angryBirdLarge(21, 105) <= 5; angryBirdLarge(21, 106) <= 5; angryBirdLarge(21, 107) <= 5; angryBirdLarge(21, 108) <= 0; angryBirdLarge(21, 109) <= 0; angryBirdLarge(21, 110) <= 0; angryBirdLarge(21, 111) <= 0; angryBirdLarge(21, 112) <= 0; angryBirdLarge(21, 113) <= 0; angryBirdLarge(21, 114) <= 0; angryBirdLarge(21, 115) <= 0; angryBirdLarge(21, 116) <= 0; angryBirdLarge(21, 117) <= 0; angryBirdLarge(21, 118) <= 0; angryBirdLarge(21, 119) <= 0; angryBirdLarge(21, 120) <= 0; angryBirdLarge(21, 121) <= 0; angryBirdLarge(21, 122) <= 0; angryBirdLarge(21, 123) <= 0; angryBirdLarge(21, 124) <= 0; angryBirdLarge(21, 125) <= 0; angryBirdLarge(21, 126) <= 0; angryBirdLarge(21, 127) <= 0; angryBirdLarge(21, 128) <= 0; angryBirdLarge(21, 129) <= 0; angryBirdLarge(21, 130) <= 0; angryBirdLarge(21, 131) <= 0; angryBirdLarge(21, 132) <= 0; angryBirdLarge(21, 133) <= 0; angryBirdLarge(21, 134) <= 0; angryBirdLarge(21, 135) <= 0; angryBirdLarge(21, 136) <= 0; angryBirdLarge(21, 137) <= 0; angryBirdLarge(21, 138) <= 0; angryBirdLarge(21, 139) <= 0; angryBirdLarge(21, 140) <= 0; angryBirdLarge(21, 141) <= 0; angryBirdLarge(21, 142) <= 0; angryBirdLarge(21, 143) <= 0; angryBirdLarge(21, 144) <= 0; angryBirdLarge(21, 145) <= 0; angryBirdLarge(21, 146) <= 0; angryBirdLarge(21, 147) <= 0; angryBirdLarge(21, 148) <= 0; angryBirdLarge(21, 149) <= 0; 
angryBirdLarge(22, 0) <= 0; angryBirdLarge(22, 1) <= 0; angryBirdLarge(22, 2) <= 0; angryBirdLarge(22, 3) <= 0; angryBirdLarge(22, 4) <= 0; angryBirdLarge(22, 5) <= 0; angryBirdLarge(22, 6) <= 0; angryBirdLarge(22, 7) <= 0; angryBirdLarge(22, 8) <= 0; angryBirdLarge(22, 9) <= 0; angryBirdLarge(22, 10) <= 0; angryBirdLarge(22, 11) <= 0; angryBirdLarge(22, 12) <= 0; angryBirdLarge(22, 13) <= 0; angryBirdLarge(22, 14) <= 0; angryBirdLarge(22, 15) <= 0; angryBirdLarge(22, 16) <= 0; angryBirdLarge(22, 17) <= 0; angryBirdLarge(22, 18) <= 0; angryBirdLarge(22, 19) <= 0; angryBirdLarge(22, 20) <= 0; angryBirdLarge(22, 21) <= 0; angryBirdLarge(22, 22) <= 0; angryBirdLarge(22, 23) <= 0; angryBirdLarge(22, 24) <= 0; angryBirdLarge(22, 25) <= 0; angryBirdLarge(22, 26) <= 0; angryBirdLarge(22, 27) <= 0; angryBirdLarge(22, 28) <= 0; angryBirdLarge(22, 29) <= 0; angryBirdLarge(22, 30) <= 0; angryBirdLarge(22, 31) <= 0; angryBirdLarge(22, 32) <= 0; angryBirdLarge(22, 33) <= 0; angryBirdLarge(22, 34) <= 0; angryBirdLarge(22, 35) <= 0; angryBirdLarge(22, 36) <= 0; angryBirdLarge(22, 37) <= 0; angryBirdLarge(22, 38) <= 0; angryBirdLarge(22, 39) <= 0; angryBirdLarge(22, 40) <= 0; angryBirdLarge(22, 41) <= 0; angryBirdLarge(22, 42) <= 5; angryBirdLarge(22, 43) <= 5; angryBirdLarge(22, 44) <= 5; angryBirdLarge(22, 45) <= 5; angryBirdLarge(22, 46) <= 5; angryBirdLarge(22, 47) <= 5; angryBirdLarge(22, 48) <= 4; angryBirdLarge(22, 49) <= 4; angryBirdLarge(22, 50) <= 4; angryBirdLarge(22, 51) <= 4; angryBirdLarge(22, 52) <= 4; angryBirdLarge(22, 53) <= 4; angryBirdLarge(22, 54) <= 4; angryBirdLarge(22, 55) <= 4; angryBirdLarge(22, 56) <= 4; angryBirdLarge(22, 57) <= 4; angryBirdLarge(22, 58) <= 4; angryBirdLarge(22, 59) <= 4; angryBirdLarge(22, 60) <= 4; angryBirdLarge(22, 61) <= 4; angryBirdLarge(22, 62) <= 4; angryBirdLarge(22, 63) <= 4; angryBirdLarge(22, 64) <= 4; angryBirdLarge(22, 65) <= 4; angryBirdLarge(22, 66) <= 4; angryBirdLarge(22, 67) <= 4; angryBirdLarge(22, 68) <= 4; angryBirdLarge(22, 69) <= 4; angryBirdLarge(22, 70) <= 4; angryBirdLarge(22, 71) <= 4; angryBirdLarge(22, 72) <= 4; angryBirdLarge(22, 73) <= 4; angryBirdLarge(22, 74) <= 4; angryBirdLarge(22, 75) <= 4; angryBirdLarge(22, 76) <= 4; angryBirdLarge(22, 77) <= 4; angryBirdLarge(22, 78) <= 4; angryBirdLarge(22, 79) <= 4; angryBirdLarge(22, 80) <= 4; angryBirdLarge(22, 81) <= 4; angryBirdLarge(22, 82) <= 4; angryBirdLarge(22, 83) <= 4; angryBirdLarge(22, 84) <= 4; angryBirdLarge(22, 85) <= 4; angryBirdLarge(22, 86) <= 4; angryBirdLarge(22, 87) <= 4; angryBirdLarge(22, 88) <= 4; angryBirdLarge(22, 89) <= 4; angryBirdLarge(22, 90) <= 4; angryBirdLarge(22, 91) <= 4; angryBirdLarge(22, 92) <= 4; angryBirdLarge(22, 93) <= 4; angryBirdLarge(22, 94) <= 4; angryBirdLarge(22, 95) <= 4; angryBirdLarge(22, 96) <= 4; angryBirdLarge(22, 97) <= 4; angryBirdLarge(22, 98) <= 4; angryBirdLarge(22, 99) <= 4; angryBirdLarge(22, 100) <= 4; angryBirdLarge(22, 101) <= 4; angryBirdLarge(22, 102) <= 5; angryBirdLarge(22, 103) <= 5; angryBirdLarge(22, 104) <= 5; angryBirdLarge(22, 105) <= 5; angryBirdLarge(22, 106) <= 5; angryBirdLarge(22, 107) <= 5; angryBirdLarge(22, 108) <= 0; angryBirdLarge(22, 109) <= 0; angryBirdLarge(22, 110) <= 0; angryBirdLarge(22, 111) <= 0; angryBirdLarge(22, 112) <= 0; angryBirdLarge(22, 113) <= 0; angryBirdLarge(22, 114) <= 0; angryBirdLarge(22, 115) <= 0; angryBirdLarge(22, 116) <= 0; angryBirdLarge(22, 117) <= 0; angryBirdLarge(22, 118) <= 0; angryBirdLarge(22, 119) <= 0; angryBirdLarge(22, 120) <= 0; angryBirdLarge(22, 121) <= 0; angryBirdLarge(22, 122) <= 0; angryBirdLarge(22, 123) <= 0; angryBirdLarge(22, 124) <= 0; angryBirdLarge(22, 125) <= 0; angryBirdLarge(22, 126) <= 0; angryBirdLarge(22, 127) <= 0; angryBirdLarge(22, 128) <= 0; angryBirdLarge(22, 129) <= 0; angryBirdLarge(22, 130) <= 0; angryBirdLarge(22, 131) <= 0; angryBirdLarge(22, 132) <= 0; angryBirdLarge(22, 133) <= 0; angryBirdLarge(22, 134) <= 0; angryBirdLarge(22, 135) <= 0; angryBirdLarge(22, 136) <= 0; angryBirdLarge(22, 137) <= 0; angryBirdLarge(22, 138) <= 0; angryBirdLarge(22, 139) <= 0; angryBirdLarge(22, 140) <= 0; angryBirdLarge(22, 141) <= 0; angryBirdLarge(22, 142) <= 0; angryBirdLarge(22, 143) <= 0; angryBirdLarge(22, 144) <= 0; angryBirdLarge(22, 145) <= 0; angryBirdLarge(22, 146) <= 0; angryBirdLarge(22, 147) <= 0; angryBirdLarge(22, 148) <= 0; angryBirdLarge(22, 149) <= 0; 
angryBirdLarge(23, 0) <= 0; angryBirdLarge(23, 1) <= 0; angryBirdLarge(23, 2) <= 0; angryBirdLarge(23, 3) <= 0; angryBirdLarge(23, 4) <= 0; angryBirdLarge(23, 5) <= 0; angryBirdLarge(23, 6) <= 0; angryBirdLarge(23, 7) <= 0; angryBirdLarge(23, 8) <= 0; angryBirdLarge(23, 9) <= 0; angryBirdLarge(23, 10) <= 0; angryBirdLarge(23, 11) <= 0; angryBirdLarge(23, 12) <= 0; angryBirdLarge(23, 13) <= 0; angryBirdLarge(23, 14) <= 0; angryBirdLarge(23, 15) <= 0; angryBirdLarge(23, 16) <= 0; angryBirdLarge(23, 17) <= 0; angryBirdLarge(23, 18) <= 0; angryBirdLarge(23, 19) <= 0; angryBirdLarge(23, 20) <= 0; angryBirdLarge(23, 21) <= 0; angryBirdLarge(23, 22) <= 0; angryBirdLarge(23, 23) <= 0; angryBirdLarge(23, 24) <= 0; angryBirdLarge(23, 25) <= 0; angryBirdLarge(23, 26) <= 0; angryBirdLarge(23, 27) <= 0; angryBirdLarge(23, 28) <= 0; angryBirdLarge(23, 29) <= 0; angryBirdLarge(23, 30) <= 0; angryBirdLarge(23, 31) <= 0; angryBirdLarge(23, 32) <= 0; angryBirdLarge(23, 33) <= 0; angryBirdLarge(23, 34) <= 0; angryBirdLarge(23, 35) <= 0; angryBirdLarge(23, 36) <= 0; angryBirdLarge(23, 37) <= 0; angryBirdLarge(23, 38) <= 0; angryBirdLarge(23, 39) <= 0; angryBirdLarge(23, 40) <= 0; angryBirdLarge(23, 41) <= 0; angryBirdLarge(23, 42) <= 5; angryBirdLarge(23, 43) <= 5; angryBirdLarge(23, 44) <= 5; angryBirdLarge(23, 45) <= 5; angryBirdLarge(23, 46) <= 5; angryBirdLarge(23, 47) <= 5; angryBirdLarge(23, 48) <= 4; angryBirdLarge(23, 49) <= 4; angryBirdLarge(23, 50) <= 4; angryBirdLarge(23, 51) <= 4; angryBirdLarge(23, 52) <= 4; angryBirdLarge(23, 53) <= 4; angryBirdLarge(23, 54) <= 4; angryBirdLarge(23, 55) <= 4; angryBirdLarge(23, 56) <= 4; angryBirdLarge(23, 57) <= 4; angryBirdLarge(23, 58) <= 4; angryBirdLarge(23, 59) <= 4; angryBirdLarge(23, 60) <= 4; angryBirdLarge(23, 61) <= 4; angryBirdLarge(23, 62) <= 4; angryBirdLarge(23, 63) <= 4; angryBirdLarge(23, 64) <= 4; angryBirdLarge(23, 65) <= 4; angryBirdLarge(23, 66) <= 4; angryBirdLarge(23, 67) <= 4; angryBirdLarge(23, 68) <= 4; angryBirdLarge(23, 69) <= 4; angryBirdLarge(23, 70) <= 4; angryBirdLarge(23, 71) <= 4; angryBirdLarge(23, 72) <= 4; angryBirdLarge(23, 73) <= 4; angryBirdLarge(23, 74) <= 4; angryBirdLarge(23, 75) <= 4; angryBirdLarge(23, 76) <= 4; angryBirdLarge(23, 77) <= 4; angryBirdLarge(23, 78) <= 4; angryBirdLarge(23, 79) <= 4; angryBirdLarge(23, 80) <= 4; angryBirdLarge(23, 81) <= 4; angryBirdLarge(23, 82) <= 4; angryBirdLarge(23, 83) <= 4; angryBirdLarge(23, 84) <= 4; angryBirdLarge(23, 85) <= 4; angryBirdLarge(23, 86) <= 4; angryBirdLarge(23, 87) <= 4; angryBirdLarge(23, 88) <= 4; angryBirdLarge(23, 89) <= 4; angryBirdLarge(23, 90) <= 4; angryBirdLarge(23, 91) <= 4; angryBirdLarge(23, 92) <= 4; angryBirdLarge(23, 93) <= 4; angryBirdLarge(23, 94) <= 4; angryBirdLarge(23, 95) <= 4; angryBirdLarge(23, 96) <= 4; angryBirdLarge(23, 97) <= 4; angryBirdLarge(23, 98) <= 4; angryBirdLarge(23, 99) <= 4; angryBirdLarge(23, 100) <= 4; angryBirdLarge(23, 101) <= 4; angryBirdLarge(23, 102) <= 5; angryBirdLarge(23, 103) <= 5; angryBirdLarge(23, 104) <= 5; angryBirdLarge(23, 105) <= 5; angryBirdLarge(23, 106) <= 5; angryBirdLarge(23, 107) <= 5; angryBirdLarge(23, 108) <= 0; angryBirdLarge(23, 109) <= 0; angryBirdLarge(23, 110) <= 0; angryBirdLarge(23, 111) <= 0; angryBirdLarge(23, 112) <= 0; angryBirdLarge(23, 113) <= 0; angryBirdLarge(23, 114) <= 0; angryBirdLarge(23, 115) <= 0; angryBirdLarge(23, 116) <= 0; angryBirdLarge(23, 117) <= 0; angryBirdLarge(23, 118) <= 0; angryBirdLarge(23, 119) <= 0; angryBirdLarge(23, 120) <= 0; angryBirdLarge(23, 121) <= 0; angryBirdLarge(23, 122) <= 0; angryBirdLarge(23, 123) <= 0; angryBirdLarge(23, 124) <= 0; angryBirdLarge(23, 125) <= 0; angryBirdLarge(23, 126) <= 0; angryBirdLarge(23, 127) <= 0; angryBirdLarge(23, 128) <= 0; angryBirdLarge(23, 129) <= 0; angryBirdLarge(23, 130) <= 0; angryBirdLarge(23, 131) <= 0; angryBirdLarge(23, 132) <= 0; angryBirdLarge(23, 133) <= 0; angryBirdLarge(23, 134) <= 0; angryBirdLarge(23, 135) <= 0; angryBirdLarge(23, 136) <= 0; angryBirdLarge(23, 137) <= 0; angryBirdLarge(23, 138) <= 0; angryBirdLarge(23, 139) <= 0; angryBirdLarge(23, 140) <= 0; angryBirdLarge(23, 141) <= 0; angryBirdLarge(23, 142) <= 0; angryBirdLarge(23, 143) <= 0; angryBirdLarge(23, 144) <= 0; angryBirdLarge(23, 145) <= 0; angryBirdLarge(23, 146) <= 0; angryBirdLarge(23, 147) <= 0; angryBirdLarge(23, 148) <= 0; angryBirdLarge(23, 149) <= 0; 
angryBirdLarge(24, 0) <= 0; angryBirdLarge(24, 1) <= 0; angryBirdLarge(24, 2) <= 0; angryBirdLarge(24, 3) <= 0; angryBirdLarge(24, 4) <= 0; angryBirdLarge(24, 5) <= 0; angryBirdLarge(24, 6) <= 0; angryBirdLarge(24, 7) <= 0; angryBirdLarge(24, 8) <= 0; angryBirdLarge(24, 9) <= 0; angryBirdLarge(24, 10) <= 0; angryBirdLarge(24, 11) <= 0; angryBirdLarge(24, 12) <= 0; angryBirdLarge(24, 13) <= 0; angryBirdLarge(24, 14) <= 0; angryBirdLarge(24, 15) <= 0; angryBirdLarge(24, 16) <= 0; angryBirdLarge(24, 17) <= 0; angryBirdLarge(24, 18) <= 0; angryBirdLarge(24, 19) <= 0; angryBirdLarge(24, 20) <= 0; angryBirdLarge(24, 21) <= 0; angryBirdLarge(24, 22) <= 0; angryBirdLarge(24, 23) <= 0; angryBirdLarge(24, 24) <= 0; angryBirdLarge(24, 25) <= 0; angryBirdLarge(24, 26) <= 0; angryBirdLarge(24, 27) <= 0; angryBirdLarge(24, 28) <= 0; angryBirdLarge(24, 29) <= 0; angryBirdLarge(24, 30) <= 0; angryBirdLarge(24, 31) <= 0; angryBirdLarge(24, 32) <= 0; angryBirdLarge(24, 33) <= 0; angryBirdLarge(24, 34) <= 0; angryBirdLarge(24, 35) <= 0; angryBirdLarge(24, 36) <= 0; angryBirdLarge(24, 37) <= 0; angryBirdLarge(24, 38) <= 0; angryBirdLarge(24, 39) <= 0; angryBirdLarge(24, 40) <= 0; angryBirdLarge(24, 41) <= 0; angryBirdLarge(24, 42) <= 5; angryBirdLarge(24, 43) <= 5; angryBirdLarge(24, 44) <= 5; angryBirdLarge(24, 45) <= 5; angryBirdLarge(24, 46) <= 5; angryBirdLarge(24, 47) <= 5; angryBirdLarge(24, 48) <= 4; angryBirdLarge(24, 49) <= 4; angryBirdLarge(24, 50) <= 4; angryBirdLarge(24, 51) <= 4; angryBirdLarge(24, 52) <= 4; angryBirdLarge(24, 53) <= 4; angryBirdLarge(24, 54) <= 4; angryBirdLarge(24, 55) <= 4; angryBirdLarge(24, 56) <= 4; angryBirdLarge(24, 57) <= 4; angryBirdLarge(24, 58) <= 4; angryBirdLarge(24, 59) <= 4; angryBirdLarge(24, 60) <= 4; angryBirdLarge(24, 61) <= 4; angryBirdLarge(24, 62) <= 4; angryBirdLarge(24, 63) <= 4; angryBirdLarge(24, 64) <= 4; angryBirdLarge(24, 65) <= 4; angryBirdLarge(24, 66) <= 4; angryBirdLarge(24, 67) <= 4; angryBirdLarge(24, 68) <= 4; angryBirdLarge(24, 69) <= 4; angryBirdLarge(24, 70) <= 4; angryBirdLarge(24, 71) <= 4; angryBirdLarge(24, 72) <= 4; angryBirdLarge(24, 73) <= 4; angryBirdLarge(24, 74) <= 4; angryBirdLarge(24, 75) <= 4; angryBirdLarge(24, 76) <= 4; angryBirdLarge(24, 77) <= 4; angryBirdLarge(24, 78) <= 4; angryBirdLarge(24, 79) <= 4; angryBirdLarge(24, 80) <= 4; angryBirdLarge(24, 81) <= 4; angryBirdLarge(24, 82) <= 4; angryBirdLarge(24, 83) <= 4; angryBirdLarge(24, 84) <= 4; angryBirdLarge(24, 85) <= 4; angryBirdLarge(24, 86) <= 4; angryBirdLarge(24, 87) <= 4; angryBirdLarge(24, 88) <= 4; angryBirdLarge(24, 89) <= 4; angryBirdLarge(24, 90) <= 4; angryBirdLarge(24, 91) <= 4; angryBirdLarge(24, 92) <= 4; angryBirdLarge(24, 93) <= 4; angryBirdLarge(24, 94) <= 4; angryBirdLarge(24, 95) <= 4; angryBirdLarge(24, 96) <= 4; angryBirdLarge(24, 97) <= 4; angryBirdLarge(24, 98) <= 4; angryBirdLarge(24, 99) <= 4; angryBirdLarge(24, 100) <= 4; angryBirdLarge(24, 101) <= 4; angryBirdLarge(24, 102) <= 4; angryBirdLarge(24, 103) <= 4; angryBirdLarge(24, 104) <= 4; angryBirdLarge(24, 105) <= 4; angryBirdLarge(24, 106) <= 4; angryBirdLarge(24, 107) <= 4; angryBirdLarge(24, 108) <= 5; angryBirdLarge(24, 109) <= 5; angryBirdLarge(24, 110) <= 5; angryBirdLarge(24, 111) <= 5; angryBirdLarge(24, 112) <= 5; angryBirdLarge(24, 113) <= 5; angryBirdLarge(24, 114) <= 0; angryBirdLarge(24, 115) <= 0; angryBirdLarge(24, 116) <= 0; angryBirdLarge(24, 117) <= 0; angryBirdLarge(24, 118) <= 0; angryBirdLarge(24, 119) <= 0; angryBirdLarge(24, 120) <= 0; angryBirdLarge(24, 121) <= 0; angryBirdLarge(24, 122) <= 0; angryBirdLarge(24, 123) <= 0; angryBirdLarge(24, 124) <= 0; angryBirdLarge(24, 125) <= 0; angryBirdLarge(24, 126) <= 0; angryBirdLarge(24, 127) <= 0; angryBirdLarge(24, 128) <= 0; angryBirdLarge(24, 129) <= 0; angryBirdLarge(24, 130) <= 0; angryBirdLarge(24, 131) <= 0; angryBirdLarge(24, 132) <= 0; angryBirdLarge(24, 133) <= 0; angryBirdLarge(24, 134) <= 0; angryBirdLarge(24, 135) <= 0; angryBirdLarge(24, 136) <= 0; angryBirdLarge(24, 137) <= 0; angryBirdLarge(24, 138) <= 0; angryBirdLarge(24, 139) <= 0; angryBirdLarge(24, 140) <= 0; angryBirdLarge(24, 141) <= 0; angryBirdLarge(24, 142) <= 0; angryBirdLarge(24, 143) <= 0; angryBirdLarge(24, 144) <= 0; angryBirdLarge(24, 145) <= 0; angryBirdLarge(24, 146) <= 0; angryBirdLarge(24, 147) <= 0; angryBirdLarge(24, 148) <= 0; angryBirdLarge(24, 149) <= 0; 
angryBirdLarge(25, 0) <= 0; angryBirdLarge(25, 1) <= 0; angryBirdLarge(25, 2) <= 0; angryBirdLarge(25, 3) <= 0; angryBirdLarge(25, 4) <= 0; angryBirdLarge(25, 5) <= 0; angryBirdLarge(25, 6) <= 0; angryBirdLarge(25, 7) <= 0; angryBirdLarge(25, 8) <= 0; angryBirdLarge(25, 9) <= 0; angryBirdLarge(25, 10) <= 0; angryBirdLarge(25, 11) <= 0; angryBirdLarge(25, 12) <= 0; angryBirdLarge(25, 13) <= 0; angryBirdLarge(25, 14) <= 0; angryBirdLarge(25, 15) <= 0; angryBirdLarge(25, 16) <= 0; angryBirdLarge(25, 17) <= 0; angryBirdLarge(25, 18) <= 0; angryBirdLarge(25, 19) <= 0; angryBirdLarge(25, 20) <= 0; angryBirdLarge(25, 21) <= 0; angryBirdLarge(25, 22) <= 0; angryBirdLarge(25, 23) <= 0; angryBirdLarge(25, 24) <= 0; angryBirdLarge(25, 25) <= 0; angryBirdLarge(25, 26) <= 0; angryBirdLarge(25, 27) <= 0; angryBirdLarge(25, 28) <= 0; angryBirdLarge(25, 29) <= 0; angryBirdLarge(25, 30) <= 0; angryBirdLarge(25, 31) <= 0; angryBirdLarge(25, 32) <= 0; angryBirdLarge(25, 33) <= 0; angryBirdLarge(25, 34) <= 0; angryBirdLarge(25, 35) <= 0; angryBirdLarge(25, 36) <= 0; angryBirdLarge(25, 37) <= 0; angryBirdLarge(25, 38) <= 0; angryBirdLarge(25, 39) <= 0; angryBirdLarge(25, 40) <= 0; angryBirdLarge(25, 41) <= 0; angryBirdLarge(25, 42) <= 5; angryBirdLarge(25, 43) <= 5; angryBirdLarge(25, 44) <= 5; angryBirdLarge(25, 45) <= 5; angryBirdLarge(25, 46) <= 5; angryBirdLarge(25, 47) <= 5; angryBirdLarge(25, 48) <= 4; angryBirdLarge(25, 49) <= 4; angryBirdLarge(25, 50) <= 4; angryBirdLarge(25, 51) <= 4; angryBirdLarge(25, 52) <= 4; angryBirdLarge(25, 53) <= 4; angryBirdLarge(25, 54) <= 4; angryBirdLarge(25, 55) <= 4; angryBirdLarge(25, 56) <= 4; angryBirdLarge(25, 57) <= 4; angryBirdLarge(25, 58) <= 4; angryBirdLarge(25, 59) <= 4; angryBirdLarge(25, 60) <= 4; angryBirdLarge(25, 61) <= 4; angryBirdLarge(25, 62) <= 4; angryBirdLarge(25, 63) <= 4; angryBirdLarge(25, 64) <= 4; angryBirdLarge(25, 65) <= 4; angryBirdLarge(25, 66) <= 4; angryBirdLarge(25, 67) <= 4; angryBirdLarge(25, 68) <= 4; angryBirdLarge(25, 69) <= 4; angryBirdLarge(25, 70) <= 4; angryBirdLarge(25, 71) <= 4; angryBirdLarge(25, 72) <= 4; angryBirdLarge(25, 73) <= 4; angryBirdLarge(25, 74) <= 4; angryBirdLarge(25, 75) <= 4; angryBirdLarge(25, 76) <= 4; angryBirdLarge(25, 77) <= 4; angryBirdLarge(25, 78) <= 4; angryBirdLarge(25, 79) <= 4; angryBirdLarge(25, 80) <= 4; angryBirdLarge(25, 81) <= 4; angryBirdLarge(25, 82) <= 4; angryBirdLarge(25, 83) <= 4; angryBirdLarge(25, 84) <= 4; angryBirdLarge(25, 85) <= 4; angryBirdLarge(25, 86) <= 4; angryBirdLarge(25, 87) <= 4; angryBirdLarge(25, 88) <= 4; angryBirdLarge(25, 89) <= 4; angryBirdLarge(25, 90) <= 4; angryBirdLarge(25, 91) <= 4; angryBirdLarge(25, 92) <= 4; angryBirdLarge(25, 93) <= 4; angryBirdLarge(25, 94) <= 4; angryBirdLarge(25, 95) <= 4; angryBirdLarge(25, 96) <= 4; angryBirdLarge(25, 97) <= 4; angryBirdLarge(25, 98) <= 4; angryBirdLarge(25, 99) <= 4; angryBirdLarge(25, 100) <= 4; angryBirdLarge(25, 101) <= 4; angryBirdLarge(25, 102) <= 4; angryBirdLarge(25, 103) <= 4; angryBirdLarge(25, 104) <= 4; angryBirdLarge(25, 105) <= 4; angryBirdLarge(25, 106) <= 4; angryBirdLarge(25, 107) <= 4; angryBirdLarge(25, 108) <= 5; angryBirdLarge(25, 109) <= 5; angryBirdLarge(25, 110) <= 5; angryBirdLarge(25, 111) <= 5; angryBirdLarge(25, 112) <= 5; angryBirdLarge(25, 113) <= 5; angryBirdLarge(25, 114) <= 0; angryBirdLarge(25, 115) <= 0; angryBirdLarge(25, 116) <= 0; angryBirdLarge(25, 117) <= 0; angryBirdLarge(25, 118) <= 0; angryBirdLarge(25, 119) <= 0; angryBirdLarge(25, 120) <= 0; angryBirdLarge(25, 121) <= 0; angryBirdLarge(25, 122) <= 0; angryBirdLarge(25, 123) <= 0; angryBirdLarge(25, 124) <= 0; angryBirdLarge(25, 125) <= 0; angryBirdLarge(25, 126) <= 0; angryBirdLarge(25, 127) <= 0; angryBirdLarge(25, 128) <= 0; angryBirdLarge(25, 129) <= 0; angryBirdLarge(25, 130) <= 0; angryBirdLarge(25, 131) <= 0; angryBirdLarge(25, 132) <= 0; angryBirdLarge(25, 133) <= 0; angryBirdLarge(25, 134) <= 0; angryBirdLarge(25, 135) <= 0; angryBirdLarge(25, 136) <= 0; angryBirdLarge(25, 137) <= 0; angryBirdLarge(25, 138) <= 0; angryBirdLarge(25, 139) <= 0; angryBirdLarge(25, 140) <= 0; angryBirdLarge(25, 141) <= 0; angryBirdLarge(25, 142) <= 0; angryBirdLarge(25, 143) <= 0; angryBirdLarge(25, 144) <= 0; angryBirdLarge(25, 145) <= 0; angryBirdLarge(25, 146) <= 0; angryBirdLarge(25, 147) <= 0; angryBirdLarge(25, 148) <= 0; angryBirdLarge(25, 149) <= 0; 
angryBirdLarge(26, 0) <= 0; angryBirdLarge(26, 1) <= 0; angryBirdLarge(26, 2) <= 0; angryBirdLarge(26, 3) <= 0; angryBirdLarge(26, 4) <= 0; angryBirdLarge(26, 5) <= 0; angryBirdLarge(26, 6) <= 0; angryBirdLarge(26, 7) <= 0; angryBirdLarge(26, 8) <= 0; angryBirdLarge(26, 9) <= 0; angryBirdLarge(26, 10) <= 0; angryBirdLarge(26, 11) <= 0; angryBirdLarge(26, 12) <= 0; angryBirdLarge(26, 13) <= 0; angryBirdLarge(26, 14) <= 0; angryBirdLarge(26, 15) <= 0; angryBirdLarge(26, 16) <= 0; angryBirdLarge(26, 17) <= 0; angryBirdLarge(26, 18) <= 0; angryBirdLarge(26, 19) <= 0; angryBirdLarge(26, 20) <= 0; angryBirdLarge(26, 21) <= 0; angryBirdLarge(26, 22) <= 0; angryBirdLarge(26, 23) <= 0; angryBirdLarge(26, 24) <= 0; angryBirdLarge(26, 25) <= 0; angryBirdLarge(26, 26) <= 0; angryBirdLarge(26, 27) <= 0; angryBirdLarge(26, 28) <= 0; angryBirdLarge(26, 29) <= 0; angryBirdLarge(26, 30) <= 0; angryBirdLarge(26, 31) <= 0; angryBirdLarge(26, 32) <= 0; angryBirdLarge(26, 33) <= 0; angryBirdLarge(26, 34) <= 0; angryBirdLarge(26, 35) <= 0; angryBirdLarge(26, 36) <= 0; angryBirdLarge(26, 37) <= 0; angryBirdLarge(26, 38) <= 0; angryBirdLarge(26, 39) <= 0; angryBirdLarge(26, 40) <= 0; angryBirdLarge(26, 41) <= 0; angryBirdLarge(26, 42) <= 5; angryBirdLarge(26, 43) <= 5; angryBirdLarge(26, 44) <= 5; angryBirdLarge(26, 45) <= 5; angryBirdLarge(26, 46) <= 5; angryBirdLarge(26, 47) <= 5; angryBirdLarge(26, 48) <= 4; angryBirdLarge(26, 49) <= 4; angryBirdLarge(26, 50) <= 4; angryBirdLarge(26, 51) <= 4; angryBirdLarge(26, 52) <= 4; angryBirdLarge(26, 53) <= 4; angryBirdLarge(26, 54) <= 4; angryBirdLarge(26, 55) <= 4; angryBirdLarge(26, 56) <= 4; angryBirdLarge(26, 57) <= 4; angryBirdLarge(26, 58) <= 4; angryBirdLarge(26, 59) <= 4; angryBirdLarge(26, 60) <= 4; angryBirdLarge(26, 61) <= 4; angryBirdLarge(26, 62) <= 4; angryBirdLarge(26, 63) <= 4; angryBirdLarge(26, 64) <= 4; angryBirdLarge(26, 65) <= 4; angryBirdLarge(26, 66) <= 4; angryBirdLarge(26, 67) <= 4; angryBirdLarge(26, 68) <= 4; angryBirdLarge(26, 69) <= 4; angryBirdLarge(26, 70) <= 4; angryBirdLarge(26, 71) <= 4; angryBirdLarge(26, 72) <= 4; angryBirdLarge(26, 73) <= 4; angryBirdLarge(26, 74) <= 4; angryBirdLarge(26, 75) <= 4; angryBirdLarge(26, 76) <= 4; angryBirdLarge(26, 77) <= 4; angryBirdLarge(26, 78) <= 4; angryBirdLarge(26, 79) <= 4; angryBirdLarge(26, 80) <= 4; angryBirdLarge(26, 81) <= 4; angryBirdLarge(26, 82) <= 4; angryBirdLarge(26, 83) <= 4; angryBirdLarge(26, 84) <= 4; angryBirdLarge(26, 85) <= 4; angryBirdLarge(26, 86) <= 4; angryBirdLarge(26, 87) <= 4; angryBirdLarge(26, 88) <= 4; angryBirdLarge(26, 89) <= 4; angryBirdLarge(26, 90) <= 4; angryBirdLarge(26, 91) <= 4; angryBirdLarge(26, 92) <= 4; angryBirdLarge(26, 93) <= 4; angryBirdLarge(26, 94) <= 4; angryBirdLarge(26, 95) <= 4; angryBirdLarge(26, 96) <= 4; angryBirdLarge(26, 97) <= 4; angryBirdLarge(26, 98) <= 4; angryBirdLarge(26, 99) <= 4; angryBirdLarge(26, 100) <= 4; angryBirdLarge(26, 101) <= 4; angryBirdLarge(26, 102) <= 4; angryBirdLarge(26, 103) <= 4; angryBirdLarge(26, 104) <= 4; angryBirdLarge(26, 105) <= 4; angryBirdLarge(26, 106) <= 4; angryBirdLarge(26, 107) <= 4; angryBirdLarge(26, 108) <= 5; angryBirdLarge(26, 109) <= 5; angryBirdLarge(26, 110) <= 5; angryBirdLarge(26, 111) <= 5; angryBirdLarge(26, 112) <= 5; angryBirdLarge(26, 113) <= 5; angryBirdLarge(26, 114) <= 0; angryBirdLarge(26, 115) <= 0; angryBirdLarge(26, 116) <= 0; angryBirdLarge(26, 117) <= 0; angryBirdLarge(26, 118) <= 0; angryBirdLarge(26, 119) <= 0; angryBirdLarge(26, 120) <= 0; angryBirdLarge(26, 121) <= 0; angryBirdLarge(26, 122) <= 0; angryBirdLarge(26, 123) <= 0; angryBirdLarge(26, 124) <= 0; angryBirdLarge(26, 125) <= 0; angryBirdLarge(26, 126) <= 0; angryBirdLarge(26, 127) <= 0; angryBirdLarge(26, 128) <= 0; angryBirdLarge(26, 129) <= 0; angryBirdLarge(26, 130) <= 0; angryBirdLarge(26, 131) <= 0; angryBirdLarge(26, 132) <= 0; angryBirdLarge(26, 133) <= 0; angryBirdLarge(26, 134) <= 0; angryBirdLarge(26, 135) <= 0; angryBirdLarge(26, 136) <= 0; angryBirdLarge(26, 137) <= 0; angryBirdLarge(26, 138) <= 0; angryBirdLarge(26, 139) <= 0; angryBirdLarge(26, 140) <= 0; angryBirdLarge(26, 141) <= 0; angryBirdLarge(26, 142) <= 0; angryBirdLarge(26, 143) <= 0; angryBirdLarge(26, 144) <= 0; angryBirdLarge(26, 145) <= 0; angryBirdLarge(26, 146) <= 0; angryBirdLarge(26, 147) <= 0; angryBirdLarge(26, 148) <= 0; angryBirdLarge(26, 149) <= 0; 
angryBirdLarge(27, 0) <= 0; angryBirdLarge(27, 1) <= 0; angryBirdLarge(27, 2) <= 0; angryBirdLarge(27, 3) <= 0; angryBirdLarge(27, 4) <= 0; angryBirdLarge(27, 5) <= 0; angryBirdLarge(27, 6) <= 0; angryBirdLarge(27, 7) <= 0; angryBirdLarge(27, 8) <= 0; angryBirdLarge(27, 9) <= 0; angryBirdLarge(27, 10) <= 0; angryBirdLarge(27, 11) <= 0; angryBirdLarge(27, 12) <= 0; angryBirdLarge(27, 13) <= 0; angryBirdLarge(27, 14) <= 0; angryBirdLarge(27, 15) <= 0; angryBirdLarge(27, 16) <= 0; angryBirdLarge(27, 17) <= 0; angryBirdLarge(27, 18) <= 0; angryBirdLarge(27, 19) <= 0; angryBirdLarge(27, 20) <= 0; angryBirdLarge(27, 21) <= 0; angryBirdLarge(27, 22) <= 0; angryBirdLarge(27, 23) <= 0; angryBirdLarge(27, 24) <= 0; angryBirdLarge(27, 25) <= 0; angryBirdLarge(27, 26) <= 0; angryBirdLarge(27, 27) <= 0; angryBirdLarge(27, 28) <= 0; angryBirdLarge(27, 29) <= 0; angryBirdLarge(27, 30) <= 0; angryBirdLarge(27, 31) <= 0; angryBirdLarge(27, 32) <= 0; angryBirdLarge(27, 33) <= 0; angryBirdLarge(27, 34) <= 0; angryBirdLarge(27, 35) <= 0; angryBirdLarge(27, 36) <= 0; angryBirdLarge(27, 37) <= 0; angryBirdLarge(27, 38) <= 0; angryBirdLarge(27, 39) <= 0; angryBirdLarge(27, 40) <= 0; angryBirdLarge(27, 41) <= 0; angryBirdLarge(27, 42) <= 5; angryBirdLarge(27, 43) <= 5; angryBirdLarge(27, 44) <= 5; angryBirdLarge(27, 45) <= 5; angryBirdLarge(27, 46) <= 5; angryBirdLarge(27, 47) <= 5; angryBirdLarge(27, 48) <= 4; angryBirdLarge(27, 49) <= 4; angryBirdLarge(27, 50) <= 4; angryBirdLarge(27, 51) <= 4; angryBirdLarge(27, 52) <= 4; angryBirdLarge(27, 53) <= 4; angryBirdLarge(27, 54) <= 4; angryBirdLarge(27, 55) <= 4; angryBirdLarge(27, 56) <= 4; angryBirdLarge(27, 57) <= 4; angryBirdLarge(27, 58) <= 4; angryBirdLarge(27, 59) <= 4; angryBirdLarge(27, 60) <= 4; angryBirdLarge(27, 61) <= 4; angryBirdLarge(27, 62) <= 4; angryBirdLarge(27, 63) <= 4; angryBirdLarge(27, 64) <= 4; angryBirdLarge(27, 65) <= 4; angryBirdLarge(27, 66) <= 4; angryBirdLarge(27, 67) <= 4; angryBirdLarge(27, 68) <= 4; angryBirdLarge(27, 69) <= 4; angryBirdLarge(27, 70) <= 4; angryBirdLarge(27, 71) <= 4; angryBirdLarge(27, 72) <= 4; angryBirdLarge(27, 73) <= 4; angryBirdLarge(27, 74) <= 4; angryBirdLarge(27, 75) <= 4; angryBirdLarge(27, 76) <= 4; angryBirdLarge(27, 77) <= 4; angryBirdLarge(27, 78) <= 4; angryBirdLarge(27, 79) <= 4; angryBirdLarge(27, 80) <= 4; angryBirdLarge(27, 81) <= 4; angryBirdLarge(27, 82) <= 4; angryBirdLarge(27, 83) <= 4; angryBirdLarge(27, 84) <= 4; angryBirdLarge(27, 85) <= 4; angryBirdLarge(27, 86) <= 4; angryBirdLarge(27, 87) <= 4; angryBirdLarge(27, 88) <= 4; angryBirdLarge(27, 89) <= 4; angryBirdLarge(27, 90) <= 4; angryBirdLarge(27, 91) <= 4; angryBirdLarge(27, 92) <= 4; angryBirdLarge(27, 93) <= 4; angryBirdLarge(27, 94) <= 4; angryBirdLarge(27, 95) <= 4; angryBirdLarge(27, 96) <= 4; angryBirdLarge(27, 97) <= 4; angryBirdLarge(27, 98) <= 4; angryBirdLarge(27, 99) <= 4; angryBirdLarge(27, 100) <= 4; angryBirdLarge(27, 101) <= 4; angryBirdLarge(27, 102) <= 4; angryBirdLarge(27, 103) <= 4; angryBirdLarge(27, 104) <= 4; angryBirdLarge(27, 105) <= 4; angryBirdLarge(27, 106) <= 4; angryBirdLarge(27, 107) <= 4; angryBirdLarge(27, 108) <= 5; angryBirdLarge(27, 109) <= 5; angryBirdLarge(27, 110) <= 5; angryBirdLarge(27, 111) <= 5; angryBirdLarge(27, 112) <= 5; angryBirdLarge(27, 113) <= 5; angryBirdLarge(27, 114) <= 0; angryBirdLarge(27, 115) <= 0; angryBirdLarge(27, 116) <= 0; angryBirdLarge(27, 117) <= 0; angryBirdLarge(27, 118) <= 0; angryBirdLarge(27, 119) <= 0; angryBirdLarge(27, 120) <= 0; angryBirdLarge(27, 121) <= 0; angryBirdLarge(27, 122) <= 0; angryBirdLarge(27, 123) <= 0; angryBirdLarge(27, 124) <= 0; angryBirdLarge(27, 125) <= 0; angryBirdLarge(27, 126) <= 0; angryBirdLarge(27, 127) <= 0; angryBirdLarge(27, 128) <= 0; angryBirdLarge(27, 129) <= 0; angryBirdLarge(27, 130) <= 0; angryBirdLarge(27, 131) <= 0; angryBirdLarge(27, 132) <= 0; angryBirdLarge(27, 133) <= 0; angryBirdLarge(27, 134) <= 0; angryBirdLarge(27, 135) <= 0; angryBirdLarge(27, 136) <= 0; angryBirdLarge(27, 137) <= 0; angryBirdLarge(27, 138) <= 0; angryBirdLarge(27, 139) <= 0; angryBirdLarge(27, 140) <= 0; angryBirdLarge(27, 141) <= 0; angryBirdLarge(27, 142) <= 0; angryBirdLarge(27, 143) <= 0; angryBirdLarge(27, 144) <= 0; angryBirdLarge(27, 145) <= 0; angryBirdLarge(27, 146) <= 0; angryBirdLarge(27, 147) <= 0; angryBirdLarge(27, 148) <= 0; angryBirdLarge(27, 149) <= 0; 
angryBirdLarge(28, 0) <= 0; angryBirdLarge(28, 1) <= 0; angryBirdLarge(28, 2) <= 0; angryBirdLarge(28, 3) <= 0; angryBirdLarge(28, 4) <= 0; angryBirdLarge(28, 5) <= 0; angryBirdLarge(28, 6) <= 0; angryBirdLarge(28, 7) <= 0; angryBirdLarge(28, 8) <= 0; angryBirdLarge(28, 9) <= 0; angryBirdLarge(28, 10) <= 0; angryBirdLarge(28, 11) <= 0; angryBirdLarge(28, 12) <= 0; angryBirdLarge(28, 13) <= 0; angryBirdLarge(28, 14) <= 0; angryBirdLarge(28, 15) <= 0; angryBirdLarge(28, 16) <= 0; angryBirdLarge(28, 17) <= 0; angryBirdLarge(28, 18) <= 0; angryBirdLarge(28, 19) <= 0; angryBirdLarge(28, 20) <= 0; angryBirdLarge(28, 21) <= 0; angryBirdLarge(28, 22) <= 0; angryBirdLarge(28, 23) <= 0; angryBirdLarge(28, 24) <= 0; angryBirdLarge(28, 25) <= 0; angryBirdLarge(28, 26) <= 0; angryBirdLarge(28, 27) <= 0; angryBirdLarge(28, 28) <= 0; angryBirdLarge(28, 29) <= 0; angryBirdLarge(28, 30) <= 0; angryBirdLarge(28, 31) <= 0; angryBirdLarge(28, 32) <= 0; angryBirdLarge(28, 33) <= 0; angryBirdLarge(28, 34) <= 0; angryBirdLarge(28, 35) <= 0; angryBirdLarge(28, 36) <= 0; angryBirdLarge(28, 37) <= 0; angryBirdLarge(28, 38) <= 0; angryBirdLarge(28, 39) <= 0; angryBirdLarge(28, 40) <= 0; angryBirdLarge(28, 41) <= 0; angryBirdLarge(28, 42) <= 5; angryBirdLarge(28, 43) <= 5; angryBirdLarge(28, 44) <= 5; angryBirdLarge(28, 45) <= 5; angryBirdLarge(28, 46) <= 5; angryBirdLarge(28, 47) <= 5; angryBirdLarge(28, 48) <= 4; angryBirdLarge(28, 49) <= 4; angryBirdLarge(28, 50) <= 4; angryBirdLarge(28, 51) <= 4; angryBirdLarge(28, 52) <= 4; angryBirdLarge(28, 53) <= 4; angryBirdLarge(28, 54) <= 4; angryBirdLarge(28, 55) <= 4; angryBirdLarge(28, 56) <= 4; angryBirdLarge(28, 57) <= 4; angryBirdLarge(28, 58) <= 4; angryBirdLarge(28, 59) <= 4; angryBirdLarge(28, 60) <= 4; angryBirdLarge(28, 61) <= 4; angryBirdLarge(28, 62) <= 4; angryBirdLarge(28, 63) <= 4; angryBirdLarge(28, 64) <= 4; angryBirdLarge(28, 65) <= 4; angryBirdLarge(28, 66) <= 4; angryBirdLarge(28, 67) <= 4; angryBirdLarge(28, 68) <= 4; angryBirdLarge(28, 69) <= 4; angryBirdLarge(28, 70) <= 4; angryBirdLarge(28, 71) <= 4; angryBirdLarge(28, 72) <= 4; angryBirdLarge(28, 73) <= 4; angryBirdLarge(28, 74) <= 4; angryBirdLarge(28, 75) <= 4; angryBirdLarge(28, 76) <= 4; angryBirdLarge(28, 77) <= 4; angryBirdLarge(28, 78) <= 4; angryBirdLarge(28, 79) <= 4; angryBirdLarge(28, 80) <= 4; angryBirdLarge(28, 81) <= 4; angryBirdLarge(28, 82) <= 4; angryBirdLarge(28, 83) <= 4; angryBirdLarge(28, 84) <= 4; angryBirdLarge(28, 85) <= 4; angryBirdLarge(28, 86) <= 4; angryBirdLarge(28, 87) <= 4; angryBirdLarge(28, 88) <= 4; angryBirdLarge(28, 89) <= 4; angryBirdLarge(28, 90) <= 4; angryBirdLarge(28, 91) <= 4; angryBirdLarge(28, 92) <= 4; angryBirdLarge(28, 93) <= 4; angryBirdLarge(28, 94) <= 4; angryBirdLarge(28, 95) <= 4; angryBirdLarge(28, 96) <= 4; angryBirdLarge(28, 97) <= 4; angryBirdLarge(28, 98) <= 4; angryBirdLarge(28, 99) <= 4; angryBirdLarge(28, 100) <= 4; angryBirdLarge(28, 101) <= 4; angryBirdLarge(28, 102) <= 4; angryBirdLarge(28, 103) <= 4; angryBirdLarge(28, 104) <= 4; angryBirdLarge(28, 105) <= 4; angryBirdLarge(28, 106) <= 4; angryBirdLarge(28, 107) <= 4; angryBirdLarge(28, 108) <= 5; angryBirdLarge(28, 109) <= 5; angryBirdLarge(28, 110) <= 5; angryBirdLarge(28, 111) <= 5; angryBirdLarge(28, 112) <= 5; angryBirdLarge(28, 113) <= 5; angryBirdLarge(28, 114) <= 0; angryBirdLarge(28, 115) <= 0; angryBirdLarge(28, 116) <= 0; angryBirdLarge(28, 117) <= 0; angryBirdLarge(28, 118) <= 0; angryBirdLarge(28, 119) <= 0; angryBirdLarge(28, 120) <= 0; angryBirdLarge(28, 121) <= 0; angryBirdLarge(28, 122) <= 0; angryBirdLarge(28, 123) <= 0; angryBirdLarge(28, 124) <= 0; angryBirdLarge(28, 125) <= 0; angryBirdLarge(28, 126) <= 0; angryBirdLarge(28, 127) <= 0; angryBirdLarge(28, 128) <= 0; angryBirdLarge(28, 129) <= 0; angryBirdLarge(28, 130) <= 0; angryBirdLarge(28, 131) <= 0; angryBirdLarge(28, 132) <= 0; angryBirdLarge(28, 133) <= 0; angryBirdLarge(28, 134) <= 0; angryBirdLarge(28, 135) <= 0; angryBirdLarge(28, 136) <= 0; angryBirdLarge(28, 137) <= 0; angryBirdLarge(28, 138) <= 0; angryBirdLarge(28, 139) <= 0; angryBirdLarge(28, 140) <= 0; angryBirdLarge(28, 141) <= 0; angryBirdLarge(28, 142) <= 0; angryBirdLarge(28, 143) <= 0; angryBirdLarge(28, 144) <= 0; angryBirdLarge(28, 145) <= 0; angryBirdLarge(28, 146) <= 0; angryBirdLarge(28, 147) <= 0; angryBirdLarge(28, 148) <= 0; angryBirdLarge(28, 149) <= 0; 
angryBirdLarge(29, 0) <= 0; angryBirdLarge(29, 1) <= 0; angryBirdLarge(29, 2) <= 0; angryBirdLarge(29, 3) <= 0; angryBirdLarge(29, 4) <= 0; angryBirdLarge(29, 5) <= 0; angryBirdLarge(29, 6) <= 0; angryBirdLarge(29, 7) <= 0; angryBirdLarge(29, 8) <= 0; angryBirdLarge(29, 9) <= 0; angryBirdLarge(29, 10) <= 0; angryBirdLarge(29, 11) <= 0; angryBirdLarge(29, 12) <= 0; angryBirdLarge(29, 13) <= 0; angryBirdLarge(29, 14) <= 0; angryBirdLarge(29, 15) <= 0; angryBirdLarge(29, 16) <= 0; angryBirdLarge(29, 17) <= 0; angryBirdLarge(29, 18) <= 0; angryBirdLarge(29, 19) <= 0; angryBirdLarge(29, 20) <= 0; angryBirdLarge(29, 21) <= 0; angryBirdLarge(29, 22) <= 0; angryBirdLarge(29, 23) <= 0; angryBirdLarge(29, 24) <= 0; angryBirdLarge(29, 25) <= 0; angryBirdLarge(29, 26) <= 0; angryBirdLarge(29, 27) <= 0; angryBirdLarge(29, 28) <= 0; angryBirdLarge(29, 29) <= 0; angryBirdLarge(29, 30) <= 0; angryBirdLarge(29, 31) <= 0; angryBirdLarge(29, 32) <= 0; angryBirdLarge(29, 33) <= 0; angryBirdLarge(29, 34) <= 0; angryBirdLarge(29, 35) <= 0; angryBirdLarge(29, 36) <= 0; angryBirdLarge(29, 37) <= 0; angryBirdLarge(29, 38) <= 0; angryBirdLarge(29, 39) <= 0; angryBirdLarge(29, 40) <= 0; angryBirdLarge(29, 41) <= 0; angryBirdLarge(29, 42) <= 5; angryBirdLarge(29, 43) <= 5; angryBirdLarge(29, 44) <= 5; angryBirdLarge(29, 45) <= 5; angryBirdLarge(29, 46) <= 5; angryBirdLarge(29, 47) <= 5; angryBirdLarge(29, 48) <= 4; angryBirdLarge(29, 49) <= 4; angryBirdLarge(29, 50) <= 4; angryBirdLarge(29, 51) <= 4; angryBirdLarge(29, 52) <= 4; angryBirdLarge(29, 53) <= 4; angryBirdLarge(29, 54) <= 4; angryBirdLarge(29, 55) <= 4; angryBirdLarge(29, 56) <= 4; angryBirdLarge(29, 57) <= 4; angryBirdLarge(29, 58) <= 4; angryBirdLarge(29, 59) <= 4; angryBirdLarge(29, 60) <= 4; angryBirdLarge(29, 61) <= 4; angryBirdLarge(29, 62) <= 4; angryBirdLarge(29, 63) <= 4; angryBirdLarge(29, 64) <= 4; angryBirdLarge(29, 65) <= 4; angryBirdLarge(29, 66) <= 4; angryBirdLarge(29, 67) <= 4; angryBirdLarge(29, 68) <= 4; angryBirdLarge(29, 69) <= 4; angryBirdLarge(29, 70) <= 4; angryBirdLarge(29, 71) <= 4; angryBirdLarge(29, 72) <= 4; angryBirdLarge(29, 73) <= 4; angryBirdLarge(29, 74) <= 4; angryBirdLarge(29, 75) <= 4; angryBirdLarge(29, 76) <= 4; angryBirdLarge(29, 77) <= 4; angryBirdLarge(29, 78) <= 4; angryBirdLarge(29, 79) <= 4; angryBirdLarge(29, 80) <= 4; angryBirdLarge(29, 81) <= 4; angryBirdLarge(29, 82) <= 4; angryBirdLarge(29, 83) <= 4; angryBirdLarge(29, 84) <= 4; angryBirdLarge(29, 85) <= 4; angryBirdLarge(29, 86) <= 4; angryBirdLarge(29, 87) <= 4; angryBirdLarge(29, 88) <= 4; angryBirdLarge(29, 89) <= 4; angryBirdLarge(29, 90) <= 4; angryBirdLarge(29, 91) <= 4; angryBirdLarge(29, 92) <= 4; angryBirdLarge(29, 93) <= 4; angryBirdLarge(29, 94) <= 4; angryBirdLarge(29, 95) <= 4; angryBirdLarge(29, 96) <= 4; angryBirdLarge(29, 97) <= 4; angryBirdLarge(29, 98) <= 4; angryBirdLarge(29, 99) <= 4; angryBirdLarge(29, 100) <= 4; angryBirdLarge(29, 101) <= 4; angryBirdLarge(29, 102) <= 4; angryBirdLarge(29, 103) <= 4; angryBirdLarge(29, 104) <= 4; angryBirdLarge(29, 105) <= 4; angryBirdLarge(29, 106) <= 4; angryBirdLarge(29, 107) <= 4; angryBirdLarge(29, 108) <= 5; angryBirdLarge(29, 109) <= 5; angryBirdLarge(29, 110) <= 5; angryBirdLarge(29, 111) <= 5; angryBirdLarge(29, 112) <= 5; angryBirdLarge(29, 113) <= 5; angryBirdLarge(29, 114) <= 0; angryBirdLarge(29, 115) <= 0; angryBirdLarge(29, 116) <= 0; angryBirdLarge(29, 117) <= 0; angryBirdLarge(29, 118) <= 0; angryBirdLarge(29, 119) <= 0; angryBirdLarge(29, 120) <= 0; angryBirdLarge(29, 121) <= 0; angryBirdLarge(29, 122) <= 0; angryBirdLarge(29, 123) <= 0; angryBirdLarge(29, 124) <= 0; angryBirdLarge(29, 125) <= 0; angryBirdLarge(29, 126) <= 0; angryBirdLarge(29, 127) <= 0; angryBirdLarge(29, 128) <= 0; angryBirdLarge(29, 129) <= 0; angryBirdLarge(29, 130) <= 0; angryBirdLarge(29, 131) <= 0; angryBirdLarge(29, 132) <= 0; angryBirdLarge(29, 133) <= 0; angryBirdLarge(29, 134) <= 0; angryBirdLarge(29, 135) <= 0; angryBirdLarge(29, 136) <= 0; angryBirdLarge(29, 137) <= 0; angryBirdLarge(29, 138) <= 0; angryBirdLarge(29, 139) <= 0; angryBirdLarge(29, 140) <= 0; angryBirdLarge(29, 141) <= 0; angryBirdLarge(29, 142) <= 0; angryBirdLarge(29, 143) <= 0; angryBirdLarge(29, 144) <= 0; angryBirdLarge(29, 145) <= 0; angryBirdLarge(29, 146) <= 0; angryBirdLarge(29, 147) <= 0; angryBirdLarge(29, 148) <= 0; angryBirdLarge(29, 149) <= 0; 
angryBirdLarge(30, 0) <= 0; angryBirdLarge(30, 1) <= 0; angryBirdLarge(30, 2) <= 0; angryBirdLarge(30, 3) <= 0; angryBirdLarge(30, 4) <= 0; angryBirdLarge(30, 5) <= 0; angryBirdLarge(30, 6) <= 0; angryBirdLarge(30, 7) <= 0; angryBirdLarge(30, 8) <= 0; angryBirdLarge(30, 9) <= 0; angryBirdLarge(30, 10) <= 0; angryBirdLarge(30, 11) <= 0; angryBirdLarge(30, 12) <= 0; angryBirdLarge(30, 13) <= 0; angryBirdLarge(30, 14) <= 0; angryBirdLarge(30, 15) <= 0; angryBirdLarge(30, 16) <= 0; angryBirdLarge(30, 17) <= 0; angryBirdLarge(30, 18) <= 0; angryBirdLarge(30, 19) <= 0; angryBirdLarge(30, 20) <= 0; angryBirdLarge(30, 21) <= 0; angryBirdLarge(30, 22) <= 0; angryBirdLarge(30, 23) <= 0; angryBirdLarge(30, 24) <= 0; angryBirdLarge(30, 25) <= 0; angryBirdLarge(30, 26) <= 0; angryBirdLarge(30, 27) <= 0; angryBirdLarge(30, 28) <= 0; angryBirdLarge(30, 29) <= 0; angryBirdLarge(30, 30) <= 0; angryBirdLarge(30, 31) <= 0; angryBirdLarge(30, 32) <= 0; angryBirdLarge(30, 33) <= 0; angryBirdLarge(30, 34) <= 0; angryBirdLarge(30, 35) <= 0; angryBirdLarge(30, 36) <= 0; angryBirdLarge(30, 37) <= 0; angryBirdLarge(30, 38) <= 0; angryBirdLarge(30, 39) <= 0; angryBirdLarge(30, 40) <= 0; angryBirdLarge(30, 41) <= 0; angryBirdLarge(30, 42) <= 0; angryBirdLarge(30, 43) <= 0; angryBirdLarge(30, 44) <= 0; angryBirdLarge(30, 45) <= 0; angryBirdLarge(30, 46) <= 0; angryBirdLarge(30, 47) <= 0; angryBirdLarge(30, 48) <= 5; angryBirdLarge(30, 49) <= 5; angryBirdLarge(30, 50) <= 5; angryBirdLarge(30, 51) <= 5; angryBirdLarge(30, 52) <= 5; angryBirdLarge(30, 53) <= 5; angryBirdLarge(30, 54) <= 5; angryBirdLarge(30, 55) <= 5; angryBirdLarge(30, 56) <= 5; angryBirdLarge(30, 57) <= 5; angryBirdLarge(30, 58) <= 5; angryBirdLarge(30, 59) <= 5; angryBirdLarge(30, 60) <= 5; angryBirdLarge(30, 61) <= 5; angryBirdLarge(30, 62) <= 5; angryBirdLarge(30, 63) <= 5; angryBirdLarge(30, 64) <= 5; angryBirdLarge(30, 65) <= 5; angryBirdLarge(30, 66) <= 4; angryBirdLarge(30, 67) <= 4; angryBirdLarge(30, 68) <= 4; angryBirdLarge(30, 69) <= 4; angryBirdLarge(30, 70) <= 4; angryBirdLarge(30, 71) <= 4; angryBirdLarge(30, 72) <= 4; angryBirdLarge(30, 73) <= 4; angryBirdLarge(30, 74) <= 4; angryBirdLarge(30, 75) <= 4; angryBirdLarge(30, 76) <= 4; angryBirdLarge(30, 77) <= 4; angryBirdLarge(30, 78) <= 4; angryBirdLarge(30, 79) <= 4; angryBirdLarge(30, 80) <= 4; angryBirdLarge(30, 81) <= 4; angryBirdLarge(30, 82) <= 4; angryBirdLarge(30, 83) <= 4; angryBirdLarge(30, 84) <= 4; angryBirdLarge(30, 85) <= 4; angryBirdLarge(30, 86) <= 4; angryBirdLarge(30, 87) <= 4; angryBirdLarge(30, 88) <= 4; angryBirdLarge(30, 89) <= 4; angryBirdLarge(30, 90) <= 4; angryBirdLarge(30, 91) <= 4; angryBirdLarge(30, 92) <= 4; angryBirdLarge(30, 93) <= 4; angryBirdLarge(30, 94) <= 4; angryBirdLarge(30, 95) <= 4; angryBirdLarge(30, 96) <= 4; angryBirdLarge(30, 97) <= 4; angryBirdLarge(30, 98) <= 4; angryBirdLarge(30, 99) <= 4; angryBirdLarge(30, 100) <= 4; angryBirdLarge(30, 101) <= 4; angryBirdLarge(30, 102) <= 4; angryBirdLarge(30, 103) <= 4; angryBirdLarge(30, 104) <= 4; angryBirdLarge(30, 105) <= 4; angryBirdLarge(30, 106) <= 4; angryBirdLarge(30, 107) <= 4; angryBirdLarge(30, 108) <= 4; angryBirdLarge(30, 109) <= 4; angryBirdLarge(30, 110) <= 4; angryBirdLarge(30, 111) <= 4; angryBirdLarge(30, 112) <= 4; angryBirdLarge(30, 113) <= 4; angryBirdLarge(30, 114) <= 5; angryBirdLarge(30, 115) <= 5; angryBirdLarge(30, 116) <= 5; angryBirdLarge(30, 117) <= 5; angryBirdLarge(30, 118) <= 5; angryBirdLarge(30, 119) <= 5; angryBirdLarge(30, 120) <= 0; angryBirdLarge(30, 121) <= 0; angryBirdLarge(30, 122) <= 0; angryBirdLarge(30, 123) <= 0; angryBirdLarge(30, 124) <= 0; angryBirdLarge(30, 125) <= 0; angryBirdLarge(30, 126) <= 0; angryBirdLarge(30, 127) <= 0; angryBirdLarge(30, 128) <= 0; angryBirdLarge(30, 129) <= 0; angryBirdLarge(30, 130) <= 0; angryBirdLarge(30, 131) <= 0; angryBirdLarge(30, 132) <= 0; angryBirdLarge(30, 133) <= 0; angryBirdLarge(30, 134) <= 0; angryBirdLarge(30, 135) <= 0; angryBirdLarge(30, 136) <= 0; angryBirdLarge(30, 137) <= 0; angryBirdLarge(30, 138) <= 0; angryBirdLarge(30, 139) <= 0; angryBirdLarge(30, 140) <= 0; angryBirdLarge(30, 141) <= 0; angryBirdLarge(30, 142) <= 0; angryBirdLarge(30, 143) <= 0; angryBirdLarge(30, 144) <= 0; angryBirdLarge(30, 145) <= 0; angryBirdLarge(30, 146) <= 0; angryBirdLarge(30, 147) <= 0; angryBirdLarge(30, 148) <= 0; angryBirdLarge(30, 149) <= 0; 
angryBirdLarge(31, 0) <= 0; angryBirdLarge(31, 1) <= 0; angryBirdLarge(31, 2) <= 0; angryBirdLarge(31, 3) <= 0; angryBirdLarge(31, 4) <= 0; angryBirdLarge(31, 5) <= 0; angryBirdLarge(31, 6) <= 0; angryBirdLarge(31, 7) <= 0; angryBirdLarge(31, 8) <= 0; angryBirdLarge(31, 9) <= 0; angryBirdLarge(31, 10) <= 0; angryBirdLarge(31, 11) <= 0; angryBirdLarge(31, 12) <= 0; angryBirdLarge(31, 13) <= 0; angryBirdLarge(31, 14) <= 0; angryBirdLarge(31, 15) <= 0; angryBirdLarge(31, 16) <= 0; angryBirdLarge(31, 17) <= 0; angryBirdLarge(31, 18) <= 0; angryBirdLarge(31, 19) <= 0; angryBirdLarge(31, 20) <= 0; angryBirdLarge(31, 21) <= 0; angryBirdLarge(31, 22) <= 0; angryBirdLarge(31, 23) <= 0; angryBirdLarge(31, 24) <= 0; angryBirdLarge(31, 25) <= 0; angryBirdLarge(31, 26) <= 0; angryBirdLarge(31, 27) <= 0; angryBirdLarge(31, 28) <= 0; angryBirdLarge(31, 29) <= 0; angryBirdLarge(31, 30) <= 0; angryBirdLarge(31, 31) <= 0; angryBirdLarge(31, 32) <= 0; angryBirdLarge(31, 33) <= 0; angryBirdLarge(31, 34) <= 0; angryBirdLarge(31, 35) <= 0; angryBirdLarge(31, 36) <= 0; angryBirdLarge(31, 37) <= 0; angryBirdLarge(31, 38) <= 0; angryBirdLarge(31, 39) <= 0; angryBirdLarge(31, 40) <= 0; angryBirdLarge(31, 41) <= 0; angryBirdLarge(31, 42) <= 0; angryBirdLarge(31, 43) <= 0; angryBirdLarge(31, 44) <= 0; angryBirdLarge(31, 45) <= 0; angryBirdLarge(31, 46) <= 0; angryBirdLarge(31, 47) <= 0; angryBirdLarge(31, 48) <= 5; angryBirdLarge(31, 49) <= 5; angryBirdLarge(31, 50) <= 5; angryBirdLarge(31, 51) <= 5; angryBirdLarge(31, 52) <= 5; angryBirdLarge(31, 53) <= 5; angryBirdLarge(31, 54) <= 5; angryBirdLarge(31, 55) <= 5; angryBirdLarge(31, 56) <= 5; angryBirdLarge(31, 57) <= 5; angryBirdLarge(31, 58) <= 5; angryBirdLarge(31, 59) <= 5; angryBirdLarge(31, 60) <= 5; angryBirdLarge(31, 61) <= 5; angryBirdLarge(31, 62) <= 5; angryBirdLarge(31, 63) <= 5; angryBirdLarge(31, 64) <= 5; angryBirdLarge(31, 65) <= 5; angryBirdLarge(31, 66) <= 4; angryBirdLarge(31, 67) <= 4; angryBirdLarge(31, 68) <= 4; angryBirdLarge(31, 69) <= 4; angryBirdLarge(31, 70) <= 4; angryBirdLarge(31, 71) <= 4; angryBirdLarge(31, 72) <= 4; angryBirdLarge(31, 73) <= 4; angryBirdLarge(31, 74) <= 4; angryBirdLarge(31, 75) <= 4; angryBirdLarge(31, 76) <= 4; angryBirdLarge(31, 77) <= 4; angryBirdLarge(31, 78) <= 4; angryBirdLarge(31, 79) <= 4; angryBirdLarge(31, 80) <= 4; angryBirdLarge(31, 81) <= 4; angryBirdLarge(31, 82) <= 4; angryBirdLarge(31, 83) <= 4; angryBirdLarge(31, 84) <= 4; angryBirdLarge(31, 85) <= 4; angryBirdLarge(31, 86) <= 4; angryBirdLarge(31, 87) <= 4; angryBirdLarge(31, 88) <= 4; angryBirdLarge(31, 89) <= 4; angryBirdLarge(31, 90) <= 4; angryBirdLarge(31, 91) <= 4; angryBirdLarge(31, 92) <= 4; angryBirdLarge(31, 93) <= 4; angryBirdLarge(31, 94) <= 4; angryBirdLarge(31, 95) <= 4; angryBirdLarge(31, 96) <= 4; angryBirdLarge(31, 97) <= 4; angryBirdLarge(31, 98) <= 4; angryBirdLarge(31, 99) <= 4; angryBirdLarge(31, 100) <= 4; angryBirdLarge(31, 101) <= 4; angryBirdLarge(31, 102) <= 4; angryBirdLarge(31, 103) <= 4; angryBirdLarge(31, 104) <= 4; angryBirdLarge(31, 105) <= 4; angryBirdLarge(31, 106) <= 4; angryBirdLarge(31, 107) <= 4; angryBirdLarge(31, 108) <= 4; angryBirdLarge(31, 109) <= 4; angryBirdLarge(31, 110) <= 4; angryBirdLarge(31, 111) <= 4; angryBirdLarge(31, 112) <= 4; angryBirdLarge(31, 113) <= 4; angryBirdLarge(31, 114) <= 5; angryBirdLarge(31, 115) <= 5; angryBirdLarge(31, 116) <= 5; angryBirdLarge(31, 117) <= 5; angryBirdLarge(31, 118) <= 5; angryBirdLarge(31, 119) <= 5; angryBirdLarge(31, 120) <= 0; angryBirdLarge(31, 121) <= 0; angryBirdLarge(31, 122) <= 0; angryBirdLarge(31, 123) <= 0; angryBirdLarge(31, 124) <= 0; angryBirdLarge(31, 125) <= 0; angryBirdLarge(31, 126) <= 0; angryBirdLarge(31, 127) <= 0; angryBirdLarge(31, 128) <= 0; angryBirdLarge(31, 129) <= 0; angryBirdLarge(31, 130) <= 0; angryBirdLarge(31, 131) <= 0; angryBirdLarge(31, 132) <= 0; angryBirdLarge(31, 133) <= 0; angryBirdLarge(31, 134) <= 0; angryBirdLarge(31, 135) <= 0; angryBirdLarge(31, 136) <= 0; angryBirdLarge(31, 137) <= 0; angryBirdLarge(31, 138) <= 0; angryBirdLarge(31, 139) <= 0; angryBirdLarge(31, 140) <= 0; angryBirdLarge(31, 141) <= 0; angryBirdLarge(31, 142) <= 0; angryBirdLarge(31, 143) <= 0; angryBirdLarge(31, 144) <= 0; angryBirdLarge(31, 145) <= 0; angryBirdLarge(31, 146) <= 0; angryBirdLarge(31, 147) <= 0; angryBirdLarge(31, 148) <= 0; angryBirdLarge(31, 149) <= 0; 
angryBirdLarge(32, 0) <= 0; angryBirdLarge(32, 1) <= 0; angryBirdLarge(32, 2) <= 0; angryBirdLarge(32, 3) <= 0; angryBirdLarge(32, 4) <= 0; angryBirdLarge(32, 5) <= 0; angryBirdLarge(32, 6) <= 0; angryBirdLarge(32, 7) <= 0; angryBirdLarge(32, 8) <= 0; angryBirdLarge(32, 9) <= 0; angryBirdLarge(32, 10) <= 0; angryBirdLarge(32, 11) <= 0; angryBirdLarge(32, 12) <= 0; angryBirdLarge(32, 13) <= 0; angryBirdLarge(32, 14) <= 0; angryBirdLarge(32, 15) <= 0; angryBirdLarge(32, 16) <= 0; angryBirdLarge(32, 17) <= 0; angryBirdLarge(32, 18) <= 0; angryBirdLarge(32, 19) <= 0; angryBirdLarge(32, 20) <= 0; angryBirdLarge(32, 21) <= 0; angryBirdLarge(32, 22) <= 0; angryBirdLarge(32, 23) <= 0; angryBirdLarge(32, 24) <= 0; angryBirdLarge(32, 25) <= 0; angryBirdLarge(32, 26) <= 0; angryBirdLarge(32, 27) <= 0; angryBirdLarge(32, 28) <= 0; angryBirdLarge(32, 29) <= 0; angryBirdLarge(32, 30) <= 0; angryBirdLarge(32, 31) <= 0; angryBirdLarge(32, 32) <= 0; angryBirdLarge(32, 33) <= 0; angryBirdLarge(32, 34) <= 0; angryBirdLarge(32, 35) <= 0; angryBirdLarge(32, 36) <= 0; angryBirdLarge(32, 37) <= 0; angryBirdLarge(32, 38) <= 0; angryBirdLarge(32, 39) <= 0; angryBirdLarge(32, 40) <= 0; angryBirdLarge(32, 41) <= 0; angryBirdLarge(32, 42) <= 0; angryBirdLarge(32, 43) <= 0; angryBirdLarge(32, 44) <= 0; angryBirdLarge(32, 45) <= 0; angryBirdLarge(32, 46) <= 0; angryBirdLarge(32, 47) <= 0; angryBirdLarge(32, 48) <= 5; angryBirdLarge(32, 49) <= 5; angryBirdLarge(32, 50) <= 5; angryBirdLarge(32, 51) <= 5; angryBirdLarge(32, 52) <= 5; angryBirdLarge(32, 53) <= 5; angryBirdLarge(32, 54) <= 5; angryBirdLarge(32, 55) <= 5; angryBirdLarge(32, 56) <= 5; angryBirdLarge(32, 57) <= 5; angryBirdLarge(32, 58) <= 5; angryBirdLarge(32, 59) <= 5; angryBirdLarge(32, 60) <= 5; angryBirdLarge(32, 61) <= 5; angryBirdLarge(32, 62) <= 5; angryBirdLarge(32, 63) <= 5; angryBirdLarge(32, 64) <= 5; angryBirdLarge(32, 65) <= 5; angryBirdLarge(32, 66) <= 4; angryBirdLarge(32, 67) <= 4; angryBirdLarge(32, 68) <= 4; angryBirdLarge(32, 69) <= 4; angryBirdLarge(32, 70) <= 4; angryBirdLarge(32, 71) <= 4; angryBirdLarge(32, 72) <= 4; angryBirdLarge(32, 73) <= 4; angryBirdLarge(32, 74) <= 4; angryBirdLarge(32, 75) <= 4; angryBirdLarge(32, 76) <= 4; angryBirdLarge(32, 77) <= 4; angryBirdLarge(32, 78) <= 4; angryBirdLarge(32, 79) <= 4; angryBirdLarge(32, 80) <= 4; angryBirdLarge(32, 81) <= 4; angryBirdLarge(32, 82) <= 4; angryBirdLarge(32, 83) <= 4; angryBirdLarge(32, 84) <= 4; angryBirdLarge(32, 85) <= 4; angryBirdLarge(32, 86) <= 4; angryBirdLarge(32, 87) <= 4; angryBirdLarge(32, 88) <= 4; angryBirdLarge(32, 89) <= 4; angryBirdLarge(32, 90) <= 4; angryBirdLarge(32, 91) <= 4; angryBirdLarge(32, 92) <= 4; angryBirdLarge(32, 93) <= 4; angryBirdLarge(32, 94) <= 4; angryBirdLarge(32, 95) <= 4; angryBirdLarge(32, 96) <= 4; angryBirdLarge(32, 97) <= 4; angryBirdLarge(32, 98) <= 4; angryBirdLarge(32, 99) <= 4; angryBirdLarge(32, 100) <= 4; angryBirdLarge(32, 101) <= 4; angryBirdLarge(32, 102) <= 4; angryBirdLarge(32, 103) <= 4; angryBirdLarge(32, 104) <= 4; angryBirdLarge(32, 105) <= 4; angryBirdLarge(32, 106) <= 4; angryBirdLarge(32, 107) <= 4; angryBirdLarge(32, 108) <= 4; angryBirdLarge(32, 109) <= 4; angryBirdLarge(32, 110) <= 4; angryBirdLarge(32, 111) <= 4; angryBirdLarge(32, 112) <= 4; angryBirdLarge(32, 113) <= 4; angryBirdLarge(32, 114) <= 5; angryBirdLarge(32, 115) <= 5; angryBirdLarge(32, 116) <= 5; angryBirdLarge(32, 117) <= 5; angryBirdLarge(32, 118) <= 5; angryBirdLarge(32, 119) <= 5; angryBirdLarge(32, 120) <= 0; angryBirdLarge(32, 121) <= 0; angryBirdLarge(32, 122) <= 0; angryBirdLarge(32, 123) <= 0; angryBirdLarge(32, 124) <= 0; angryBirdLarge(32, 125) <= 0; angryBirdLarge(32, 126) <= 0; angryBirdLarge(32, 127) <= 0; angryBirdLarge(32, 128) <= 0; angryBirdLarge(32, 129) <= 0; angryBirdLarge(32, 130) <= 0; angryBirdLarge(32, 131) <= 0; angryBirdLarge(32, 132) <= 0; angryBirdLarge(32, 133) <= 0; angryBirdLarge(32, 134) <= 0; angryBirdLarge(32, 135) <= 0; angryBirdLarge(32, 136) <= 0; angryBirdLarge(32, 137) <= 0; angryBirdLarge(32, 138) <= 0; angryBirdLarge(32, 139) <= 0; angryBirdLarge(32, 140) <= 0; angryBirdLarge(32, 141) <= 0; angryBirdLarge(32, 142) <= 0; angryBirdLarge(32, 143) <= 0; angryBirdLarge(32, 144) <= 0; angryBirdLarge(32, 145) <= 0; angryBirdLarge(32, 146) <= 0; angryBirdLarge(32, 147) <= 0; angryBirdLarge(32, 148) <= 0; angryBirdLarge(32, 149) <= 0; 
angryBirdLarge(33, 0) <= 0; angryBirdLarge(33, 1) <= 0; angryBirdLarge(33, 2) <= 0; angryBirdLarge(33, 3) <= 0; angryBirdLarge(33, 4) <= 0; angryBirdLarge(33, 5) <= 0; angryBirdLarge(33, 6) <= 0; angryBirdLarge(33, 7) <= 0; angryBirdLarge(33, 8) <= 0; angryBirdLarge(33, 9) <= 0; angryBirdLarge(33, 10) <= 0; angryBirdLarge(33, 11) <= 0; angryBirdLarge(33, 12) <= 0; angryBirdLarge(33, 13) <= 0; angryBirdLarge(33, 14) <= 0; angryBirdLarge(33, 15) <= 0; angryBirdLarge(33, 16) <= 0; angryBirdLarge(33, 17) <= 0; angryBirdLarge(33, 18) <= 0; angryBirdLarge(33, 19) <= 0; angryBirdLarge(33, 20) <= 0; angryBirdLarge(33, 21) <= 0; angryBirdLarge(33, 22) <= 0; angryBirdLarge(33, 23) <= 0; angryBirdLarge(33, 24) <= 0; angryBirdLarge(33, 25) <= 0; angryBirdLarge(33, 26) <= 0; angryBirdLarge(33, 27) <= 0; angryBirdLarge(33, 28) <= 0; angryBirdLarge(33, 29) <= 0; angryBirdLarge(33, 30) <= 0; angryBirdLarge(33, 31) <= 0; angryBirdLarge(33, 32) <= 0; angryBirdLarge(33, 33) <= 0; angryBirdLarge(33, 34) <= 0; angryBirdLarge(33, 35) <= 0; angryBirdLarge(33, 36) <= 0; angryBirdLarge(33, 37) <= 0; angryBirdLarge(33, 38) <= 0; angryBirdLarge(33, 39) <= 0; angryBirdLarge(33, 40) <= 0; angryBirdLarge(33, 41) <= 0; angryBirdLarge(33, 42) <= 0; angryBirdLarge(33, 43) <= 0; angryBirdLarge(33, 44) <= 0; angryBirdLarge(33, 45) <= 0; angryBirdLarge(33, 46) <= 0; angryBirdLarge(33, 47) <= 0; angryBirdLarge(33, 48) <= 5; angryBirdLarge(33, 49) <= 5; angryBirdLarge(33, 50) <= 5; angryBirdLarge(33, 51) <= 5; angryBirdLarge(33, 52) <= 5; angryBirdLarge(33, 53) <= 5; angryBirdLarge(33, 54) <= 5; angryBirdLarge(33, 55) <= 5; angryBirdLarge(33, 56) <= 5; angryBirdLarge(33, 57) <= 5; angryBirdLarge(33, 58) <= 5; angryBirdLarge(33, 59) <= 5; angryBirdLarge(33, 60) <= 5; angryBirdLarge(33, 61) <= 5; angryBirdLarge(33, 62) <= 5; angryBirdLarge(33, 63) <= 5; angryBirdLarge(33, 64) <= 5; angryBirdLarge(33, 65) <= 5; angryBirdLarge(33, 66) <= 4; angryBirdLarge(33, 67) <= 4; angryBirdLarge(33, 68) <= 4; angryBirdLarge(33, 69) <= 4; angryBirdLarge(33, 70) <= 4; angryBirdLarge(33, 71) <= 4; angryBirdLarge(33, 72) <= 4; angryBirdLarge(33, 73) <= 4; angryBirdLarge(33, 74) <= 4; angryBirdLarge(33, 75) <= 4; angryBirdLarge(33, 76) <= 4; angryBirdLarge(33, 77) <= 4; angryBirdLarge(33, 78) <= 4; angryBirdLarge(33, 79) <= 4; angryBirdLarge(33, 80) <= 4; angryBirdLarge(33, 81) <= 4; angryBirdLarge(33, 82) <= 4; angryBirdLarge(33, 83) <= 4; angryBirdLarge(33, 84) <= 4; angryBirdLarge(33, 85) <= 4; angryBirdLarge(33, 86) <= 4; angryBirdLarge(33, 87) <= 4; angryBirdLarge(33, 88) <= 4; angryBirdLarge(33, 89) <= 4; angryBirdLarge(33, 90) <= 4; angryBirdLarge(33, 91) <= 4; angryBirdLarge(33, 92) <= 4; angryBirdLarge(33, 93) <= 4; angryBirdLarge(33, 94) <= 4; angryBirdLarge(33, 95) <= 4; angryBirdLarge(33, 96) <= 4; angryBirdLarge(33, 97) <= 4; angryBirdLarge(33, 98) <= 4; angryBirdLarge(33, 99) <= 4; angryBirdLarge(33, 100) <= 4; angryBirdLarge(33, 101) <= 4; angryBirdLarge(33, 102) <= 4; angryBirdLarge(33, 103) <= 4; angryBirdLarge(33, 104) <= 4; angryBirdLarge(33, 105) <= 4; angryBirdLarge(33, 106) <= 4; angryBirdLarge(33, 107) <= 4; angryBirdLarge(33, 108) <= 4; angryBirdLarge(33, 109) <= 4; angryBirdLarge(33, 110) <= 4; angryBirdLarge(33, 111) <= 4; angryBirdLarge(33, 112) <= 4; angryBirdLarge(33, 113) <= 4; angryBirdLarge(33, 114) <= 5; angryBirdLarge(33, 115) <= 5; angryBirdLarge(33, 116) <= 5; angryBirdLarge(33, 117) <= 5; angryBirdLarge(33, 118) <= 5; angryBirdLarge(33, 119) <= 5; angryBirdLarge(33, 120) <= 0; angryBirdLarge(33, 121) <= 0; angryBirdLarge(33, 122) <= 0; angryBirdLarge(33, 123) <= 0; angryBirdLarge(33, 124) <= 0; angryBirdLarge(33, 125) <= 0; angryBirdLarge(33, 126) <= 0; angryBirdLarge(33, 127) <= 0; angryBirdLarge(33, 128) <= 0; angryBirdLarge(33, 129) <= 0; angryBirdLarge(33, 130) <= 0; angryBirdLarge(33, 131) <= 0; angryBirdLarge(33, 132) <= 0; angryBirdLarge(33, 133) <= 0; angryBirdLarge(33, 134) <= 0; angryBirdLarge(33, 135) <= 0; angryBirdLarge(33, 136) <= 0; angryBirdLarge(33, 137) <= 0; angryBirdLarge(33, 138) <= 0; angryBirdLarge(33, 139) <= 0; angryBirdLarge(33, 140) <= 0; angryBirdLarge(33, 141) <= 0; angryBirdLarge(33, 142) <= 0; angryBirdLarge(33, 143) <= 0; angryBirdLarge(33, 144) <= 0; angryBirdLarge(33, 145) <= 0; angryBirdLarge(33, 146) <= 0; angryBirdLarge(33, 147) <= 0; angryBirdLarge(33, 148) <= 0; angryBirdLarge(33, 149) <= 0; 
angryBirdLarge(34, 0) <= 0; angryBirdLarge(34, 1) <= 0; angryBirdLarge(34, 2) <= 0; angryBirdLarge(34, 3) <= 0; angryBirdLarge(34, 4) <= 0; angryBirdLarge(34, 5) <= 0; angryBirdLarge(34, 6) <= 0; angryBirdLarge(34, 7) <= 0; angryBirdLarge(34, 8) <= 0; angryBirdLarge(34, 9) <= 0; angryBirdLarge(34, 10) <= 0; angryBirdLarge(34, 11) <= 0; angryBirdLarge(34, 12) <= 0; angryBirdLarge(34, 13) <= 0; angryBirdLarge(34, 14) <= 0; angryBirdLarge(34, 15) <= 0; angryBirdLarge(34, 16) <= 0; angryBirdLarge(34, 17) <= 0; angryBirdLarge(34, 18) <= 0; angryBirdLarge(34, 19) <= 0; angryBirdLarge(34, 20) <= 0; angryBirdLarge(34, 21) <= 0; angryBirdLarge(34, 22) <= 0; angryBirdLarge(34, 23) <= 0; angryBirdLarge(34, 24) <= 0; angryBirdLarge(34, 25) <= 0; angryBirdLarge(34, 26) <= 0; angryBirdLarge(34, 27) <= 0; angryBirdLarge(34, 28) <= 0; angryBirdLarge(34, 29) <= 0; angryBirdLarge(34, 30) <= 0; angryBirdLarge(34, 31) <= 0; angryBirdLarge(34, 32) <= 0; angryBirdLarge(34, 33) <= 0; angryBirdLarge(34, 34) <= 0; angryBirdLarge(34, 35) <= 0; angryBirdLarge(34, 36) <= 0; angryBirdLarge(34, 37) <= 0; angryBirdLarge(34, 38) <= 0; angryBirdLarge(34, 39) <= 0; angryBirdLarge(34, 40) <= 0; angryBirdLarge(34, 41) <= 0; angryBirdLarge(34, 42) <= 0; angryBirdLarge(34, 43) <= 0; angryBirdLarge(34, 44) <= 0; angryBirdLarge(34, 45) <= 0; angryBirdLarge(34, 46) <= 0; angryBirdLarge(34, 47) <= 0; angryBirdLarge(34, 48) <= 5; angryBirdLarge(34, 49) <= 5; angryBirdLarge(34, 50) <= 5; angryBirdLarge(34, 51) <= 5; angryBirdLarge(34, 52) <= 5; angryBirdLarge(34, 53) <= 5; angryBirdLarge(34, 54) <= 5; angryBirdLarge(34, 55) <= 5; angryBirdLarge(34, 56) <= 5; angryBirdLarge(34, 57) <= 5; angryBirdLarge(34, 58) <= 5; angryBirdLarge(34, 59) <= 5; angryBirdLarge(34, 60) <= 5; angryBirdLarge(34, 61) <= 5; angryBirdLarge(34, 62) <= 5; angryBirdLarge(34, 63) <= 5; angryBirdLarge(34, 64) <= 5; angryBirdLarge(34, 65) <= 5; angryBirdLarge(34, 66) <= 4; angryBirdLarge(34, 67) <= 4; angryBirdLarge(34, 68) <= 4; angryBirdLarge(34, 69) <= 4; angryBirdLarge(34, 70) <= 4; angryBirdLarge(34, 71) <= 4; angryBirdLarge(34, 72) <= 4; angryBirdLarge(34, 73) <= 4; angryBirdLarge(34, 74) <= 4; angryBirdLarge(34, 75) <= 4; angryBirdLarge(34, 76) <= 4; angryBirdLarge(34, 77) <= 4; angryBirdLarge(34, 78) <= 4; angryBirdLarge(34, 79) <= 4; angryBirdLarge(34, 80) <= 4; angryBirdLarge(34, 81) <= 4; angryBirdLarge(34, 82) <= 4; angryBirdLarge(34, 83) <= 4; angryBirdLarge(34, 84) <= 4; angryBirdLarge(34, 85) <= 4; angryBirdLarge(34, 86) <= 4; angryBirdLarge(34, 87) <= 4; angryBirdLarge(34, 88) <= 4; angryBirdLarge(34, 89) <= 4; angryBirdLarge(34, 90) <= 4; angryBirdLarge(34, 91) <= 4; angryBirdLarge(34, 92) <= 4; angryBirdLarge(34, 93) <= 4; angryBirdLarge(34, 94) <= 4; angryBirdLarge(34, 95) <= 4; angryBirdLarge(34, 96) <= 4; angryBirdLarge(34, 97) <= 4; angryBirdLarge(34, 98) <= 4; angryBirdLarge(34, 99) <= 4; angryBirdLarge(34, 100) <= 4; angryBirdLarge(34, 101) <= 4; angryBirdLarge(34, 102) <= 4; angryBirdLarge(34, 103) <= 4; angryBirdLarge(34, 104) <= 4; angryBirdLarge(34, 105) <= 4; angryBirdLarge(34, 106) <= 4; angryBirdLarge(34, 107) <= 4; angryBirdLarge(34, 108) <= 4; angryBirdLarge(34, 109) <= 4; angryBirdLarge(34, 110) <= 4; angryBirdLarge(34, 111) <= 4; angryBirdLarge(34, 112) <= 4; angryBirdLarge(34, 113) <= 4; angryBirdLarge(34, 114) <= 5; angryBirdLarge(34, 115) <= 5; angryBirdLarge(34, 116) <= 5; angryBirdLarge(34, 117) <= 5; angryBirdLarge(34, 118) <= 5; angryBirdLarge(34, 119) <= 5; angryBirdLarge(34, 120) <= 0; angryBirdLarge(34, 121) <= 0; angryBirdLarge(34, 122) <= 0; angryBirdLarge(34, 123) <= 0; angryBirdLarge(34, 124) <= 0; angryBirdLarge(34, 125) <= 0; angryBirdLarge(34, 126) <= 0; angryBirdLarge(34, 127) <= 0; angryBirdLarge(34, 128) <= 0; angryBirdLarge(34, 129) <= 0; angryBirdLarge(34, 130) <= 0; angryBirdLarge(34, 131) <= 0; angryBirdLarge(34, 132) <= 0; angryBirdLarge(34, 133) <= 0; angryBirdLarge(34, 134) <= 0; angryBirdLarge(34, 135) <= 0; angryBirdLarge(34, 136) <= 0; angryBirdLarge(34, 137) <= 0; angryBirdLarge(34, 138) <= 0; angryBirdLarge(34, 139) <= 0; angryBirdLarge(34, 140) <= 0; angryBirdLarge(34, 141) <= 0; angryBirdLarge(34, 142) <= 0; angryBirdLarge(34, 143) <= 0; angryBirdLarge(34, 144) <= 0; angryBirdLarge(34, 145) <= 0; angryBirdLarge(34, 146) <= 0; angryBirdLarge(34, 147) <= 0; angryBirdLarge(34, 148) <= 0; angryBirdLarge(34, 149) <= 0; 
angryBirdLarge(35, 0) <= 0; angryBirdLarge(35, 1) <= 0; angryBirdLarge(35, 2) <= 0; angryBirdLarge(35, 3) <= 0; angryBirdLarge(35, 4) <= 0; angryBirdLarge(35, 5) <= 0; angryBirdLarge(35, 6) <= 0; angryBirdLarge(35, 7) <= 0; angryBirdLarge(35, 8) <= 0; angryBirdLarge(35, 9) <= 0; angryBirdLarge(35, 10) <= 0; angryBirdLarge(35, 11) <= 0; angryBirdLarge(35, 12) <= 0; angryBirdLarge(35, 13) <= 0; angryBirdLarge(35, 14) <= 0; angryBirdLarge(35, 15) <= 0; angryBirdLarge(35, 16) <= 0; angryBirdLarge(35, 17) <= 0; angryBirdLarge(35, 18) <= 0; angryBirdLarge(35, 19) <= 0; angryBirdLarge(35, 20) <= 0; angryBirdLarge(35, 21) <= 0; angryBirdLarge(35, 22) <= 0; angryBirdLarge(35, 23) <= 0; angryBirdLarge(35, 24) <= 0; angryBirdLarge(35, 25) <= 0; angryBirdLarge(35, 26) <= 0; angryBirdLarge(35, 27) <= 0; angryBirdLarge(35, 28) <= 0; angryBirdLarge(35, 29) <= 0; angryBirdLarge(35, 30) <= 0; angryBirdLarge(35, 31) <= 0; angryBirdLarge(35, 32) <= 0; angryBirdLarge(35, 33) <= 0; angryBirdLarge(35, 34) <= 0; angryBirdLarge(35, 35) <= 0; angryBirdLarge(35, 36) <= 0; angryBirdLarge(35, 37) <= 0; angryBirdLarge(35, 38) <= 0; angryBirdLarge(35, 39) <= 0; angryBirdLarge(35, 40) <= 0; angryBirdLarge(35, 41) <= 0; angryBirdLarge(35, 42) <= 0; angryBirdLarge(35, 43) <= 0; angryBirdLarge(35, 44) <= 0; angryBirdLarge(35, 45) <= 0; angryBirdLarge(35, 46) <= 0; angryBirdLarge(35, 47) <= 0; angryBirdLarge(35, 48) <= 5; angryBirdLarge(35, 49) <= 5; angryBirdLarge(35, 50) <= 5; angryBirdLarge(35, 51) <= 5; angryBirdLarge(35, 52) <= 5; angryBirdLarge(35, 53) <= 5; angryBirdLarge(35, 54) <= 5; angryBirdLarge(35, 55) <= 5; angryBirdLarge(35, 56) <= 5; angryBirdLarge(35, 57) <= 5; angryBirdLarge(35, 58) <= 5; angryBirdLarge(35, 59) <= 5; angryBirdLarge(35, 60) <= 5; angryBirdLarge(35, 61) <= 5; angryBirdLarge(35, 62) <= 5; angryBirdLarge(35, 63) <= 5; angryBirdLarge(35, 64) <= 5; angryBirdLarge(35, 65) <= 5; angryBirdLarge(35, 66) <= 4; angryBirdLarge(35, 67) <= 4; angryBirdLarge(35, 68) <= 4; angryBirdLarge(35, 69) <= 4; angryBirdLarge(35, 70) <= 4; angryBirdLarge(35, 71) <= 4; angryBirdLarge(35, 72) <= 4; angryBirdLarge(35, 73) <= 4; angryBirdLarge(35, 74) <= 4; angryBirdLarge(35, 75) <= 4; angryBirdLarge(35, 76) <= 4; angryBirdLarge(35, 77) <= 4; angryBirdLarge(35, 78) <= 4; angryBirdLarge(35, 79) <= 4; angryBirdLarge(35, 80) <= 4; angryBirdLarge(35, 81) <= 4; angryBirdLarge(35, 82) <= 4; angryBirdLarge(35, 83) <= 4; angryBirdLarge(35, 84) <= 4; angryBirdLarge(35, 85) <= 4; angryBirdLarge(35, 86) <= 4; angryBirdLarge(35, 87) <= 4; angryBirdLarge(35, 88) <= 4; angryBirdLarge(35, 89) <= 4; angryBirdLarge(35, 90) <= 4; angryBirdLarge(35, 91) <= 4; angryBirdLarge(35, 92) <= 4; angryBirdLarge(35, 93) <= 4; angryBirdLarge(35, 94) <= 4; angryBirdLarge(35, 95) <= 4; angryBirdLarge(35, 96) <= 4; angryBirdLarge(35, 97) <= 4; angryBirdLarge(35, 98) <= 4; angryBirdLarge(35, 99) <= 4; angryBirdLarge(35, 100) <= 4; angryBirdLarge(35, 101) <= 4; angryBirdLarge(35, 102) <= 4; angryBirdLarge(35, 103) <= 4; angryBirdLarge(35, 104) <= 4; angryBirdLarge(35, 105) <= 4; angryBirdLarge(35, 106) <= 4; angryBirdLarge(35, 107) <= 4; angryBirdLarge(35, 108) <= 4; angryBirdLarge(35, 109) <= 4; angryBirdLarge(35, 110) <= 4; angryBirdLarge(35, 111) <= 4; angryBirdLarge(35, 112) <= 4; angryBirdLarge(35, 113) <= 4; angryBirdLarge(35, 114) <= 5; angryBirdLarge(35, 115) <= 5; angryBirdLarge(35, 116) <= 5; angryBirdLarge(35, 117) <= 5; angryBirdLarge(35, 118) <= 5; angryBirdLarge(35, 119) <= 5; angryBirdLarge(35, 120) <= 0; angryBirdLarge(35, 121) <= 0; angryBirdLarge(35, 122) <= 0; angryBirdLarge(35, 123) <= 0; angryBirdLarge(35, 124) <= 0; angryBirdLarge(35, 125) <= 0; angryBirdLarge(35, 126) <= 0; angryBirdLarge(35, 127) <= 0; angryBirdLarge(35, 128) <= 0; angryBirdLarge(35, 129) <= 0; angryBirdLarge(35, 130) <= 0; angryBirdLarge(35, 131) <= 0; angryBirdLarge(35, 132) <= 0; angryBirdLarge(35, 133) <= 0; angryBirdLarge(35, 134) <= 0; angryBirdLarge(35, 135) <= 0; angryBirdLarge(35, 136) <= 0; angryBirdLarge(35, 137) <= 0; angryBirdLarge(35, 138) <= 0; angryBirdLarge(35, 139) <= 0; angryBirdLarge(35, 140) <= 0; angryBirdLarge(35, 141) <= 0; angryBirdLarge(35, 142) <= 0; angryBirdLarge(35, 143) <= 0; angryBirdLarge(35, 144) <= 0; angryBirdLarge(35, 145) <= 0; angryBirdLarge(35, 146) <= 0; angryBirdLarge(35, 147) <= 0; angryBirdLarge(35, 148) <= 0; angryBirdLarge(35, 149) <= 0; 
angryBirdLarge(36, 0) <= 0; angryBirdLarge(36, 1) <= 0; angryBirdLarge(36, 2) <= 0; angryBirdLarge(36, 3) <= 0; angryBirdLarge(36, 4) <= 0; angryBirdLarge(36, 5) <= 0; angryBirdLarge(36, 6) <= 0; angryBirdLarge(36, 7) <= 0; angryBirdLarge(36, 8) <= 0; angryBirdLarge(36, 9) <= 0; angryBirdLarge(36, 10) <= 0; angryBirdLarge(36, 11) <= 0; angryBirdLarge(36, 12) <= 0; angryBirdLarge(36, 13) <= 0; angryBirdLarge(36, 14) <= 0; angryBirdLarge(36, 15) <= 0; angryBirdLarge(36, 16) <= 0; angryBirdLarge(36, 17) <= 0; angryBirdLarge(36, 18) <= 0; angryBirdLarge(36, 19) <= 0; angryBirdLarge(36, 20) <= 0; angryBirdLarge(36, 21) <= 0; angryBirdLarge(36, 22) <= 0; angryBirdLarge(36, 23) <= 0; angryBirdLarge(36, 24) <= 0; angryBirdLarge(36, 25) <= 0; angryBirdLarge(36, 26) <= 0; angryBirdLarge(36, 27) <= 0; angryBirdLarge(36, 28) <= 0; angryBirdLarge(36, 29) <= 0; angryBirdLarge(36, 30) <= 0; angryBirdLarge(36, 31) <= 0; angryBirdLarge(36, 32) <= 0; angryBirdLarge(36, 33) <= 0; angryBirdLarge(36, 34) <= 0; angryBirdLarge(36, 35) <= 0; angryBirdLarge(36, 36) <= 0; angryBirdLarge(36, 37) <= 0; angryBirdLarge(36, 38) <= 0; angryBirdLarge(36, 39) <= 0; angryBirdLarge(36, 40) <= 0; angryBirdLarge(36, 41) <= 0; angryBirdLarge(36, 42) <= 5; angryBirdLarge(36, 43) <= 5; angryBirdLarge(36, 44) <= 5; angryBirdLarge(36, 45) <= 5; angryBirdLarge(36, 46) <= 5; angryBirdLarge(36, 47) <= 5; angryBirdLarge(36, 48) <= 4; angryBirdLarge(36, 49) <= 4; angryBirdLarge(36, 50) <= 4; angryBirdLarge(36, 51) <= 4; angryBirdLarge(36, 52) <= 4; angryBirdLarge(36, 53) <= 4; angryBirdLarge(36, 54) <= 4; angryBirdLarge(36, 55) <= 4; angryBirdLarge(36, 56) <= 4; angryBirdLarge(36, 57) <= 4; angryBirdLarge(36, 58) <= 4; angryBirdLarge(36, 59) <= 4; angryBirdLarge(36, 60) <= 4; angryBirdLarge(36, 61) <= 4; angryBirdLarge(36, 62) <= 4; angryBirdLarge(36, 63) <= 4; angryBirdLarge(36, 64) <= 4; angryBirdLarge(36, 65) <= 4; angryBirdLarge(36, 66) <= 4; angryBirdLarge(36, 67) <= 4; angryBirdLarge(36, 68) <= 4; angryBirdLarge(36, 69) <= 4; angryBirdLarge(36, 70) <= 4; angryBirdLarge(36, 71) <= 4; angryBirdLarge(36, 72) <= 4; angryBirdLarge(36, 73) <= 4; angryBirdLarge(36, 74) <= 4; angryBirdLarge(36, 75) <= 4; angryBirdLarge(36, 76) <= 4; angryBirdLarge(36, 77) <= 4; angryBirdLarge(36, 78) <= 4; angryBirdLarge(36, 79) <= 4; angryBirdLarge(36, 80) <= 4; angryBirdLarge(36, 81) <= 4; angryBirdLarge(36, 82) <= 4; angryBirdLarge(36, 83) <= 4; angryBirdLarge(36, 84) <= 4; angryBirdLarge(36, 85) <= 4; angryBirdLarge(36, 86) <= 4; angryBirdLarge(36, 87) <= 4; angryBirdLarge(36, 88) <= 4; angryBirdLarge(36, 89) <= 4; angryBirdLarge(36, 90) <= 4; angryBirdLarge(36, 91) <= 4; angryBirdLarge(36, 92) <= 4; angryBirdLarge(36, 93) <= 4; angryBirdLarge(36, 94) <= 4; angryBirdLarge(36, 95) <= 4; angryBirdLarge(36, 96) <= 4; angryBirdLarge(36, 97) <= 4; angryBirdLarge(36, 98) <= 4; angryBirdLarge(36, 99) <= 4; angryBirdLarge(36, 100) <= 4; angryBirdLarge(36, 101) <= 4; angryBirdLarge(36, 102) <= 4; angryBirdLarge(36, 103) <= 4; angryBirdLarge(36, 104) <= 4; angryBirdLarge(36, 105) <= 4; angryBirdLarge(36, 106) <= 4; angryBirdLarge(36, 107) <= 4; angryBirdLarge(36, 108) <= 4; angryBirdLarge(36, 109) <= 4; angryBirdLarge(36, 110) <= 4; angryBirdLarge(36, 111) <= 4; angryBirdLarge(36, 112) <= 4; angryBirdLarge(36, 113) <= 4; angryBirdLarge(36, 114) <= 4; angryBirdLarge(36, 115) <= 4; angryBirdLarge(36, 116) <= 4; angryBirdLarge(36, 117) <= 4; angryBirdLarge(36, 118) <= 4; angryBirdLarge(36, 119) <= 4; angryBirdLarge(36, 120) <= 5; angryBirdLarge(36, 121) <= 5; angryBirdLarge(36, 122) <= 5; angryBirdLarge(36, 123) <= 5; angryBirdLarge(36, 124) <= 5; angryBirdLarge(36, 125) <= 5; angryBirdLarge(36, 126) <= 0; angryBirdLarge(36, 127) <= 0; angryBirdLarge(36, 128) <= 0; angryBirdLarge(36, 129) <= 0; angryBirdLarge(36, 130) <= 0; angryBirdLarge(36, 131) <= 0; angryBirdLarge(36, 132) <= 0; angryBirdLarge(36, 133) <= 0; angryBirdLarge(36, 134) <= 0; angryBirdLarge(36, 135) <= 0; angryBirdLarge(36, 136) <= 0; angryBirdLarge(36, 137) <= 0; angryBirdLarge(36, 138) <= 0; angryBirdLarge(36, 139) <= 0; angryBirdLarge(36, 140) <= 0; angryBirdLarge(36, 141) <= 0; angryBirdLarge(36, 142) <= 0; angryBirdLarge(36, 143) <= 0; angryBirdLarge(36, 144) <= 0; angryBirdLarge(36, 145) <= 0; angryBirdLarge(36, 146) <= 0; angryBirdLarge(36, 147) <= 0; angryBirdLarge(36, 148) <= 0; angryBirdLarge(36, 149) <= 0; 
angryBirdLarge(37, 0) <= 0; angryBirdLarge(37, 1) <= 0; angryBirdLarge(37, 2) <= 0; angryBirdLarge(37, 3) <= 0; angryBirdLarge(37, 4) <= 0; angryBirdLarge(37, 5) <= 0; angryBirdLarge(37, 6) <= 0; angryBirdLarge(37, 7) <= 0; angryBirdLarge(37, 8) <= 0; angryBirdLarge(37, 9) <= 0; angryBirdLarge(37, 10) <= 0; angryBirdLarge(37, 11) <= 0; angryBirdLarge(37, 12) <= 0; angryBirdLarge(37, 13) <= 0; angryBirdLarge(37, 14) <= 0; angryBirdLarge(37, 15) <= 0; angryBirdLarge(37, 16) <= 0; angryBirdLarge(37, 17) <= 0; angryBirdLarge(37, 18) <= 0; angryBirdLarge(37, 19) <= 0; angryBirdLarge(37, 20) <= 0; angryBirdLarge(37, 21) <= 0; angryBirdLarge(37, 22) <= 0; angryBirdLarge(37, 23) <= 0; angryBirdLarge(37, 24) <= 0; angryBirdLarge(37, 25) <= 0; angryBirdLarge(37, 26) <= 0; angryBirdLarge(37, 27) <= 0; angryBirdLarge(37, 28) <= 0; angryBirdLarge(37, 29) <= 0; angryBirdLarge(37, 30) <= 0; angryBirdLarge(37, 31) <= 0; angryBirdLarge(37, 32) <= 0; angryBirdLarge(37, 33) <= 0; angryBirdLarge(37, 34) <= 0; angryBirdLarge(37, 35) <= 0; angryBirdLarge(37, 36) <= 0; angryBirdLarge(37, 37) <= 0; angryBirdLarge(37, 38) <= 0; angryBirdLarge(37, 39) <= 0; angryBirdLarge(37, 40) <= 0; angryBirdLarge(37, 41) <= 0; angryBirdLarge(37, 42) <= 5; angryBirdLarge(37, 43) <= 5; angryBirdLarge(37, 44) <= 5; angryBirdLarge(37, 45) <= 5; angryBirdLarge(37, 46) <= 5; angryBirdLarge(37, 47) <= 5; angryBirdLarge(37, 48) <= 4; angryBirdLarge(37, 49) <= 4; angryBirdLarge(37, 50) <= 4; angryBirdLarge(37, 51) <= 4; angryBirdLarge(37, 52) <= 4; angryBirdLarge(37, 53) <= 4; angryBirdLarge(37, 54) <= 4; angryBirdLarge(37, 55) <= 4; angryBirdLarge(37, 56) <= 4; angryBirdLarge(37, 57) <= 4; angryBirdLarge(37, 58) <= 4; angryBirdLarge(37, 59) <= 4; angryBirdLarge(37, 60) <= 4; angryBirdLarge(37, 61) <= 4; angryBirdLarge(37, 62) <= 4; angryBirdLarge(37, 63) <= 4; angryBirdLarge(37, 64) <= 4; angryBirdLarge(37, 65) <= 4; angryBirdLarge(37, 66) <= 4; angryBirdLarge(37, 67) <= 4; angryBirdLarge(37, 68) <= 4; angryBirdLarge(37, 69) <= 4; angryBirdLarge(37, 70) <= 4; angryBirdLarge(37, 71) <= 4; angryBirdLarge(37, 72) <= 4; angryBirdLarge(37, 73) <= 4; angryBirdLarge(37, 74) <= 4; angryBirdLarge(37, 75) <= 4; angryBirdLarge(37, 76) <= 4; angryBirdLarge(37, 77) <= 4; angryBirdLarge(37, 78) <= 4; angryBirdLarge(37, 79) <= 4; angryBirdLarge(37, 80) <= 4; angryBirdLarge(37, 81) <= 4; angryBirdLarge(37, 82) <= 4; angryBirdLarge(37, 83) <= 4; angryBirdLarge(37, 84) <= 4; angryBirdLarge(37, 85) <= 4; angryBirdLarge(37, 86) <= 4; angryBirdLarge(37, 87) <= 4; angryBirdLarge(37, 88) <= 4; angryBirdLarge(37, 89) <= 4; angryBirdLarge(37, 90) <= 4; angryBirdLarge(37, 91) <= 4; angryBirdLarge(37, 92) <= 4; angryBirdLarge(37, 93) <= 4; angryBirdLarge(37, 94) <= 4; angryBirdLarge(37, 95) <= 4; angryBirdLarge(37, 96) <= 4; angryBirdLarge(37, 97) <= 4; angryBirdLarge(37, 98) <= 4; angryBirdLarge(37, 99) <= 4; angryBirdLarge(37, 100) <= 4; angryBirdLarge(37, 101) <= 4; angryBirdLarge(37, 102) <= 4; angryBirdLarge(37, 103) <= 4; angryBirdLarge(37, 104) <= 4; angryBirdLarge(37, 105) <= 4; angryBirdLarge(37, 106) <= 4; angryBirdLarge(37, 107) <= 4; angryBirdLarge(37, 108) <= 4; angryBirdLarge(37, 109) <= 4; angryBirdLarge(37, 110) <= 4; angryBirdLarge(37, 111) <= 4; angryBirdLarge(37, 112) <= 4; angryBirdLarge(37, 113) <= 4; angryBirdLarge(37, 114) <= 4; angryBirdLarge(37, 115) <= 4; angryBirdLarge(37, 116) <= 4; angryBirdLarge(37, 117) <= 4; angryBirdLarge(37, 118) <= 4; angryBirdLarge(37, 119) <= 4; angryBirdLarge(37, 120) <= 5; angryBirdLarge(37, 121) <= 5; angryBirdLarge(37, 122) <= 5; angryBirdLarge(37, 123) <= 5; angryBirdLarge(37, 124) <= 5; angryBirdLarge(37, 125) <= 5; angryBirdLarge(37, 126) <= 0; angryBirdLarge(37, 127) <= 0; angryBirdLarge(37, 128) <= 0; angryBirdLarge(37, 129) <= 0; angryBirdLarge(37, 130) <= 0; angryBirdLarge(37, 131) <= 0; angryBirdLarge(37, 132) <= 0; angryBirdLarge(37, 133) <= 0; angryBirdLarge(37, 134) <= 0; angryBirdLarge(37, 135) <= 0; angryBirdLarge(37, 136) <= 0; angryBirdLarge(37, 137) <= 0; angryBirdLarge(37, 138) <= 0; angryBirdLarge(37, 139) <= 0; angryBirdLarge(37, 140) <= 0; angryBirdLarge(37, 141) <= 0; angryBirdLarge(37, 142) <= 0; angryBirdLarge(37, 143) <= 0; angryBirdLarge(37, 144) <= 0; angryBirdLarge(37, 145) <= 0; angryBirdLarge(37, 146) <= 0; angryBirdLarge(37, 147) <= 0; angryBirdLarge(37, 148) <= 0; angryBirdLarge(37, 149) <= 0; 
angryBirdLarge(38, 0) <= 0; angryBirdLarge(38, 1) <= 0; angryBirdLarge(38, 2) <= 0; angryBirdLarge(38, 3) <= 0; angryBirdLarge(38, 4) <= 0; angryBirdLarge(38, 5) <= 0; angryBirdLarge(38, 6) <= 0; angryBirdLarge(38, 7) <= 0; angryBirdLarge(38, 8) <= 0; angryBirdLarge(38, 9) <= 0; angryBirdLarge(38, 10) <= 0; angryBirdLarge(38, 11) <= 0; angryBirdLarge(38, 12) <= 0; angryBirdLarge(38, 13) <= 0; angryBirdLarge(38, 14) <= 0; angryBirdLarge(38, 15) <= 0; angryBirdLarge(38, 16) <= 0; angryBirdLarge(38, 17) <= 0; angryBirdLarge(38, 18) <= 0; angryBirdLarge(38, 19) <= 0; angryBirdLarge(38, 20) <= 0; angryBirdLarge(38, 21) <= 0; angryBirdLarge(38, 22) <= 0; angryBirdLarge(38, 23) <= 0; angryBirdLarge(38, 24) <= 0; angryBirdLarge(38, 25) <= 0; angryBirdLarge(38, 26) <= 0; angryBirdLarge(38, 27) <= 0; angryBirdLarge(38, 28) <= 0; angryBirdLarge(38, 29) <= 0; angryBirdLarge(38, 30) <= 0; angryBirdLarge(38, 31) <= 0; angryBirdLarge(38, 32) <= 0; angryBirdLarge(38, 33) <= 0; angryBirdLarge(38, 34) <= 0; angryBirdLarge(38, 35) <= 0; angryBirdLarge(38, 36) <= 0; angryBirdLarge(38, 37) <= 0; angryBirdLarge(38, 38) <= 0; angryBirdLarge(38, 39) <= 0; angryBirdLarge(38, 40) <= 0; angryBirdLarge(38, 41) <= 0; angryBirdLarge(38, 42) <= 5; angryBirdLarge(38, 43) <= 5; angryBirdLarge(38, 44) <= 5; angryBirdLarge(38, 45) <= 5; angryBirdLarge(38, 46) <= 5; angryBirdLarge(38, 47) <= 5; angryBirdLarge(38, 48) <= 4; angryBirdLarge(38, 49) <= 4; angryBirdLarge(38, 50) <= 4; angryBirdLarge(38, 51) <= 4; angryBirdLarge(38, 52) <= 4; angryBirdLarge(38, 53) <= 4; angryBirdLarge(38, 54) <= 4; angryBirdLarge(38, 55) <= 4; angryBirdLarge(38, 56) <= 4; angryBirdLarge(38, 57) <= 4; angryBirdLarge(38, 58) <= 4; angryBirdLarge(38, 59) <= 4; angryBirdLarge(38, 60) <= 4; angryBirdLarge(38, 61) <= 4; angryBirdLarge(38, 62) <= 4; angryBirdLarge(38, 63) <= 4; angryBirdLarge(38, 64) <= 4; angryBirdLarge(38, 65) <= 4; angryBirdLarge(38, 66) <= 4; angryBirdLarge(38, 67) <= 4; angryBirdLarge(38, 68) <= 4; angryBirdLarge(38, 69) <= 4; angryBirdLarge(38, 70) <= 4; angryBirdLarge(38, 71) <= 4; angryBirdLarge(38, 72) <= 4; angryBirdLarge(38, 73) <= 4; angryBirdLarge(38, 74) <= 4; angryBirdLarge(38, 75) <= 4; angryBirdLarge(38, 76) <= 4; angryBirdLarge(38, 77) <= 4; angryBirdLarge(38, 78) <= 4; angryBirdLarge(38, 79) <= 4; angryBirdLarge(38, 80) <= 4; angryBirdLarge(38, 81) <= 4; angryBirdLarge(38, 82) <= 4; angryBirdLarge(38, 83) <= 4; angryBirdLarge(38, 84) <= 4; angryBirdLarge(38, 85) <= 4; angryBirdLarge(38, 86) <= 4; angryBirdLarge(38, 87) <= 4; angryBirdLarge(38, 88) <= 4; angryBirdLarge(38, 89) <= 4; angryBirdLarge(38, 90) <= 4; angryBirdLarge(38, 91) <= 4; angryBirdLarge(38, 92) <= 4; angryBirdLarge(38, 93) <= 4; angryBirdLarge(38, 94) <= 4; angryBirdLarge(38, 95) <= 4; angryBirdLarge(38, 96) <= 4; angryBirdLarge(38, 97) <= 4; angryBirdLarge(38, 98) <= 4; angryBirdLarge(38, 99) <= 4; angryBirdLarge(38, 100) <= 4; angryBirdLarge(38, 101) <= 4; angryBirdLarge(38, 102) <= 4; angryBirdLarge(38, 103) <= 4; angryBirdLarge(38, 104) <= 4; angryBirdLarge(38, 105) <= 4; angryBirdLarge(38, 106) <= 4; angryBirdLarge(38, 107) <= 4; angryBirdLarge(38, 108) <= 4; angryBirdLarge(38, 109) <= 4; angryBirdLarge(38, 110) <= 4; angryBirdLarge(38, 111) <= 4; angryBirdLarge(38, 112) <= 4; angryBirdLarge(38, 113) <= 4; angryBirdLarge(38, 114) <= 4; angryBirdLarge(38, 115) <= 4; angryBirdLarge(38, 116) <= 4; angryBirdLarge(38, 117) <= 4; angryBirdLarge(38, 118) <= 4; angryBirdLarge(38, 119) <= 4; angryBirdLarge(38, 120) <= 5; angryBirdLarge(38, 121) <= 5; angryBirdLarge(38, 122) <= 5; angryBirdLarge(38, 123) <= 5; angryBirdLarge(38, 124) <= 5; angryBirdLarge(38, 125) <= 5; angryBirdLarge(38, 126) <= 0; angryBirdLarge(38, 127) <= 0; angryBirdLarge(38, 128) <= 0; angryBirdLarge(38, 129) <= 0; angryBirdLarge(38, 130) <= 0; angryBirdLarge(38, 131) <= 0; angryBirdLarge(38, 132) <= 0; angryBirdLarge(38, 133) <= 0; angryBirdLarge(38, 134) <= 0; angryBirdLarge(38, 135) <= 0; angryBirdLarge(38, 136) <= 0; angryBirdLarge(38, 137) <= 0; angryBirdLarge(38, 138) <= 0; angryBirdLarge(38, 139) <= 0; angryBirdLarge(38, 140) <= 0; angryBirdLarge(38, 141) <= 0; angryBirdLarge(38, 142) <= 0; angryBirdLarge(38, 143) <= 0; angryBirdLarge(38, 144) <= 0; angryBirdLarge(38, 145) <= 0; angryBirdLarge(38, 146) <= 0; angryBirdLarge(38, 147) <= 0; angryBirdLarge(38, 148) <= 0; angryBirdLarge(38, 149) <= 0; 
angryBirdLarge(39, 0) <= 0; angryBirdLarge(39, 1) <= 0; angryBirdLarge(39, 2) <= 0; angryBirdLarge(39, 3) <= 0; angryBirdLarge(39, 4) <= 0; angryBirdLarge(39, 5) <= 0; angryBirdLarge(39, 6) <= 0; angryBirdLarge(39, 7) <= 0; angryBirdLarge(39, 8) <= 0; angryBirdLarge(39, 9) <= 0; angryBirdLarge(39, 10) <= 0; angryBirdLarge(39, 11) <= 0; angryBirdLarge(39, 12) <= 0; angryBirdLarge(39, 13) <= 0; angryBirdLarge(39, 14) <= 0; angryBirdLarge(39, 15) <= 0; angryBirdLarge(39, 16) <= 0; angryBirdLarge(39, 17) <= 0; angryBirdLarge(39, 18) <= 0; angryBirdLarge(39, 19) <= 0; angryBirdLarge(39, 20) <= 0; angryBirdLarge(39, 21) <= 0; angryBirdLarge(39, 22) <= 0; angryBirdLarge(39, 23) <= 0; angryBirdLarge(39, 24) <= 0; angryBirdLarge(39, 25) <= 0; angryBirdLarge(39, 26) <= 0; angryBirdLarge(39, 27) <= 0; angryBirdLarge(39, 28) <= 0; angryBirdLarge(39, 29) <= 0; angryBirdLarge(39, 30) <= 0; angryBirdLarge(39, 31) <= 0; angryBirdLarge(39, 32) <= 0; angryBirdLarge(39, 33) <= 0; angryBirdLarge(39, 34) <= 0; angryBirdLarge(39, 35) <= 0; angryBirdLarge(39, 36) <= 0; angryBirdLarge(39, 37) <= 0; angryBirdLarge(39, 38) <= 0; angryBirdLarge(39, 39) <= 0; angryBirdLarge(39, 40) <= 0; angryBirdLarge(39, 41) <= 0; angryBirdLarge(39, 42) <= 5; angryBirdLarge(39, 43) <= 5; angryBirdLarge(39, 44) <= 5; angryBirdLarge(39, 45) <= 5; angryBirdLarge(39, 46) <= 5; angryBirdLarge(39, 47) <= 5; angryBirdLarge(39, 48) <= 4; angryBirdLarge(39, 49) <= 4; angryBirdLarge(39, 50) <= 4; angryBirdLarge(39, 51) <= 4; angryBirdLarge(39, 52) <= 4; angryBirdLarge(39, 53) <= 4; angryBirdLarge(39, 54) <= 4; angryBirdLarge(39, 55) <= 4; angryBirdLarge(39, 56) <= 4; angryBirdLarge(39, 57) <= 4; angryBirdLarge(39, 58) <= 4; angryBirdLarge(39, 59) <= 4; angryBirdLarge(39, 60) <= 4; angryBirdLarge(39, 61) <= 4; angryBirdLarge(39, 62) <= 4; angryBirdLarge(39, 63) <= 4; angryBirdLarge(39, 64) <= 4; angryBirdLarge(39, 65) <= 4; angryBirdLarge(39, 66) <= 4; angryBirdLarge(39, 67) <= 4; angryBirdLarge(39, 68) <= 4; angryBirdLarge(39, 69) <= 4; angryBirdLarge(39, 70) <= 4; angryBirdLarge(39, 71) <= 4; angryBirdLarge(39, 72) <= 4; angryBirdLarge(39, 73) <= 4; angryBirdLarge(39, 74) <= 4; angryBirdLarge(39, 75) <= 4; angryBirdLarge(39, 76) <= 4; angryBirdLarge(39, 77) <= 4; angryBirdLarge(39, 78) <= 4; angryBirdLarge(39, 79) <= 4; angryBirdLarge(39, 80) <= 4; angryBirdLarge(39, 81) <= 4; angryBirdLarge(39, 82) <= 4; angryBirdLarge(39, 83) <= 4; angryBirdLarge(39, 84) <= 4; angryBirdLarge(39, 85) <= 4; angryBirdLarge(39, 86) <= 4; angryBirdLarge(39, 87) <= 4; angryBirdLarge(39, 88) <= 4; angryBirdLarge(39, 89) <= 4; angryBirdLarge(39, 90) <= 4; angryBirdLarge(39, 91) <= 4; angryBirdLarge(39, 92) <= 4; angryBirdLarge(39, 93) <= 4; angryBirdLarge(39, 94) <= 4; angryBirdLarge(39, 95) <= 4; angryBirdLarge(39, 96) <= 4; angryBirdLarge(39, 97) <= 4; angryBirdLarge(39, 98) <= 4; angryBirdLarge(39, 99) <= 4; angryBirdLarge(39, 100) <= 4; angryBirdLarge(39, 101) <= 4; angryBirdLarge(39, 102) <= 4; angryBirdLarge(39, 103) <= 4; angryBirdLarge(39, 104) <= 4; angryBirdLarge(39, 105) <= 4; angryBirdLarge(39, 106) <= 4; angryBirdLarge(39, 107) <= 4; angryBirdLarge(39, 108) <= 4; angryBirdLarge(39, 109) <= 4; angryBirdLarge(39, 110) <= 4; angryBirdLarge(39, 111) <= 4; angryBirdLarge(39, 112) <= 4; angryBirdLarge(39, 113) <= 4; angryBirdLarge(39, 114) <= 4; angryBirdLarge(39, 115) <= 4; angryBirdLarge(39, 116) <= 4; angryBirdLarge(39, 117) <= 4; angryBirdLarge(39, 118) <= 4; angryBirdLarge(39, 119) <= 4; angryBirdLarge(39, 120) <= 5; angryBirdLarge(39, 121) <= 5; angryBirdLarge(39, 122) <= 5; angryBirdLarge(39, 123) <= 5; angryBirdLarge(39, 124) <= 5; angryBirdLarge(39, 125) <= 5; angryBirdLarge(39, 126) <= 0; angryBirdLarge(39, 127) <= 0; angryBirdLarge(39, 128) <= 0; angryBirdLarge(39, 129) <= 0; angryBirdLarge(39, 130) <= 0; angryBirdLarge(39, 131) <= 0; angryBirdLarge(39, 132) <= 0; angryBirdLarge(39, 133) <= 0; angryBirdLarge(39, 134) <= 0; angryBirdLarge(39, 135) <= 0; angryBirdLarge(39, 136) <= 0; angryBirdLarge(39, 137) <= 0; angryBirdLarge(39, 138) <= 0; angryBirdLarge(39, 139) <= 0; angryBirdLarge(39, 140) <= 0; angryBirdLarge(39, 141) <= 0; angryBirdLarge(39, 142) <= 0; angryBirdLarge(39, 143) <= 0; angryBirdLarge(39, 144) <= 0; angryBirdLarge(39, 145) <= 0; angryBirdLarge(39, 146) <= 0; angryBirdLarge(39, 147) <= 0; angryBirdLarge(39, 148) <= 0; angryBirdLarge(39, 149) <= 0; 
angryBirdLarge(40, 0) <= 0; angryBirdLarge(40, 1) <= 0; angryBirdLarge(40, 2) <= 0; angryBirdLarge(40, 3) <= 0; angryBirdLarge(40, 4) <= 0; angryBirdLarge(40, 5) <= 0; angryBirdLarge(40, 6) <= 0; angryBirdLarge(40, 7) <= 0; angryBirdLarge(40, 8) <= 0; angryBirdLarge(40, 9) <= 0; angryBirdLarge(40, 10) <= 0; angryBirdLarge(40, 11) <= 0; angryBirdLarge(40, 12) <= 0; angryBirdLarge(40, 13) <= 0; angryBirdLarge(40, 14) <= 0; angryBirdLarge(40, 15) <= 0; angryBirdLarge(40, 16) <= 0; angryBirdLarge(40, 17) <= 0; angryBirdLarge(40, 18) <= 0; angryBirdLarge(40, 19) <= 0; angryBirdLarge(40, 20) <= 0; angryBirdLarge(40, 21) <= 0; angryBirdLarge(40, 22) <= 0; angryBirdLarge(40, 23) <= 0; angryBirdLarge(40, 24) <= 0; angryBirdLarge(40, 25) <= 0; angryBirdLarge(40, 26) <= 0; angryBirdLarge(40, 27) <= 0; angryBirdLarge(40, 28) <= 0; angryBirdLarge(40, 29) <= 0; angryBirdLarge(40, 30) <= 0; angryBirdLarge(40, 31) <= 0; angryBirdLarge(40, 32) <= 0; angryBirdLarge(40, 33) <= 0; angryBirdLarge(40, 34) <= 0; angryBirdLarge(40, 35) <= 0; angryBirdLarge(40, 36) <= 0; angryBirdLarge(40, 37) <= 0; angryBirdLarge(40, 38) <= 0; angryBirdLarge(40, 39) <= 0; angryBirdLarge(40, 40) <= 0; angryBirdLarge(40, 41) <= 0; angryBirdLarge(40, 42) <= 5; angryBirdLarge(40, 43) <= 5; angryBirdLarge(40, 44) <= 5; angryBirdLarge(40, 45) <= 5; angryBirdLarge(40, 46) <= 5; angryBirdLarge(40, 47) <= 5; angryBirdLarge(40, 48) <= 4; angryBirdLarge(40, 49) <= 4; angryBirdLarge(40, 50) <= 4; angryBirdLarge(40, 51) <= 4; angryBirdLarge(40, 52) <= 4; angryBirdLarge(40, 53) <= 4; angryBirdLarge(40, 54) <= 4; angryBirdLarge(40, 55) <= 4; angryBirdLarge(40, 56) <= 4; angryBirdLarge(40, 57) <= 4; angryBirdLarge(40, 58) <= 4; angryBirdLarge(40, 59) <= 4; angryBirdLarge(40, 60) <= 4; angryBirdLarge(40, 61) <= 4; angryBirdLarge(40, 62) <= 4; angryBirdLarge(40, 63) <= 4; angryBirdLarge(40, 64) <= 4; angryBirdLarge(40, 65) <= 4; angryBirdLarge(40, 66) <= 4; angryBirdLarge(40, 67) <= 4; angryBirdLarge(40, 68) <= 4; angryBirdLarge(40, 69) <= 4; angryBirdLarge(40, 70) <= 4; angryBirdLarge(40, 71) <= 4; angryBirdLarge(40, 72) <= 4; angryBirdLarge(40, 73) <= 4; angryBirdLarge(40, 74) <= 4; angryBirdLarge(40, 75) <= 4; angryBirdLarge(40, 76) <= 4; angryBirdLarge(40, 77) <= 4; angryBirdLarge(40, 78) <= 4; angryBirdLarge(40, 79) <= 4; angryBirdLarge(40, 80) <= 4; angryBirdLarge(40, 81) <= 4; angryBirdLarge(40, 82) <= 4; angryBirdLarge(40, 83) <= 4; angryBirdLarge(40, 84) <= 4; angryBirdLarge(40, 85) <= 4; angryBirdLarge(40, 86) <= 4; angryBirdLarge(40, 87) <= 4; angryBirdLarge(40, 88) <= 4; angryBirdLarge(40, 89) <= 4; angryBirdLarge(40, 90) <= 4; angryBirdLarge(40, 91) <= 4; angryBirdLarge(40, 92) <= 4; angryBirdLarge(40, 93) <= 4; angryBirdLarge(40, 94) <= 4; angryBirdLarge(40, 95) <= 4; angryBirdLarge(40, 96) <= 4; angryBirdLarge(40, 97) <= 4; angryBirdLarge(40, 98) <= 4; angryBirdLarge(40, 99) <= 4; angryBirdLarge(40, 100) <= 4; angryBirdLarge(40, 101) <= 4; angryBirdLarge(40, 102) <= 4; angryBirdLarge(40, 103) <= 4; angryBirdLarge(40, 104) <= 4; angryBirdLarge(40, 105) <= 4; angryBirdLarge(40, 106) <= 4; angryBirdLarge(40, 107) <= 4; angryBirdLarge(40, 108) <= 4; angryBirdLarge(40, 109) <= 4; angryBirdLarge(40, 110) <= 4; angryBirdLarge(40, 111) <= 4; angryBirdLarge(40, 112) <= 4; angryBirdLarge(40, 113) <= 4; angryBirdLarge(40, 114) <= 4; angryBirdLarge(40, 115) <= 4; angryBirdLarge(40, 116) <= 4; angryBirdLarge(40, 117) <= 4; angryBirdLarge(40, 118) <= 4; angryBirdLarge(40, 119) <= 4; angryBirdLarge(40, 120) <= 5; angryBirdLarge(40, 121) <= 5; angryBirdLarge(40, 122) <= 5; angryBirdLarge(40, 123) <= 5; angryBirdLarge(40, 124) <= 5; angryBirdLarge(40, 125) <= 5; angryBirdLarge(40, 126) <= 0; angryBirdLarge(40, 127) <= 0; angryBirdLarge(40, 128) <= 0; angryBirdLarge(40, 129) <= 0; angryBirdLarge(40, 130) <= 0; angryBirdLarge(40, 131) <= 0; angryBirdLarge(40, 132) <= 0; angryBirdLarge(40, 133) <= 0; angryBirdLarge(40, 134) <= 0; angryBirdLarge(40, 135) <= 0; angryBirdLarge(40, 136) <= 0; angryBirdLarge(40, 137) <= 0; angryBirdLarge(40, 138) <= 0; angryBirdLarge(40, 139) <= 0; angryBirdLarge(40, 140) <= 0; angryBirdLarge(40, 141) <= 0; angryBirdLarge(40, 142) <= 0; angryBirdLarge(40, 143) <= 0; angryBirdLarge(40, 144) <= 0; angryBirdLarge(40, 145) <= 0; angryBirdLarge(40, 146) <= 0; angryBirdLarge(40, 147) <= 0; angryBirdLarge(40, 148) <= 0; angryBirdLarge(40, 149) <= 0; 
angryBirdLarge(41, 0) <= 0; angryBirdLarge(41, 1) <= 0; angryBirdLarge(41, 2) <= 0; angryBirdLarge(41, 3) <= 0; angryBirdLarge(41, 4) <= 0; angryBirdLarge(41, 5) <= 0; angryBirdLarge(41, 6) <= 0; angryBirdLarge(41, 7) <= 0; angryBirdLarge(41, 8) <= 0; angryBirdLarge(41, 9) <= 0; angryBirdLarge(41, 10) <= 0; angryBirdLarge(41, 11) <= 0; angryBirdLarge(41, 12) <= 0; angryBirdLarge(41, 13) <= 0; angryBirdLarge(41, 14) <= 0; angryBirdLarge(41, 15) <= 0; angryBirdLarge(41, 16) <= 0; angryBirdLarge(41, 17) <= 0; angryBirdLarge(41, 18) <= 0; angryBirdLarge(41, 19) <= 0; angryBirdLarge(41, 20) <= 0; angryBirdLarge(41, 21) <= 0; angryBirdLarge(41, 22) <= 0; angryBirdLarge(41, 23) <= 0; angryBirdLarge(41, 24) <= 0; angryBirdLarge(41, 25) <= 0; angryBirdLarge(41, 26) <= 0; angryBirdLarge(41, 27) <= 0; angryBirdLarge(41, 28) <= 0; angryBirdLarge(41, 29) <= 0; angryBirdLarge(41, 30) <= 0; angryBirdLarge(41, 31) <= 0; angryBirdLarge(41, 32) <= 0; angryBirdLarge(41, 33) <= 0; angryBirdLarge(41, 34) <= 0; angryBirdLarge(41, 35) <= 0; angryBirdLarge(41, 36) <= 0; angryBirdLarge(41, 37) <= 0; angryBirdLarge(41, 38) <= 0; angryBirdLarge(41, 39) <= 0; angryBirdLarge(41, 40) <= 0; angryBirdLarge(41, 41) <= 0; angryBirdLarge(41, 42) <= 5; angryBirdLarge(41, 43) <= 5; angryBirdLarge(41, 44) <= 5; angryBirdLarge(41, 45) <= 5; angryBirdLarge(41, 46) <= 5; angryBirdLarge(41, 47) <= 5; angryBirdLarge(41, 48) <= 4; angryBirdLarge(41, 49) <= 4; angryBirdLarge(41, 50) <= 4; angryBirdLarge(41, 51) <= 4; angryBirdLarge(41, 52) <= 4; angryBirdLarge(41, 53) <= 4; angryBirdLarge(41, 54) <= 4; angryBirdLarge(41, 55) <= 4; angryBirdLarge(41, 56) <= 4; angryBirdLarge(41, 57) <= 4; angryBirdLarge(41, 58) <= 4; angryBirdLarge(41, 59) <= 4; angryBirdLarge(41, 60) <= 4; angryBirdLarge(41, 61) <= 4; angryBirdLarge(41, 62) <= 4; angryBirdLarge(41, 63) <= 4; angryBirdLarge(41, 64) <= 4; angryBirdLarge(41, 65) <= 4; angryBirdLarge(41, 66) <= 4; angryBirdLarge(41, 67) <= 4; angryBirdLarge(41, 68) <= 4; angryBirdLarge(41, 69) <= 4; angryBirdLarge(41, 70) <= 4; angryBirdLarge(41, 71) <= 4; angryBirdLarge(41, 72) <= 4; angryBirdLarge(41, 73) <= 4; angryBirdLarge(41, 74) <= 4; angryBirdLarge(41, 75) <= 4; angryBirdLarge(41, 76) <= 4; angryBirdLarge(41, 77) <= 4; angryBirdLarge(41, 78) <= 4; angryBirdLarge(41, 79) <= 4; angryBirdLarge(41, 80) <= 4; angryBirdLarge(41, 81) <= 4; angryBirdLarge(41, 82) <= 4; angryBirdLarge(41, 83) <= 4; angryBirdLarge(41, 84) <= 4; angryBirdLarge(41, 85) <= 4; angryBirdLarge(41, 86) <= 4; angryBirdLarge(41, 87) <= 4; angryBirdLarge(41, 88) <= 4; angryBirdLarge(41, 89) <= 4; angryBirdLarge(41, 90) <= 4; angryBirdLarge(41, 91) <= 4; angryBirdLarge(41, 92) <= 4; angryBirdLarge(41, 93) <= 4; angryBirdLarge(41, 94) <= 4; angryBirdLarge(41, 95) <= 4; angryBirdLarge(41, 96) <= 4; angryBirdLarge(41, 97) <= 4; angryBirdLarge(41, 98) <= 4; angryBirdLarge(41, 99) <= 4; angryBirdLarge(41, 100) <= 4; angryBirdLarge(41, 101) <= 4; angryBirdLarge(41, 102) <= 4; angryBirdLarge(41, 103) <= 4; angryBirdLarge(41, 104) <= 4; angryBirdLarge(41, 105) <= 4; angryBirdLarge(41, 106) <= 4; angryBirdLarge(41, 107) <= 4; angryBirdLarge(41, 108) <= 4; angryBirdLarge(41, 109) <= 4; angryBirdLarge(41, 110) <= 4; angryBirdLarge(41, 111) <= 4; angryBirdLarge(41, 112) <= 4; angryBirdLarge(41, 113) <= 4; angryBirdLarge(41, 114) <= 4; angryBirdLarge(41, 115) <= 4; angryBirdLarge(41, 116) <= 4; angryBirdLarge(41, 117) <= 4; angryBirdLarge(41, 118) <= 4; angryBirdLarge(41, 119) <= 4; angryBirdLarge(41, 120) <= 5; angryBirdLarge(41, 121) <= 5; angryBirdLarge(41, 122) <= 5; angryBirdLarge(41, 123) <= 5; angryBirdLarge(41, 124) <= 5; angryBirdLarge(41, 125) <= 5; angryBirdLarge(41, 126) <= 0; angryBirdLarge(41, 127) <= 0; angryBirdLarge(41, 128) <= 0; angryBirdLarge(41, 129) <= 0; angryBirdLarge(41, 130) <= 0; angryBirdLarge(41, 131) <= 0; angryBirdLarge(41, 132) <= 0; angryBirdLarge(41, 133) <= 0; angryBirdLarge(41, 134) <= 0; angryBirdLarge(41, 135) <= 0; angryBirdLarge(41, 136) <= 0; angryBirdLarge(41, 137) <= 0; angryBirdLarge(41, 138) <= 0; angryBirdLarge(41, 139) <= 0; angryBirdLarge(41, 140) <= 0; angryBirdLarge(41, 141) <= 0; angryBirdLarge(41, 142) <= 0; angryBirdLarge(41, 143) <= 0; angryBirdLarge(41, 144) <= 0; angryBirdLarge(41, 145) <= 0; angryBirdLarge(41, 146) <= 0; angryBirdLarge(41, 147) <= 0; angryBirdLarge(41, 148) <= 0; angryBirdLarge(41, 149) <= 0; 
angryBirdLarge(42, 0) <= 0; angryBirdLarge(42, 1) <= 0; angryBirdLarge(42, 2) <= 0; angryBirdLarge(42, 3) <= 0; angryBirdLarge(42, 4) <= 0; angryBirdLarge(42, 5) <= 0; angryBirdLarge(42, 6) <= 0; angryBirdLarge(42, 7) <= 0; angryBirdLarge(42, 8) <= 0; angryBirdLarge(42, 9) <= 0; angryBirdLarge(42, 10) <= 0; angryBirdLarge(42, 11) <= 0; angryBirdLarge(42, 12) <= 0; angryBirdLarge(42, 13) <= 0; angryBirdLarge(42, 14) <= 0; angryBirdLarge(42, 15) <= 0; angryBirdLarge(42, 16) <= 0; angryBirdLarge(42, 17) <= 0; angryBirdLarge(42, 18) <= 0; angryBirdLarge(42, 19) <= 0; angryBirdLarge(42, 20) <= 0; angryBirdLarge(42, 21) <= 0; angryBirdLarge(42, 22) <= 0; angryBirdLarge(42, 23) <= 0; angryBirdLarge(42, 24) <= 0; angryBirdLarge(42, 25) <= 0; angryBirdLarge(42, 26) <= 0; angryBirdLarge(42, 27) <= 0; angryBirdLarge(42, 28) <= 0; angryBirdLarge(42, 29) <= 0; angryBirdLarge(42, 30) <= 0; angryBirdLarge(42, 31) <= 0; angryBirdLarge(42, 32) <= 0; angryBirdLarge(42, 33) <= 0; angryBirdLarge(42, 34) <= 0; angryBirdLarge(42, 35) <= 0; angryBirdLarge(42, 36) <= 5; angryBirdLarge(42, 37) <= 5; angryBirdLarge(42, 38) <= 5; angryBirdLarge(42, 39) <= 5; angryBirdLarge(42, 40) <= 5; angryBirdLarge(42, 41) <= 5; angryBirdLarge(42, 42) <= 4; angryBirdLarge(42, 43) <= 4; angryBirdLarge(42, 44) <= 4; angryBirdLarge(42, 45) <= 4; angryBirdLarge(42, 46) <= 4; angryBirdLarge(42, 47) <= 4; angryBirdLarge(42, 48) <= 4; angryBirdLarge(42, 49) <= 4; angryBirdLarge(42, 50) <= 4; angryBirdLarge(42, 51) <= 4; angryBirdLarge(42, 52) <= 4; angryBirdLarge(42, 53) <= 4; angryBirdLarge(42, 54) <= 4; angryBirdLarge(42, 55) <= 4; angryBirdLarge(42, 56) <= 4; angryBirdLarge(42, 57) <= 4; angryBirdLarge(42, 58) <= 4; angryBirdLarge(42, 59) <= 4; angryBirdLarge(42, 60) <= 4; angryBirdLarge(42, 61) <= 4; angryBirdLarge(42, 62) <= 4; angryBirdLarge(42, 63) <= 4; angryBirdLarge(42, 64) <= 4; angryBirdLarge(42, 65) <= 4; angryBirdLarge(42, 66) <= 4; angryBirdLarge(42, 67) <= 4; angryBirdLarge(42, 68) <= 4; angryBirdLarge(42, 69) <= 4; angryBirdLarge(42, 70) <= 4; angryBirdLarge(42, 71) <= 4; angryBirdLarge(42, 72) <= 4; angryBirdLarge(42, 73) <= 4; angryBirdLarge(42, 74) <= 4; angryBirdLarge(42, 75) <= 4; angryBirdLarge(42, 76) <= 4; angryBirdLarge(42, 77) <= 4; angryBirdLarge(42, 78) <= 4; angryBirdLarge(42, 79) <= 4; angryBirdLarge(42, 80) <= 4; angryBirdLarge(42, 81) <= 4; angryBirdLarge(42, 82) <= 4; angryBirdLarge(42, 83) <= 4; angryBirdLarge(42, 84) <= 4; angryBirdLarge(42, 85) <= 4; angryBirdLarge(42, 86) <= 4; angryBirdLarge(42, 87) <= 4; angryBirdLarge(42, 88) <= 4; angryBirdLarge(42, 89) <= 4; angryBirdLarge(42, 90) <= 4; angryBirdLarge(42, 91) <= 4; angryBirdLarge(42, 92) <= 4; angryBirdLarge(42, 93) <= 4; angryBirdLarge(42, 94) <= 4; angryBirdLarge(42, 95) <= 4; angryBirdLarge(42, 96) <= 4; angryBirdLarge(42, 97) <= 4; angryBirdLarge(42, 98) <= 4; angryBirdLarge(42, 99) <= 4; angryBirdLarge(42, 100) <= 4; angryBirdLarge(42, 101) <= 4; angryBirdLarge(42, 102) <= 4; angryBirdLarge(42, 103) <= 4; angryBirdLarge(42, 104) <= 4; angryBirdLarge(42, 105) <= 4; angryBirdLarge(42, 106) <= 4; angryBirdLarge(42, 107) <= 4; angryBirdLarge(42, 108) <= 4; angryBirdLarge(42, 109) <= 4; angryBirdLarge(42, 110) <= 4; angryBirdLarge(42, 111) <= 4; angryBirdLarge(42, 112) <= 4; angryBirdLarge(42, 113) <= 4; angryBirdLarge(42, 114) <= 4; angryBirdLarge(42, 115) <= 4; angryBirdLarge(42, 116) <= 4; angryBirdLarge(42, 117) <= 4; angryBirdLarge(42, 118) <= 4; angryBirdLarge(42, 119) <= 4; angryBirdLarge(42, 120) <= 4; angryBirdLarge(42, 121) <= 4; angryBirdLarge(42, 122) <= 4; angryBirdLarge(42, 123) <= 4; angryBirdLarge(42, 124) <= 4; angryBirdLarge(42, 125) <= 4; angryBirdLarge(42, 126) <= 5; angryBirdLarge(42, 127) <= 5; angryBirdLarge(42, 128) <= 5; angryBirdLarge(42, 129) <= 5; angryBirdLarge(42, 130) <= 5; angryBirdLarge(42, 131) <= 5; angryBirdLarge(42, 132) <= 0; angryBirdLarge(42, 133) <= 0; angryBirdLarge(42, 134) <= 0; angryBirdLarge(42, 135) <= 0; angryBirdLarge(42, 136) <= 0; angryBirdLarge(42, 137) <= 0; angryBirdLarge(42, 138) <= 0; angryBirdLarge(42, 139) <= 0; angryBirdLarge(42, 140) <= 0; angryBirdLarge(42, 141) <= 0; angryBirdLarge(42, 142) <= 0; angryBirdLarge(42, 143) <= 0; angryBirdLarge(42, 144) <= 0; angryBirdLarge(42, 145) <= 0; angryBirdLarge(42, 146) <= 0; angryBirdLarge(42, 147) <= 0; angryBirdLarge(42, 148) <= 0; angryBirdLarge(42, 149) <= 0; 
angryBirdLarge(43, 0) <= 0; angryBirdLarge(43, 1) <= 0; angryBirdLarge(43, 2) <= 0; angryBirdLarge(43, 3) <= 0; angryBirdLarge(43, 4) <= 0; angryBirdLarge(43, 5) <= 0; angryBirdLarge(43, 6) <= 0; angryBirdLarge(43, 7) <= 0; angryBirdLarge(43, 8) <= 0; angryBirdLarge(43, 9) <= 0; angryBirdLarge(43, 10) <= 0; angryBirdLarge(43, 11) <= 0; angryBirdLarge(43, 12) <= 0; angryBirdLarge(43, 13) <= 0; angryBirdLarge(43, 14) <= 0; angryBirdLarge(43, 15) <= 0; angryBirdLarge(43, 16) <= 0; angryBirdLarge(43, 17) <= 0; angryBirdLarge(43, 18) <= 0; angryBirdLarge(43, 19) <= 0; angryBirdLarge(43, 20) <= 0; angryBirdLarge(43, 21) <= 0; angryBirdLarge(43, 22) <= 0; angryBirdLarge(43, 23) <= 0; angryBirdLarge(43, 24) <= 0; angryBirdLarge(43, 25) <= 0; angryBirdLarge(43, 26) <= 0; angryBirdLarge(43, 27) <= 0; angryBirdLarge(43, 28) <= 0; angryBirdLarge(43, 29) <= 0; angryBirdLarge(43, 30) <= 0; angryBirdLarge(43, 31) <= 0; angryBirdLarge(43, 32) <= 0; angryBirdLarge(43, 33) <= 0; angryBirdLarge(43, 34) <= 0; angryBirdLarge(43, 35) <= 0; angryBirdLarge(43, 36) <= 5; angryBirdLarge(43, 37) <= 5; angryBirdLarge(43, 38) <= 5; angryBirdLarge(43, 39) <= 5; angryBirdLarge(43, 40) <= 5; angryBirdLarge(43, 41) <= 5; angryBirdLarge(43, 42) <= 4; angryBirdLarge(43, 43) <= 4; angryBirdLarge(43, 44) <= 4; angryBirdLarge(43, 45) <= 4; angryBirdLarge(43, 46) <= 4; angryBirdLarge(43, 47) <= 4; angryBirdLarge(43, 48) <= 4; angryBirdLarge(43, 49) <= 4; angryBirdLarge(43, 50) <= 4; angryBirdLarge(43, 51) <= 4; angryBirdLarge(43, 52) <= 4; angryBirdLarge(43, 53) <= 4; angryBirdLarge(43, 54) <= 4; angryBirdLarge(43, 55) <= 4; angryBirdLarge(43, 56) <= 4; angryBirdLarge(43, 57) <= 4; angryBirdLarge(43, 58) <= 4; angryBirdLarge(43, 59) <= 4; angryBirdLarge(43, 60) <= 4; angryBirdLarge(43, 61) <= 4; angryBirdLarge(43, 62) <= 4; angryBirdLarge(43, 63) <= 4; angryBirdLarge(43, 64) <= 4; angryBirdLarge(43, 65) <= 4; angryBirdLarge(43, 66) <= 4; angryBirdLarge(43, 67) <= 4; angryBirdLarge(43, 68) <= 4; angryBirdLarge(43, 69) <= 4; angryBirdLarge(43, 70) <= 4; angryBirdLarge(43, 71) <= 4; angryBirdLarge(43, 72) <= 4; angryBirdLarge(43, 73) <= 4; angryBirdLarge(43, 74) <= 4; angryBirdLarge(43, 75) <= 4; angryBirdLarge(43, 76) <= 4; angryBirdLarge(43, 77) <= 4; angryBirdLarge(43, 78) <= 4; angryBirdLarge(43, 79) <= 4; angryBirdLarge(43, 80) <= 4; angryBirdLarge(43, 81) <= 4; angryBirdLarge(43, 82) <= 4; angryBirdLarge(43, 83) <= 4; angryBirdLarge(43, 84) <= 4; angryBirdLarge(43, 85) <= 4; angryBirdLarge(43, 86) <= 4; angryBirdLarge(43, 87) <= 4; angryBirdLarge(43, 88) <= 4; angryBirdLarge(43, 89) <= 4; angryBirdLarge(43, 90) <= 4; angryBirdLarge(43, 91) <= 4; angryBirdLarge(43, 92) <= 4; angryBirdLarge(43, 93) <= 4; angryBirdLarge(43, 94) <= 4; angryBirdLarge(43, 95) <= 4; angryBirdLarge(43, 96) <= 4; angryBirdLarge(43, 97) <= 4; angryBirdLarge(43, 98) <= 4; angryBirdLarge(43, 99) <= 4; angryBirdLarge(43, 100) <= 4; angryBirdLarge(43, 101) <= 4; angryBirdLarge(43, 102) <= 4; angryBirdLarge(43, 103) <= 4; angryBirdLarge(43, 104) <= 4; angryBirdLarge(43, 105) <= 4; angryBirdLarge(43, 106) <= 4; angryBirdLarge(43, 107) <= 4; angryBirdLarge(43, 108) <= 4; angryBirdLarge(43, 109) <= 4; angryBirdLarge(43, 110) <= 4; angryBirdLarge(43, 111) <= 4; angryBirdLarge(43, 112) <= 4; angryBirdLarge(43, 113) <= 4; angryBirdLarge(43, 114) <= 4; angryBirdLarge(43, 115) <= 4; angryBirdLarge(43, 116) <= 4; angryBirdLarge(43, 117) <= 4; angryBirdLarge(43, 118) <= 4; angryBirdLarge(43, 119) <= 4; angryBirdLarge(43, 120) <= 4; angryBirdLarge(43, 121) <= 4; angryBirdLarge(43, 122) <= 4; angryBirdLarge(43, 123) <= 4; angryBirdLarge(43, 124) <= 4; angryBirdLarge(43, 125) <= 4; angryBirdLarge(43, 126) <= 5; angryBirdLarge(43, 127) <= 5; angryBirdLarge(43, 128) <= 5; angryBirdLarge(43, 129) <= 5; angryBirdLarge(43, 130) <= 5; angryBirdLarge(43, 131) <= 5; angryBirdLarge(43, 132) <= 0; angryBirdLarge(43, 133) <= 0; angryBirdLarge(43, 134) <= 0; angryBirdLarge(43, 135) <= 0; angryBirdLarge(43, 136) <= 0; angryBirdLarge(43, 137) <= 0; angryBirdLarge(43, 138) <= 0; angryBirdLarge(43, 139) <= 0; angryBirdLarge(43, 140) <= 0; angryBirdLarge(43, 141) <= 0; angryBirdLarge(43, 142) <= 0; angryBirdLarge(43, 143) <= 0; angryBirdLarge(43, 144) <= 0; angryBirdLarge(43, 145) <= 0; angryBirdLarge(43, 146) <= 0; angryBirdLarge(43, 147) <= 0; angryBirdLarge(43, 148) <= 0; angryBirdLarge(43, 149) <= 0; 
angryBirdLarge(44, 0) <= 0; angryBirdLarge(44, 1) <= 0; angryBirdLarge(44, 2) <= 0; angryBirdLarge(44, 3) <= 0; angryBirdLarge(44, 4) <= 0; angryBirdLarge(44, 5) <= 0; angryBirdLarge(44, 6) <= 0; angryBirdLarge(44, 7) <= 0; angryBirdLarge(44, 8) <= 0; angryBirdLarge(44, 9) <= 0; angryBirdLarge(44, 10) <= 0; angryBirdLarge(44, 11) <= 0; angryBirdLarge(44, 12) <= 0; angryBirdLarge(44, 13) <= 0; angryBirdLarge(44, 14) <= 0; angryBirdLarge(44, 15) <= 0; angryBirdLarge(44, 16) <= 0; angryBirdLarge(44, 17) <= 0; angryBirdLarge(44, 18) <= 0; angryBirdLarge(44, 19) <= 0; angryBirdLarge(44, 20) <= 0; angryBirdLarge(44, 21) <= 0; angryBirdLarge(44, 22) <= 0; angryBirdLarge(44, 23) <= 0; angryBirdLarge(44, 24) <= 0; angryBirdLarge(44, 25) <= 0; angryBirdLarge(44, 26) <= 0; angryBirdLarge(44, 27) <= 0; angryBirdLarge(44, 28) <= 0; angryBirdLarge(44, 29) <= 0; angryBirdLarge(44, 30) <= 0; angryBirdLarge(44, 31) <= 0; angryBirdLarge(44, 32) <= 0; angryBirdLarge(44, 33) <= 0; angryBirdLarge(44, 34) <= 0; angryBirdLarge(44, 35) <= 0; angryBirdLarge(44, 36) <= 5; angryBirdLarge(44, 37) <= 5; angryBirdLarge(44, 38) <= 5; angryBirdLarge(44, 39) <= 5; angryBirdLarge(44, 40) <= 5; angryBirdLarge(44, 41) <= 5; angryBirdLarge(44, 42) <= 4; angryBirdLarge(44, 43) <= 4; angryBirdLarge(44, 44) <= 4; angryBirdLarge(44, 45) <= 4; angryBirdLarge(44, 46) <= 4; angryBirdLarge(44, 47) <= 4; angryBirdLarge(44, 48) <= 4; angryBirdLarge(44, 49) <= 4; angryBirdLarge(44, 50) <= 4; angryBirdLarge(44, 51) <= 4; angryBirdLarge(44, 52) <= 4; angryBirdLarge(44, 53) <= 4; angryBirdLarge(44, 54) <= 4; angryBirdLarge(44, 55) <= 4; angryBirdLarge(44, 56) <= 4; angryBirdLarge(44, 57) <= 4; angryBirdLarge(44, 58) <= 4; angryBirdLarge(44, 59) <= 4; angryBirdLarge(44, 60) <= 4; angryBirdLarge(44, 61) <= 4; angryBirdLarge(44, 62) <= 4; angryBirdLarge(44, 63) <= 4; angryBirdLarge(44, 64) <= 4; angryBirdLarge(44, 65) <= 4; angryBirdLarge(44, 66) <= 4; angryBirdLarge(44, 67) <= 4; angryBirdLarge(44, 68) <= 4; angryBirdLarge(44, 69) <= 4; angryBirdLarge(44, 70) <= 4; angryBirdLarge(44, 71) <= 4; angryBirdLarge(44, 72) <= 4; angryBirdLarge(44, 73) <= 4; angryBirdLarge(44, 74) <= 4; angryBirdLarge(44, 75) <= 4; angryBirdLarge(44, 76) <= 4; angryBirdLarge(44, 77) <= 4; angryBirdLarge(44, 78) <= 4; angryBirdLarge(44, 79) <= 4; angryBirdLarge(44, 80) <= 4; angryBirdLarge(44, 81) <= 4; angryBirdLarge(44, 82) <= 4; angryBirdLarge(44, 83) <= 4; angryBirdLarge(44, 84) <= 4; angryBirdLarge(44, 85) <= 4; angryBirdLarge(44, 86) <= 4; angryBirdLarge(44, 87) <= 4; angryBirdLarge(44, 88) <= 4; angryBirdLarge(44, 89) <= 4; angryBirdLarge(44, 90) <= 4; angryBirdLarge(44, 91) <= 4; angryBirdLarge(44, 92) <= 4; angryBirdLarge(44, 93) <= 4; angryBirdLarge(44, 94) <= 4; angryBirdLarge(44, 95) <= 4; angryBirdLarge(44, 96) <= 4; angryBirdLarge(44, 97) <= 4; angryBirdLarge(44, 98) <= 4; angryBirdLarge(44, 99) <= 4; angryBirdLarge(44, 100) <= 4; angryBirdLarge(44, 101) <= 4; angryBirdLarge(44, 102) <= 4; angryBirdLarge(44, 103) <= 4; angryBirdLarge(44, 104) <= 4; angryBirdLarge(44, 105) <= 4; angryBirdLarge(44, 106) <= 4; angryBirdLarge(44, 107) <= 4; angryBirdLarge(44, 108) <= 4; angryBirdLarge(44, 109) <= 4; angryBirdLarge(44, 110) <= 4; angryBirdLarge(44, 111) <= 4; angryBirdLarge(44, 112) <= 4; angryBirdLarge(44, 113) <= 4; angryBirdLarge(44, 114) <= 4; angryBirdLarge(44, 115) <= 4; angryBirdLarge(44, 116) <= 4; angryBirdLarge(44, 117) <= 4; angryBirdLarge(44, 118) <= 4; angryBirdLarge(44, 119) <= 4; angryBirdLarge(44, 120) <= 4; angryBirdLarge(44, 121) <= 4; angryBirdLarge(44, 122) <= 4; angryBirdLarge(44, 123) <= 4; angryBirdLarge(44, 124) <= 4; angryBirdLarge(44, 125) <= 4; angryBirdLarge(44, 126) <= 5; angryBirdLarge(44, 127) <= 5; angryBirdLarge(44, 128) <= 5; angryBirdLarge(44, 129) <= 5; angryBirdLarge(44, 130) <= 5; angryBirdLarge(44, 131) <= 5; angryBirdLarge(44, 132) <= 0; angryBirdLarge(44, 133) <= 0; angryBirdLarge(44, 134) <= 0; angryBirdLarge(44, 135) <= 0; angryBirdLarge(44, 136) <= 0; angryBirdLarge(44, 137) <= 0; angryBirdLarge(44, 138) <= 0; angryBirdLarge(44, 139) <= 0; angryBirdLarge(44, 140) <= 0; angryBirdLarge(44, 141) <= 0; angryBirdLarge(44, 142) <= 0; angryBirdLarge(44, 143) <= 0; angryBirdLarge(44, 144) <= 0; angryBirdLarge(44, 145) <= 0; angryBirdLarge(44, 146) <= 0; angryBirdLarge(44, 147) <= 0; angryBirdLarge(44, 148) <= 0; angryBirdLarge(44, 149) <= 0; 
angryBirdLarge(45, 0) <= 0; angryBirdLarge(45, 1) <= 0; angryBirdLarge(45, 2) <= 0; angryBirdLarge(45, 3) <= 0; angryBirdLarge(45, 4) <= 0; angryBirdLarge(45, 5) <= 0; angryBirdLarge(45, 6) <= 0; angryBirdLarge(45, 7) <= 0; angryBirdLarge(45, 8) <= 0; angryBirdLarge(45, 9) <= 0; angryBirdLarge(45, 10) <= 0; angryBirdLarge(45, 11) <= 0; angryBirdLarge(45, 12) <= 0; angryBirdLarge(45, 13) <= 0; angryBirdLarge(45, 14) <= 0; angryBirdLarge(45, 15) <= 0; angryBirdLarge(45, 16) <= 0; angryBirdLarge(45, 17) <= 0; angryBirdLarge(45, 18) <= 0; angryBirdLarge(45, 19) <= 0; angryBirdLarge(45, 20) <= 0; angryBirdLarge(45, 21) <= 0; angryBirdLarge(45, 22) <= 0; angryBirdLarge(45, 23) <= 0; angryBirdLarge(45, 24) <= 0; angryBirdLarge(45, 25) <= 0; angryBirdLarge(45, 26) <= 0; angryBirdLarge(45, 27) <= 0; angryBirdLarge(45, 28) <= 0; angryBirdLarge(45, 29) <= 0; angryBirdLarge(45, 30) <= 0; angryBirdLarge(45, 31) <= 0; angryBirdLarge(45, 32) <= 0; angryBirdLarge(45, 33) <= 0; angryBirdLarge(45, 34) <= 0; angryBirdLarge(45, 35) <= 0; angryBirdLarge(45, 36) <= 5; angryBirdLarge(45, 37) <= 5; angryBirdLarge(45, 38) <= 5; angryBirdLarge(45, 39) <= 5; angryBirdLarge(45, 40) <= 5; angryBirdLarge(45, 41) <= 5; angryBirdLarge(45, 42) <= 4; angryBirdLarge(45, 43) <= 4; angryBirdLarge(45, 44) <= 4; angryBirdLarge(45, 45) <= 4; angryBirdLarge(45, 46) <= 4; angryBirdLarge(45, 47) <= 4; angryBirdLarge(45, 48) <= 4; angryBirdLarge(45, 49) <= 4; angryBirdLarge(45, 50) <= 4; angryBirdLarge(45, 51) <= 4; angryBirdLarge(45, 52) <= 4; angryBirdLarge(45, 53) <= 4; angryBirdLarge(45, 54) <= 4; angryBirdLarge(45, 55) <= 4; angryBirdLarge(45, 56) <= 4; angryBirdLarge(45, 57) <= 4; angryBirdLarge(45, 58) <= 4; angryBirdLarge(45, 59) <= 4; angryBirdLarge(45, 60) <= 4; angryBirdLarge(45, 61) <= 4; angryBirdLarge(45, 62) <= 4; angryBirdLarge(45, 63) <= 4; angryBirdLarge(45, 64) <= 4; angryBirdLarge(45, 65) <= 4; angryBirdLarge(45, 66) <= 4; angryBirdLarge(45, 67) <= 4; angryBirdLarge(45, 68) <= 4; angryBirdLarge(45, 69) <= 4; angryBirdLarge(45, 70) <= 4; angryBirdLarge(45, 71) <= 4; angryBirdLarge(45, 72) <= 4; angryBirdLarge(45, 73) <= 4; angryBirdLarge(45, 74) <= 4; angryBirdLarge(45, 75) <= 4; angryBirdLarge(45, 76) <= 4; angryBirdLarge(45, 77) <= 4; angryBirdLarge(45, 78) <= 4; angryBirdLarge(45, 79) <= 4; angryBirdLarge(45, 80) <= 4; angryBirdLarge(45, 81) <= 4; angryBirdLarge(45, 82) <= 4; angryBirdLarge(45, 83) <= 4; angryBirdLarge(45, 84) <= 4; angryBirdLarge(45, 85) <= 4; angryBirdLarge(45, 86) <= 4; angryBirdLarge(45, 87) <= 4; angryBirdLarge(45, 88) <= 4; angryBirdLarge(45, 89) <= 4; angryBirdLarge(45, 90) <= 4; angryBirdLarge(45, 91) <= 4; angryBirdLarge(45, 92) <= 4; angryBirdLarge(45, 93) <= 4; angryBirdLarge(45, 94) <= 4; angryBirdLarge(45, 95) <= 4; angryBirdLarge(45, 96) <= 4; angryBirdLarge(45, 97) <= 4; angryBirdLarge(45, 98) <= 4; angryBirdLarge(45, 99) <= 4; angryBirdLarge(45, 100) <= 4; angryBirdLarge(45, 101) <= 4; angryBirdLarge(45, 102) <= 4; angryBirdLarge(45, 103) <= 4; angryBirdLarge(45, 104) <= 4; angryBirdLarge(45, 105) <= 4; angryBirdLarge(45, 106) <= 4; angryBirdLarge(45, 107) <= 4; angryBirdLarge(45, 108) <= 4; angryBirdLarge(45, 109) <= 4; angryBirdLarge(45, 110) <= 4; angryBirdLarge(45, 111) <= 4; angryBirdLarge(45, 112) <= 4; angryBirdLarge(45, 113) <= 4; angryBirdLarge(45, 114) <= 4; angryBirdLarge(45, 115) <= 4; angryBirdLarge(45, 116) <= 4; angryBirdLarge(45, 117) <= 4; angryBirdLarge(45, 118) <= 4; angryBirdLarge(45, 119) <= 4; angryBirdLarge(45, 120) <= 4; angryBirdLarge(45, 121) <= 4; angryBirdLarge(45, 122) <= 4; angryBirdLarge(45, 123) <= 4; angryBirdLarge(45, 124) <= 4; angryBirdLarge(45, 125) <= 4; angryBirdLarge(45, 126) <= 5; angryBirdLarge(45, 127) <= 5; angryBirdLarge(45, 128) <= 5; angryBirdLarge(45, 129) <= 5; angryBirdLarge(45, 130) <= 5; angryBirdLarge(45, 131) <= 5; angryBirdLarge(45, 132) <= 0; angryBirdLarge(45, 133) <= 0; angryBirdLarge(45, 134) <= 0; angryBirdLarge(45, 135) <= 0; angryBirdLarge(45, 136) <= 0; angryBirdLarge(45, 137) <= 0; angryBirdLarge(45, 138) <= 0; angryBirdLarge(45, 139) <= 0; angryBirdLarge(45, 140) <= 0; angryBirdLarge(45, 141) <= 0; angryBirdLarge(45, 142) <= 0; angryBirdLarge(45, 143) <= 0; angryBirdLarge(45, 144) <= 0; angryBirdLarge(45, 145) <= 0; angryBirdLarge(45, 146) <= 0; angryBirdLarge(45, 147) <= 0; angryBirdLarge(45, 148) <= 0; angryBirdLarge(45, 149) <= 0; 
angryBirdLarge(46, 0) <= 0; angryBirdLarge(46, 1) <= 0; angryBirdLarge(46, 2) <= 0; angryBirdLarge(46, 3) <= 0; angryBirdLarge(46, 4) <= 0; angryBirdLarge(46, 5) <= 0; angryBirdLarge(46, 6) <= 0; angryBirdLarge(46, 7) <= 0; angryBirdLarge(46, 8) <= 0; angryBirdLarge(46, 9) <= 0; angryBirdLarge(46, 10) <= 0; angryBirdLarge(46, 11) <= 0; angryBirdLarge(46, 12) <= 0; angryBirdLarge(46, 13) <= 0; angryBirdLarge(46, 14) <= 0; angryBirdLarge(46, 15) <= 0; angryBirdLarge(46, 16) <= 0; angryBirdLarge(46, 17) <= 0; angryBirdLarge(46, 18) <= 0; angryBirdLarge(46, 19) <= 0; angryBirdLarge(46, 20) <= 0; angryBirdLarge(46, 21) <= 0; angryBirdLarge(46, 22) <= 0; angryBirdLarge(46, 23) <= 0; angryBirdLarge(46, 24) <= 0; angryBirdLarge(46, 25) <= 0; angryBirdLarge(46, 26) <= 0; angryBirdLarge(46, 27) <= 0; angryBirdLarge(46, 28) <= 0; angryBirdLarge(46, 29) <= 0; angryBirdLarge(46, 30) <= 0; angryBirdLarge(46, 31) <= 0; angryBirdLarge(46, 32) <= 0; angryBirdLarge(46, 33) <= 0; angryBirdLarge(46, 34) <= 0; angryBirdLarge(46, 35) <= 0; angryBirdLarge(46, 36) <= 5; angryBirdLarge(46, 37) <= 5; angryBirdLarge(46, 38) <= 5; angryBirdLarge(46, 39) <= 5; angryBirdLarge(46, 40) <= 5; angryBirdLarge(46, 41) <= 5; angryBirdLarge(46, 42) <= 4; angryBirdLarge(46, 43) <= 4; angryBirdLarge(46, 44) <= 4; angryBirdLarge(46, 45) <= 4; angryBirdLarge(46, 46) <= 4; angryBirdLarge(46, 47) <= 4; angryBirdLarge(46, 48) <= 4; angryBirdLarge(46, 49) <= 4; angryBirdLarge(46, 50) <= 4; angryBirdLarge(46, 51) <= 4; angryBirdLarge(46, 52) <= 4; angryBirdLarge(46, 53) <= 4; angryBirdLarge(46, 54) <= 4; angryBirdLarge(46, 55) <= 4; angryBirdLarge(46, 56) <= 4; angryBirdLarge(46, 57) <= 4; angryBirdLarge(46, 58) <= 4; angryBirdLarge(46, 59) <= 4; angryBirdLarge(46, 60) <= 4; angryBirdLarge(46, 61) <= 4; angryBirdLarge(46, 62) <= 4; angryBirdLarge(46, 63) <= 4; angryBirdLarge(46, 64) <= 4; angryBirdLarge(46, 65) <= 4; angryBirdLarge(46, 66) <= 4; angryBirdLarge(46, 67) <= 4; angryBirdLarge(46, 68) <= 4; angryBirdLarge(46, 69) <= 4; angryBirdLarge(46, 70) <= 4; angryBirdLarge(46, 71) <= 4; angryBirdLarge(46, 72) <= 4; angryBirdLarge(46, 73) <= 4; angryBirdLarge(46, 74) <= 4; angryBirdLarge(46, 75) <= 4; angryBirdLarge(46, 76) <= 4; angryBirdLarge(46, 77) <= 4; angryBirdLarge(46, 78) <= 4; angryBirdLarge(46, 79) <= 4; angryBirdLarge(46, 80) <= 4; angryBirdLarge(46, 81) <= 4; angryBirdLarge(46, 82) <= 4; angryBirdLarge(46, 83) <= 4; angryBirdLarge(46, 84) <= 4; angryBirdLarge(46, 85) <= 4; angryBirdLarge(46, 86) <= 4; angryBirdLarge(46, 87) <= 4; angryBirdLarge(46, 88) <= 4; angryBirdLarge(46, 89) <= 4; angryBirdLarge(46, 90) <= 4; angryBirdLarge(46, 91) <= 4; angryBirdLarge(46, 92) <= 4; angryBirdLarge(46, 93) <= 4; angryBirdLarge(46, 94) <= 4; angryBirdLarge(46, 95) <= 4; angryBirdLarge(46, 96) <= 4; angryBirdLarge(46, 97) <= 4; angryBirdLarge(46, 98) <= 4; angryBirdLarge(46, 99) <= 4; angryBirdLarge(46, 100) <= 4; angryBirdLarge(46, 101) <= 4; angryBirdLarge(46, 102) <= 4; angryBirdLarge(46, 103) <= 4; angryBirdLarge(46, 104) <= 4; angryBirdLarge(46, 105) <= 4; angryBirdLarge(46, 106) <= 4; angryBirdLarge(46, 107) <= 4; angryBirdLarge(46, 108) <= 4; angryBirdLarge(46, 109) <= 4; angryBirdLarge(46, 110) <= 4; angryBirdLarge(46, 111) <= 4; angryBirdLarge(46, 112) <= 4; angryBirdLarge(46, 113) <= 4; angryBirdLarge(46, 114) <= 4; angryBirdLarge(46, 115) <= 4; angryBirdLarge(46, 116) <= 4; angryBirdLarge(46, 117) <= 4; angryBirdLarge(46, 118) <= 4; angryBirdLarge(46, 119) <= 4; angryBirdLarge(46, 120) <= 4; angryBirdLarge(46, 121) <= 4; angryBirdLarge(46, 122) <= 4; angryBirdLarge(46, 123) <= 4; angryBirdLarge(46, 124) <= 4; angryBirdLarge(46, 125) <= 4; angryBirdLarge(46, 126) <= 5; angryBirdLarge(46, 127) <= 5; angryBirdLarge(46, 128) <= 5; angryBirdLarge(46, 129) <= 5; angryBirdLarge(46, 130) <= 5; angryBirdLarge(46, 131) <= 5; angryBirdLarge(46, 132) <= 0; angryBirdLarge(46, 133) <= 0; angryBirdLarge(46, 134) <= 0; angryBirdLarge(46, 135) <= 0; angryBirdLarge(46, 136) <= 0; angryBirdLarge(46, 137) <= 0; angryBirdLarge(46, 138) <= 0; angryBirdLarge(46, 139) <= 0; angryBirdLarge(46, 140) <= 0; angryBirdLarge(46, 141) <= 0; angryBirdLarge(46, 142) <= 0; angryBirdLarge(46, 143) <= 0; angryBirdLarge(46, 144) <= 0; angryBirdLarge(46, 145) <= 0; angryBirdLarge(46, 146) <= 0; angryBirdLarge(46, 147) <= 0; angryBirdLarge(46, 148) <= 0; angryBirdLarge(46, 149) <= 0; 
angryBirdLarge(47, 0) <= 0; angryBirdLarge(47, 1) <= 0; angryBirdLarge(47, 2) <= 0; angryBirdLarge(47, 3) <= 0; angryBirdLarge(47, 4) <= 0; angryBirdLarge(47, 5) <= 0; angryBirdLarge(47, 6) <= 0; angryBirdLarge(47, 7) <= 0; angryBirdLarge(47, 8) <= 0; angryBirdLarge(47, 9) <= 0; angryBirdLarge(47, 10) <= 0; angryBirdLarge(47, 11) <= 0; angryBirdLarge(47, 12) <= 0; angryBirdLarge(47, 13) <= 0; angryBirdLarge(47, 14) <= 0; angryBirdLarge(47, 15) <= 0; angryBirdLarge(47, 16) <= 0; angryBirdLarge(47, 17) <= 0; angryBirdLarge(47, 18) <= 0; angryBirdLarge(47, 19) <= 0; angryBirdLarge(47, 20) <= 0; angryBirdLarge(47, 21) <= 0; angryBirdLarge(47, 22) <= 0; angryBirdLarge(47, 23) <= 0; angryBirdLarge(47, 24) <= 0; angryBirdLarge(47, 25) <= 0; angryBirdLarge(47, 26) <= 0; angryBirdLarge(47, 27) <= 0; angryBirdLarge(47, 28) <= 0; angryBirdLarge(47, 29) <= 0; angryBirdLarge(47, 30) <= 0; angryBirdLarge(47, 31) <= 0; angryBirdLarge(47, 32) <= 0; angryBirdLarge(47, 33) <= 0; angryBirdLarge(47, 34) <= 0; angryBirdLarge(47, 35) <= 0; angryBirdLarge(47, 36) <= 5; angryBirdLarge(47, 37) <= 5; angryBirdLarge(47, 38) <= 5; angryBirdLarge(47, 39) <= 5; angryBirdLarge(47, 40) <= 5; angryBirdLarge(47, 41) <= 5; angryBirdLarge(47, 42) <= 4; angryBirdLarge(47, 43) <= 4; angryBirdLarge(47, 44) <= 4; angryBirdLarge(47, 45) <= 4; angryBirdLarge(47, 46) <= 4; angryBirdLarge(47, 47) <= 4; angryBirdLarge(47, 48) <= 4; angryBirdLarge(47, 49) <= 4; angryBirdLarge(47, 50) <= 4; angryBirdLarge(47, 51) <= 4; angryBirdLarge(47, 52) <= 4; angryBirdLarge(47, 53) <= 4; angryBirdLarge(47, 54) <= 4; angryBirdLarge(47, 55) <= 4; angryBirdLarge(47, 56) <= 4; angryBirdLarge(47, 57) <= 4; angryBirdLarge(47, 58) <= 4; angryBirdLarge(47, 59) <= 4; angryBirdLarge(47, 60) <= 4; angryBirdLarge(47, 61) <= 4; angryBirdLarge(47, 62) <= 4; angryBirdLarge(47, 63) <= 4; angryBirdLarge(47, 64) <= 4; angryBirdLarge(47, 65) <= 4; angryBirdLarge(47, 66) <= 4; angryBirdLarge(47, 67) <= 4; angryBirdLarge(47, 68) <= 4; angryBirdLarge(47, 69) <= 4; angryBirdLarge(47, 70) <= 4; angryBirdLarge(47, 71) <= 4; angryBirdLarge(47, 72) <= 4; angryBirdLarge(47, 73) <= 4; angryBirdLarge(47, 74) <= 4; angryBirdLarge(47, 75) <= 4; angryBirdLarge(47, 76) <= 4; angryBirdLarge(47, 77) <= 4; angryBirdLarge(47, 78) <= 4; angryBirdLarge(47, 79) <= 4; angryBirdLarge(47, 80) <= 4; angryBirdLarge(47, 81) <= 4; angryBirdLarge(47, 82) <= 4; angryBirdLarge(47, 83) <= 4; angryBirdLarge(47, 84) <= 4; angryBirdLarge(47, 85) <= 4; angryBirdLarge(47, 86) <= 4; angryBirdLarge(47, 87) <= 4; angryBirdLarge(47, 88) <= 4; angryBirdLarge(47, 89) <= 4; angryBirdLarge(47, 90) <= 4; angryBirdLarge(47, 91) <= 4; angryBirdLarge(47, 92) <= 4; angryBirdLarge(47, 93) <= 4; angryBirdLarge(47, 94) <= 4; angryBirdLarge(47, 95) <= 4; angryBirdLarge(47, 96) <= 4; angryBirdLarge(47, 97) <= 4; angryBirdLarge(47, 98) <= 4; angryBirdLarge(47, 99) <= 4; angryBirdLarge(47, 100) <= 4; angryBirdLarge(47, 101) <= 4; angryBirdLarge(47, 102) <= 4; angryBirdLarge(47, 103) <= 4; angryBirdLarge(47, 104) <= 4; angryBirdLarge(47, 105) <= 4; angryBirdLarge(47, 106) <= 4; angryBirdLarge(47, 107) <= 4; angryBirdLarge(47, 108) <= 4; angryBirdLarge(47, 109) <= 4; angryBirdLarge(47, 110) <= 4; angryBirdLarge(47, 111) <= 4; angryBirdLarge(47, 112) <= 4; angryBirdLarge(47, 113) <= 4; angryBirdLarge(47, 114) <= 4; angryBirdLarge(47, 115) <= 4; angryBirdLarge(47, 116) <= 4; angryBirdLarge(47, 117) <= 4; angryBirdLarge(47, 118) <= 4; angryBirdLarge(47, 119) <= 4; angryBirdLarge(47, 120) <= 4; angryBirdLarge(47, 121) <= 4; angryBirdLarge(47, 122) <= 4; angryBirdLarge(47, 123) <= 4; angryBirdLarge(47, 124) <= 4; angryBirdLarge(47, 125) <= 4; angryBirdLarge(47, 126) <= 5; angryBirdLarge(47, 127) <= 5; angryBirdLarge(47, 128) <= 5; angryBirdLarge(47, 129) <= 5; angryBirdLarge(47, 130) <= 5; angryBirdLarge(47, 131) <= 5; angryBirdLarge(47, 132) <= 0; angryBirdLarge(47, 133) <= 0; angryBirdLarge(47, 134) <= 0; angryBirdLarge(47, 135) <= 0; angryBirdLarge(47, 136) <= 0; angryBirdLarge(47, 137) <= 0; angryBirdLarge(47, 138) <= 0; angryBirdLarge(47, 139) <= 0; angryBirdLarge(47, 140) <= 0; angryBirdLarge(47, 141) <= 0; angryBirdLarge(47, 142) <= 0; angryBirdLarge(47, 143) <= 0; angryBirdLarge(47, 144) <= 0; angryBirdLarge(47, 145) <= 0; angryBirdLarge(47, 146) <= 0; angryBirdLarge(47, 147) <= 0; angryBirdLarge(47, 148) <= 0; angryBirdLarge(47, 149) <= 0; 
angryBirdLarge(48, 0) <= 0; angryBirdLarge(48, 1) <= 0; angryBirdLarge(48, 2) <= 0; angryBirdLarge(48, 3) <= 0; angryBirdLarge(48, 4) <= 0; angryBirdLarge(48, 5) <= 0; angryBirdLarge(48, 6) <= 0; angryBirdLarge(48, 7) <= 0; angryBirdLarge(48, 8) <= 0; angryBirdLarge(48, 9) <= 0; angryBirdLarge(48, 10) <= 0; angryBirdLarge(48, 11) <= 0; angryBirdLarge(48, 12) <= 0; angryBirdLarge(48, 13) <= 0; angryBirdLarge(48, 14) <= 0; angryBirdLarge(48, 15) <= 0; angryBirdLarge(48, 16) <= 0; angryBirdLarge(48, 17) <= 0; angryBirdLarge(48, 18) <= 0; angryBirdLarge(48, 19) <= 0; angryBirdLarge(48, 20) <= 0; angryBirdLarge(48, 21) <= 0; angryBirdLarge(48, 22) <= 0; angryBirdLarge(48, 23) <= 0; angryBirdLarge(48, 24) <= 0; angryBirdLarge(48, 25) <= 0; angryBirdLarge(48, 26) <= 0; angryBirdLarge(48, 27) <= 0; angryBirdLarge(48, 28) <= 0; angryBirdLarge(48, 29) <= 0; angryBirdLarge(48, 30) <= 0; angryBirdLarge(48, 31) <= 0; angryBirdLarge(48, 32) <= 0; angryBirdLarge(48, 33) <= 0; angryBirdLarge(48, 34) <= 0; angryBirdLarge(48, 35) <= 0; angryBirdLarge(48, 36) <= 5; angryBirdLarge(48, 37) <= 5; angryBirdLarge(48, 38) <= 5; angryBirdLarge(48, 39) <= 5; angryBirdLarge(48, 40) <= 5; angryBirdLarge(48, 41) <= 5; angryBirdLarge(48, 42) <= 4; angryBirdLarge(48, 43) <= 4; angryBirdLarge(48, 44) <= 4; angryBirdLarge(48, 45) <= 4; angryBirdLarge(48, 46) <= 4; angryBirdLarge(48, 47) <= 4; angryBirdLarge(48, 48) <= 4; angryBirdLarge(48, 49) <= 4; angryBirdLarge(48, 50) <= 4; angryBirdLarge(48, 51) <= 4; angryBirdLarge(48, 52) <= 4; angryBirdLarge(48, 53) <= 4; angryBirdLarge(48, 54) <= 4; angryBirdLarge(48, 55) <= 4; angryBirdLarge(48, 56) <= 4; angryBirdLarge(48, 57) <= 4; angryBirdLarge(48, 58) <= 4; angryBirdLarge(48, 59) <= 4; angryBirdLarge(48, 60) <= 4; angryBirdLarge(48, 61) <= 4; angryBirdLarge(48, 62) <= 4; angryBirdLarge(48, 63) <= 4; angryBirdLarge(48, 64) <= 4; angryBirdLarge(48, 65) <= 4; angryBirdLarge(48, 66) <= 4; angryBirdLarge(48, 67) <= 4; angryBirdLarge(48, 68) <= 4; angryBirdLarge(48, 69) <= 4; angryBirdLarge(48, 70) <= 4; angryBirdLarge(48, 71) <= 4; angryBirdLarge(48, 72) <= 4; angryBirdLarge(48, 73) <= 4; angryBirdLarge(48, 74) <= 4; angryBirdLarge(48, 75) <= 4; angryBirdLarge(48, 76) <= 4; angryBirdLarge(48, 77) <= 4; angryBirdLarge(48, 78) <= 4; angryBirdLarge(48, 79) <= 4; angryBirdLarge(48, 80) <= 4; angryBirdLarge(48, 81) <= 4; angryBirdLarge(48, 82) <= 4; angryBirdLarge(48, 83) <= 4; angryBirdLarge(48, 84) <= 4; angryBirdLarge(48, 85) <= 4; angryBirdLarge(48, 86) <= 4; angryBirdLarge(48, 87) <= 4; angryBirdLarge(48, 88) <= 4; angryBirdLarge(48, 89) <= 4; angryBirdLarge(48, 90) <= 4; angryBirdLarge(48, 91) <= 4; angryBirdLarge(48, 92) <= 4; angryBirdLarge(48, 93) <= 4; angryBirdLarge(48, 94) <= 4; angryBirdLarge(48, 95) <= 4; angryBirdLarge(48, 96) <= 4; angryBirdLarge(48, 97) <= 4; angryBirdLarge(48, 98) <= 4; angryBirdLarge(48, 99) <= 4; angryBirdLarge(48, 100) <= 4; angryBirdLarge(48, 101) <= 4; angryBirdLarge(48, 102) <= 4; angryBirdLarge(48, 103) <= 4; angryBirdLarge(48, 104) <= 4; angryBirdLarge(48, 105) <= 4; angryBirdLarge(48, 106) <= 4; angryBirdLarge(48, 107) <= 4; angryBirdLarge(48, 108) <= 4; angryBirdLarge(48, 109) <= 4; angryBirdLarge(48, 110) <= 4; angryBirdLarge(48, 111) <= 4; angryBirdLarge(48, 112) <= 4; angryBirdLarge(48, 113) <= 4; angryBirdLarge(48, 114) <= 4; angryBirdLarge(48, 115) <= 4; angryBirdLarge(48, 116) <= 4; angryBirdLarge(48, 117) <= 4; angryBirdLarge(48, 118) <= 4; angryBirdLarge(48, 119) <= 4; angryBirdLarge(48, 120) <= 4; angryBirdLarge(48, 121) <= 4; angryBirdLarge(48, 122) <= 4; angryBirdLarge(48, 123) <= 4; angryBirdLarge(48, 124) <= 4; angryBirdLarge(48, 125) <= 4; angryBirdLarge(48, 126) <= 4; angryBirdLarge(48, 127) <= 4; angryBirdLarge(48, 128) <= 4; angryBirdLarge(48, 129) <= 4; angryBirdLarge(48, 130) <= 4; angryBirdLarge(48, 131) <= 4; angryBirdLarge(48, 132) <= 5; angryBirdLarge(48, 133) <= 5; angryBirdLarge(48, 134) <= 5; angryBirdLarge(48, 135) <= 5; angryBirdLarge(48, 136) <= 5; angryBirdLarge(48, 137) <= 5; angryBirdLarge(48, 138) <= 0; angryBirdLarge(48, 139) <= 0; angryBirdLarge(48, 140) <= 0; angryBirdLarge(48, 141) <= 0; angryBirdLarge(48, 142) <= 0; angryBirdLarge(48, 143) <= 0; angryBirdLarge(48, 144) <= 0; angryBirdLarge(48, 145) <= 0; angryBirdLarge(48, 146) <= 0; angryBirdLarge(48, 147) <= 0; angryBirdLarge(48, 148) <= 0; angryBirdLarge(48, 149) <= 0; 
angryBirdLarge(49, 0) <= 0; angryBirdLarge(49, 1) <= 0; angryBirdLarge(49, 2) <= 0; angryBirdLarge(49, 3) <= 0; angryBirdLarge(49, 4) <= 0; angryBirdLarge(49, 5) <= 0; angryBirdLarge(49, 6) <= 0; angryBirdLarge(49, 7) <= 0; angryBirdLarge(49, 8) <= 0; angryBirdLarge(49, 9) <= 0; angryBirdLarge(49, 10) <= 0; angryBirdLarge(49, 11) <= 0; angryBirdLarge(49, 12) <= 0; angryBirdLarge(49, 13) <= 0; angryBirdLarge(49, 14) <= 0; angryBirdLarge(49, 15) <= 0; angryBirdLarge(49, 16) <= 0; angryBirdLarge(49, 17) <= 0; angryBirdLarge(49, 18) <= 0; angryBirdLarge(49, 19) <= 0; angryBirdLarge(49, 20) <= 0; angryBirdLarge(49, 21) <= 0; angryBirdLarge(49, 22) <= 0; angryBirdLarge(49, 23) <= 0; angryBirdLarge(49, 24) <= 0; angryBirdLarge(49, 25) <= 0; angryBirdLarge(49, 26) <= 0; angryBirdLarge(49, 27) <= 0; angryBirdLarge(49, 28) <= 0; angryBirdLarge(49, 29) <= 0; angryBirdLarge(49, 30) <= 0; angryBirdLarge(49, 31) <= 0; angryBirdLarge(49, 32) <= 0; angryBirdLarge(49, 33) <= 0; angryBirdLarge(49, 34) <= 0; angryBirdLarge(49, 35) <= 0; angryBirdLarge(49, 36) <= 5; angryBirdLarge(49, 37) <= 5; angryBirdLarge(49, 38) <= 5; angryBirdLarge(49, 39) <= 5; angryBirdLarge(49, 40) <= 5; angryBirdLarge(49, 41) <= 5; angryBirdLarge(49, 42) <= 4; angryBirdLarge(49, 43) <= 4; angryBirdLarge(49, 44) <= 4; angryBirdLarge(49, 45) <= 4; angryBirdLarge(49, 46) <= 4; angryBirdLarge(49, 47) <= 4; angryBirdLarge(49, 48) <= 4; angryBirdLarge(49, 49) <= 4; angryBirdLarge(49, 50) <= 4; angryBirdLarge(49, 51) <= 4; angryBirdLarge(49, 52) <= 4; angryBirdLarge(49, 53) <= 4; angryBirdLarge(49, 54) <= 4; angryBirdLarge(49, 55) <= 4; angryBirdLarge(49, 56) <= 4; angryBirdLarge(49, 57) <= 4; angryBirdLarge(49, 58) <= 4; angryBirdLarge(49, 59) <= 4; angryBirdLarge(49, 60) <= 4; angryBirdLarge(49, 61) <= 4; angryBirdLarge(49, 62) <= 4; angryBirdLarge(49, 63) <= 4; angryBirdLarge(49, 64) <= 4; angryBirdLarge(49, 65) <= 4; angryBirdLarge(49, 66) <= 4; angryBirdLarge(49, 67) <= 4; angryBirdLarge(49, 68) <= 4; angryBirdLarge(49, 69) <= 4; angryBirdLarge(49, 70) <= 4; angryBirdLarge(49, 71) <= 4; angryBirdLarge(49, 72) <= 4; angryBirdLarge(49, 73) <= 4; angryBirdLarge(49, 74) <= 4; angryBirdLarge(49, 75) <= 4; angryBirdLarge(49, 76) <= 4; angryBirdLarge(49, 77) <= 4; angryBirdLarge(49, 78) <= 4; angryBirdLarge(49, 79) <= 4; angryBirdLarge(49, 80) <= 4; angryBirdLarge(49, 81) <= 4; angryBirdLarge(49, 82) <= 4; angryBirdLarge(49, 83) <= 4; angryBirdLarge(49, 84) <= 4; angryBirdLarge(49, 85) <= 4; angryBirdLarge(49, 86) <= 4; angryBirdLarge(49, 87) <= 4; angryBirdLarge(49, 88) <= 4; angryBirdLarge(49, 89) <= 4; angryBirdLarge(49, 90) <= 4; angryBirdLarge(49, 91) <= 4; angryBirdLarge(49, 92) <= 4; angryBirdLarge(49, 93) <= 4; angryBirdLarge(49, 94) <= 4; angryBirdLarge(49, 95) <= 4; angryBirdLarge(49, 96) <= 4; angryBirdLarge(49, 97) <= 4; angryBirdLarge(49, 98) <= 4; angryBirdLarge(49, 99) <= 4; angryBirdLarge(49, 100) <= 4; angryBirdLarge(49, 101) <= 4; angryBirdLarge(49, 102) <= 4; angryBirdLarge(49, 103) <= 4; angryBirdLarge(49, 104) <= 4; angryBirdLarge(49, 105) <= 4; angryBirdLarge(49, 106) <= 4; angryBirdLarge(49, 107) <= 4; angryBirdLarge(49, 108) <= 4; angryBirdLarge(49, 109) <= 4; angryBirdLarge(49, 110) <= 4; angryBirdLarge(49, 111) <= 4; angryBirdLarge(49, 112) <= 4; angryBirdLarge(49, 113) <= 4; angryBirdLarge(49, 114) <= 4; angryBirdLarge(49, 115) <= 4; angryBirdLarge(49, 116) <= 4; angryBirdLarge(49, 117) <= 4; angryBirdLarge(49, 118) <= 4; angryBirdLarge(49, 119) <= 4; angryBirdLarge(49, 120) <= 4; angryBirdLarge(49, 121) <= 4; angryBirdLarge(49, 122) <= 4; angryBirdLarge(49, 123) <= 4; angryBirdLarge(49, 124) <= 4; angryBirdLarge(49, 125) <= 4; angryBirdLarge(49, 126) <= 4; angryBirdLarge(49, 127) <= 4; angryBirdLarge(49, 128) <= 4; angryBirdLarge(49, 129) <= 4; angryBirdLarge(49, 130) <= 4; angryBirdLarge(49, 131) <= 4; angryBirdLarge(49, 132) <= 5; angryBirdLarge(49, 133) <= 5; angryBirdLarge(49, 134) <= 5; angryBirdLarge(49, 135) <= 5; angryBirdLarge(49, 136) <= 5; angryBirdLarge(49, 137) <= 5; angryBirdLarge(49, 138) <= 0; angryBirdLarge(49, 139) <= 0; angryBirdLarge(49, 140) <= 0; angryBirdLarge(49, 141) <= 0; angryBirdLarge(49, 142) <= 0; angryBirdLarge(49, 143) <= 0; angryBirdLarge(49, 144) <= 0; angryBirdLarge(49, 145) <= 0; angryBirdLarge(49, 146) <= 0; angryBirdLarge(49, 147) <= 0; angryBirdLarge(49, 148) <= 0; angryBirdLarge(49, 149) <= 0; 
angryBirdLarge(50, 0) <= 0; angryBirdLarge(50, 1) <= 0; angryBirdLarge(50, 2) <= 0; angryBirdLarge(50, 3) <= 0; angryBirdLarge(50, 4) <= 0; angryBirdLarge(50, 5) <= 0; angryBirdLarge(50, 6) <= 0; angryBirdLarge(50, 7) <= 0; angryBirdLarge(50, 8) <= 0; angryBirdLarge(50, 9) <= 0; angryBirdLarge(50, 10) <= 0; angryBirdLarge(50, 11) <= 0; angryBirdLarge(50, 12) <= 0; angryBirdLarge(50, 13) <= 0; angryBirdLarge(50, 14) <= 0; angryBirdLarge(50, 15) <= 0; angryBirdLarge(50, 16) <= 0; angryBirdLarge(50, 17) <= 0; angryBirdLarge(50, 18) <= 0; angryBirdLarge(50, 19) <= 0; angryBirdLarge(50, 20) <= 0; angryBirdLarge(50, 21) <= 0; angryBirdLarge(50, 22) <= 0; angryBirdLarge(50, 23) <= 0; angryBirdLarge(50, 24) <= 0; angryBirdLarge(50, 25) <= 0; angryBirdLarge(50, 26) <= 0; angryBirdLarge(50, 27) <= 0; angryBirdLarge(50, 28) <= 0; angryBirdLarge(50, 29) <= 0; angryBirdLarge(50, 30) <= 0; angryBirdLarge(50, 31) <= 0; angryBirdLarge(50, 32) <= 0; angryBirdLarge(50, 33) <= 0; angryBirdLarge(50, 34) <= 0; angryBirdLarge(50, 35) <= 0; angryBirdLarge(50, 36) <= 5; angryBirdLarge(50, 37) <= 5; angryBirdLarge(50, 38) <= 5; angryBirdLarge(50, 39) <= 5; angryBirdLarge(50, 40) <= 5; angryBirdLarge(50, 41) <= 5; angryBirdLarge(50, 42) <= 4; angryBirdLarge(50, 43) <= 4; angryBirdLarge(50, 44) <= 4; angryBirdLarge(50, 45) <= 4; angryBirdLarge(50, 46) <= 4; angryBirdLarge(50, 47) <= 4; angryBirdLarge(50, 48) <= 4; angryBirdLarge(50, 49) <= 4; angryBirdLarge(50, 50) <= 4; angryBirdLarge(50, 51) <= 4; angryBirdLarge(50, 52) <= 4; angryBirdLarge(50, 53) <= 4; angryBirdLarge(50, 54) <= 4; angryBirdLarge(50, 55) <= 4; angryBirdLarge(50, 56) <= 4; angryBirdLarge(50, 57) <= 4; angryBirdLarge(50, 58) <= 4; angryBirdLarge(50, 59) <= 4; angryBirdLarge(50, 60) <= 4; angryBirdLarge(50, 61) <= 4; angryBirdLarge(50, 62) <= 4; angryBirdLarge(50, 63) <= 4; angryBirdLarge(50, 64) <= 4; angryBirdLarge(50, 65) <= 4; angryBirdLarge(50, 66) <= 4; angryBirdLarge(50, 67) <= 4; angryBirdLarge(50, 68) <= 4; angryBirdLarge(50, 69) <= 4; angryBirdLarge(50, 70) <= 4; angryBirdLarge(50, 71) <= 4; angryBirdLarge(50, 72) <= 4; angryBirdLarge(50, 73) <= 4; angryBirdLarge(50, 74) <= 4; angryBirdLarge(50, 75) <= 4; angryBirdLarge(50, 76) <= 4; angryBirdLarge(50, 77) <= 4; angryBirdLarge(50, 78) <= 4; angryBirdLarge(50, 79) <= 4; angryBirdLarge(50, 80) <= 4; angryBirdLarge(50, 81) <= 4; angryBirdLarge(50, 82) <= 4; angryBirdLarge(50, 83) <= 4; angryBirdLarge(50, 84) <= 4; angryBirdLarge(50, 85) <= 4; angryBirdLarge(50, 86) <= 4; angryBirdLarge(50, 87) <= 4; angryBirdLarge(50, 88) <= 4; angryBirdLarge(50, 89) <= 4; angryBirdLarge(50, 90) <= 4; angryBirdLarge(50, 91) <= 4; angryBirdLarge(50, 92) <= 4; angryBirdLarge(50, 93) <= 4; angryBirdLarge(50, 94) <= 4; angryBirdLarge(50, 95) <= 4; angryBirdLarge(50, 96) <= 4; angryBirdLarge(50, 97) <= 4; angryBirdLarge(50, 98) <= 4; angryBirdLarge(50, 99) <= 4; angryBirdLarge(50, 100) <= 4; angryBirdLarge(50, 101) <= 4; angryBirdLarge(50, 102) <= 4; angryBirdLarge(50, 103) <= 4; angryBirdLarge(50, 104) <= 4; angryBirdLarge(50, 105) <= 4; angryBirdLarge(50, 106) <= 4; angryBirdLarge(50, 107) <= 4; angryBirdLarge(50, 108) <= 4; angryBirdLarge(50, 109) <= 4; angryBirdLarge(50, 110) <= 4; angryBirdLarge(50, 111) <= 4; angryBirdLarge(50, 112) <= 4; angryBirdLarge(50, 113) <= 4; angryBirdLarge(50, 114) <= 4; angryBirdLarge(50, 115) <= 4; angryBirdLarge(50, 116) <= 4; angryBirdLarge(50, 117) <= 4; angryBirdLarge(50, 118) <= 4; angryBirdLarge(50, 119) <= 4; angryBirdLarge(50, 120) <= 4; angryBirdLarge(50, 121) <= 4; angryBirdLarge(50, 122) <= 4; angryBirdLarge(50, 123) <= 4; angryBirdLarge(50, 124) <= 4; angryBirdLarge(50, 125) <= 4; angryBirdLarge(50, 126) <= 4; angryBirdLarge(50, 127) <= 4; angryBirdLarge(50, 128) <= 4; angryBirdLarge(50, 129) <= 4; angryBirdLarge(50, 130) <= 4; angryBirdLarge(50, 131) <= 4; angryBirdLarge(50, 132) <= 5; angryBirdLarge(50, 133) <= 5; angryBirdLarge(50, 134) <= 5; angryBirdLarge(50, 135) <= 5; angryBirdLarge(50, 136) <= 5; angryBirdLarge(50, 137) <= 5; angryBirdLarge(50, 138) <= 0; angryBirdLarge(50, 139) <= 0; angryBirdLarge(50, 140) <= 0; angryBirdLarge(50, 141) <= 0; angryBirdLarge(50, 142) <= 0; angryBirdLarge(50, 143) <= 0; angryBirdLarge(50, 144) <= 0; angryBirdLarge(50, 145) <= 0; angryBirdLarge(50, 146) <= 0; angryBirdLarge(50, 147) <= 0; angryBirdLarge(50, 148) <= 0; angryBirdLarge(50, 149) <= 0; 
angryBirdLarge(51, 0) <= 0; angryBirdLarge(51, 1) <= 0; angryBirdLarge(51, 2) <= 0; angryBirdLarge(51, 3) <= 0; angryBirdLarge(51, 4) <= 0; angryBirdLarge(51, 5) <= 0; angryBirdLarge(51, 6) <= 0; angryBirdLarge(51, 7) <= 0; angryBirdLarge(51, 8) <= 0; angryBirdLarge(51, 9) <= 0; angryBirdLarge(51, 10) <= 0; angryBirdLarge(51, 11) <= 0; angryBirdLarge(51, 12) <= 0; angryBirdLarge(51, 13) <= 0; angryBirdLarge(51, 14) <= 0; angryBirdLarge(51, 15) <= 0; angryBirdLarge(51, 16) <= 0; angryBirdLarge(51, 17) <= 0; angryBirdLarge(51, 18) <= 0; angryBirdLarge(51, 19) <= 0; angryBirdLarge(51, 20) <= 0; angryBirdLarge(51, 21) <= 0; angryBirdLarge(51, 22) <= 0; angryBirdLarge(51, 23) <= 0; angryBirdLarge(51, 24) <= 0; angryBirdLarge(51, 25) <= 0; angryBirdLarge(51, 26) <= 0; angryBirdLarge(51, 27) <= 0; angryBirdLarge(51, 28) <= 0; angryBirdLarge(51, 29) <= 0; angryBirdLarge(51, 30) <= 0; angryBirdLarge(51, 31) <= 0; angryBirdLarge(51, 32) <= 0; angryBirdLarge(51, 33) <= 0; angryBirdLarge(51, 34) <= 0; angryBirdLarge(51, 35) <= 0; angryBirdLarge(51, 36) <= 5; angryBirdLarge(51, 37) <= 5; angryBirdLarge(51, 38) <= 5; angryBirdLarge(51, 39) <= 5; angryBirdLarge(51, 40) <= 5; angryBirdLarge(51, 41) <= 5; angryBirdLarge(51, 42) <= 4; angryBirdLarge(51, 43) <= 4; angryBirdLarge(51, 44) <= 4; angryBirdLarge(51, 45) <= 4; angryBirdLarge(51, 46) <= 4; angryBirdLarge(51, 47) <= 4; angryBirdLarge(51, 48) <= 4; angryBirdLarge(51, 49) <= 4; angryBirdLarge(51, 50) <= 4; angryBirdLarge(51, 51) <= 4; angryBirdLarge(51, 52) <= 4; angryBirdLarge(51, 53) <= 4; angryBirdLarge(51, 54) <= 4; angryBirdLarge(51, 55) <= 4; angryBirdLarge(51, 56) <= 4; angryBirdLarge(51, 57) <= 4; angryBirdLarge(51, 58) <= 4; angryBirdLarge(51, 59) <= 4; angryBirdLarge(51, 60) <= 4; angryBirdLarge(51, 61) <= 4; angryBirdLarge(51, 62) <= 4; angryBirdLarge(51, 63) <= 4; angryBirdLarge(51, 64) <= 4; angryBirdLarge(51, 65) <= 4; angryBirdLarge(51, 66) <= 4; angryBirdLarge(51, 67) <= 4; angryBirdLarge(51, 68) <= 4; angryBirdLarge(51, 69) <= 4; angryBirdLarge(51, 70) <= 4; angryBirdLarge(51, 71) <= 4; angryBirdLarge(51, 72) <= 4; angryBirdLarge(51, 73) <= 4; angryBirdLarge(51, 74) <= 4; angryBirdLarge(51, 75) <= 4; angryBirdLarge(51, 76) <= 4; angryBirdLarge(51, 77) <= 4; angryBirdLarge(51, 78) <= 4; angryBirdLarge(51, 79) <= 4; angryBirdLarge(51, 80) <= 4; angryBirdLarge(51, 81) <= 4; angryBirdLarge(51, 82) <= 4; angryBirdLarge(51, 83) <= 4; angryBirdLarge(51, 84) <= 4; angryBirdLarge(51, 85) <= 4; angryBirdLarge(51, 86) <= 4; angryBirdLarge(51, 87) <= 4; angryBirdLarge(51, 88) <= 4; angryBirdLarge(51, 89) <= 4; angryBirdLarge(51, 90) <= 4; angryBirdLarge(51, 91) <= 4; angryBirdLarge(51, 92) <= 4; angryBirdLarge(51, 93) <= 4; angryBirdLarge(51, 94) <= 4; angryBirdLarge(51, 95) <= 4; angryBirdLarge(51, 96) <= 4; angryBirdLarge(51, 97) <= 4; angryBirdLarge(51, 98) <= 4; angryBirdLarge(51, 99) <= 4; angryBirdLarge(51, 100) <= 4; angryBirdLarge(51, 101) <= 4; angryBirdLarge(51, 102) <= 4; angryBirdLarge(51, 103) <= 4; angryBirdLarge(51, 104) <= 4; angryBirdLarge(51, 105) <= 4; angryBirdLarge(51, 106) <= 4; angryBirdLarge(51, 107) <= 4; angryBirdLarge(51, 108) <= 4; angryBirdLarge(51, 109) <= 4; angryBirdLarge(51, 110) <= 4; angryBirdLarge(51, 111) <= 4; angryBirdLarge(51, 112) <= 4; angryBirdLarge(51, 113) <= 4; angryBirdLarge(51, 114) <= 4; angryBirdLarge(51, 115) <= 4; angryBirdLarge(51, 116) <= 4; angryBirdLarge(51, 117) <= 4; angryBirdLarge(51, 118) <= 4; angryBirdLarge(51, 119) <= 4; angryBirdLarge(51, 120) <= 4; angryBirdLarge(51, 121) <= 4; angryBirdLarge(51, 122) <= 4; angryBirdLarge(51, 123) <= 4; angryBirdLarge(51, 124) <= 4; angryBirdLarge(51, 125) <= 4; angryBirdLarge(51, 126) <= 4; angryBirdLarge(51, 127) <= 4; angryBirdLarge(51, 128) <= 4; angryBirdLarge(51, 129) <= 4; angryBirdLarge(51, 130) <= 4; angryBirdLarge(51, 131) <= 4; angryBirdLarge(51, 132) <= 5; angryBirdLarge(51, 133) <= 5; angryBirdLarge(51, 134) <= 5; angryBirdLarge(51, 135) <= 5; angryBirdLarge(51, 136) <= 5; angryBirdLarge(51, 137) <= 5; angryBirdLarge(51, 138) <= 0; angryBirdLarge(51, 139) <= 0; angryBirdLarge(51, 140) <= 0; angryBirdLarge(51, 141) <= 0; angryBirdLarge(51, 142) <= 0; angryBirdLarge(51, 143) <= 0; angryBirdLarge(51, 144) <= 0; angryBirdLarge(51, 145) <= 0; angryBirdLarge(51, 146) <= 0; angryBirdLarge(51, 147) <= 0; angryBirdLarge(51, 148) <= 0; angryBirdLarge(51, 149) <= 0; 
angryBirdLarge(52, 0) <= 0; angryBirdLarge(52, 1) <= 0; angryBirdLarge(52, 2) <= 0; angryBirdLarge(52, 3) <= 0; angryBirdLarge(52, 4) <= 0; angryBirdLarge(52, 5) <= 0; angryBirdLarge(52, 6) <= 0; angryBirdLarge(52, 7) <= 0; angryBirdLarge(52, 8) <= 0; angryBirdLarge(52, 9) <= 0; angryBirdLarge(52, 10) <= 0; angryBirdLarge(52, 11) <= 0; angryBirdLarge(52, 12) <= 0; angryBirdLarge(52, 13) <= 0; angryBirdLarge(52, 14) <= 0; angryBirdLarge(52, 15) <= 0; angryBirdLarge(52, 16) <= 0; angryBirdLarge(52, 17) <= 0; angryBirdLarge(52, 18) <= 0; angryBirdLarge(52, 19) <= 0; angryBirdLarge(52, 20) <= 0; angryBirdLarge(52, 21) <= 0; angryBirdLarge(52, 22) <= 0; angryBirdLarge(52, 23) <= 0; angryBirdLarge(52, 24) <= 0; angryBirdLarge(52, 25) <= 0; angryBirdLarge(52, 26) <= 0; angryBirdLarge(52, 27) <= 0; angryBirdLarge(52, 28) <= 0; angryBirdLarge(52, 29) <= 0; angryBirdLarge(52, 30) <= 0; angryBirdLarge(52, 31) <= 0; angryBirdLarge(52, 32) <= 0; angryBirdLarge(52, 33) <= 0; angryBirdLarge(52, 34) <= 0; angryBirdLarge(52, 35) <= 0; angryBirdLarge(52, 36) <= 5; angryBirdLarge(52, 37) <= 5; angryBirdLarge(52, 38) <= 5; angryBirdLarge(52, 39) <= 5; angryBirdLarge(52, 40) <= 5; angryBirdLarge(52, 41) <= 5; angryBirdLarge(52, 42) <= 4; angryBirdLarge(52, 43) <= 4; angryBirdLarge(52, 44) <= 4; angryBirdLarge(52, 45) <= 4; angryBirdLarge(52, 46) <= 4; angryBirdLarge(52, 47) <= 4; angryBirdLarge(52, 48) <= 4; angryBirdLarge(52, 49) <= 4; angryBirdLarge(52, 50) <= 4; angryBirdLarge(52, 51) <= 4; angryBirdLarge(52, 52) <= 4; angryBirdLarge(52, 53) <= 4; angryBirdLarge(52, 54) <= 4; angryBirdLarge(52, 55) <= 4; angryBirdLarge(52, 56) <= 4; angryBirdLarge(52, 57) <= 4; angryBirdLarge(52, 58) <= 4; angryBirdLarge(52, 59) <= 4; angryBirdLarge(52, 60) <= 4; angryBirdLarge(52, 61) <= 4; angryBirdLarge(52, 62) <= 4; angryBirdLarge(52, 63) <= 4; angryBirdLarge(52, 64) <= 4; angryBirdLarge(52, 65) <= 4; angryBirdLarge(52, 66) <= 4; angryBirdLarge(52, 67) <= 4; angryBirdLarge(52, 68) <= 4; angryBirdLarge(52, 69) <= 4; angryBirdLarge(52, 70) <= 4; angryBirdLarge(52, 71) <= 4; angryBirdLarge(52, 72) <= 4; angryBirdLarge(52, 73) <= 4; angryBirdLarge(52, 74) <= 4; angryBirdLarge(52, 75) <= 4; angryBirdLarge(52, 76) <= 4; angryBirdLarge(52, 77) <= 4; angryBirdLarge(52, 78) <= 4; angryBirdLarge(52, 79) <= 4; angryBirdLarge(52, 80) <= 4; angryBirdLarge(52, 81) <= 4; angryBirdLarge(52, 82) <= 4; angryBirdLarge(52, 83) <= 4; angryBirdLarge(52, 84) <= 4; angryBirdLarge(52, 85) <= 4; angryBirdLarge(52, 86) <= 4; angryBirdLarge(52, 87) <= 4; angryBirdLarge(52, 88) <= 4; angryBirdLarge(52, 89) <= 4; angryBirdLarge(52, 90) <= 4; angryBirdLarge(52, 91) <= 4; angryBirdLarge(52, 92) <= 4; angryBirdLarge(52, 93) <= 4; angryBirdLarge(52, 94) <= 4; angryBirdLarge(52, 95) <= 4; angryBirdLarge(52, 96) <= 4; angryBirdLarge(52, 97) <= 4; angryBirdLarge(52, 98) <= 4; angryBirdLarge(52, 99) <= 4; angryBirdLarge(52, 100) <= 4; angryBirdLarge(52, 101) <= 4; angryBirdLarge(52, 102) <= 4; angryBirdLarge(52, 103) <= 4; angryBirdLarge(52, 104) <= 4; angryBirdLarge(52, 105) <= 4; angryBirdLarge(52, 106) <= 4; angryBirdLarge(52, 107) <= 4; angryBirdLarge(52, 108) <= 4; angryBirdLarge(52, 109) <= 4; angryBirdLarge(52, 110) <= 4; angryBirdLarge(52, 111) <= 4; angryBirdLarge(52, 112) <= 4; angryBirdLarge(52, 113) <= 4; angryBirdLarge(52, 114) <= 4; angryBirdLarge(52, 115) <= 4; angryBirdLarge(52, 116) <= 4; angryBirdLarge(52, 117) <= 4; angryBirdLarge(52, 118) <= 4; angryBirdLarge(52, 119) <= 4; angryBirdLarge(52, 120) <= 4; angryBirdLarge(52, 121) <= 4; angryBirdLarge(52, 122) <= 4; angryBirdLarge(52, 123) <= 4; angryBirdLarge(52, 124) <= 4; angryBirdLarge(52, 125) <= 4; angryBirdLarge(52, 126) <= 4; angryBirdLarge(52, 127) <= 4; angryBirdLarge(52, 128) <= 4; angryBirdLarge(52, 129) <= 4; angryBirdLarge(52, 130) <= 4; angryBirdLarge(52, 131) <= 4; angryBirdLarge(52, 132) <= 5; angryBirdLarge(52, 133) <= 5; angryBirdLarge(52, 134) <= 5; angryBirdLarge(52, 135) <= 5; angryBirdLarge(52, 136) <= 5; angryBirdLarge(52, 137) <= 5; angryBirdLarge(52, 138) <= 0; angryBirdLarge(52, 139) <= 0; angryBirdLarge(52, 140) <= 0; angryBirdLarge(52, 141) <= 0; angryBirdLarge(52, 142) <= 0; angryBirdLarge(52, 143) <= 0; angryBirdLarge(52, 144) <= 0; angryBirdLarge(52, 145) <= 0; angryBirdLarge(52, 146) <= 0; angryBirdLarge(52, 147) <= 0; angryBirdLarge(52, 148) <= 0; angryBirdLarge(52, 149) <= 0; 
angryBirdLarge(53, 0) <= 0; angryBirdLarge(53, 1) <= 0; angryBirdLarge(53, 2) <= 0; angryBirdLarge(53, 3) <= 0; angryBirdLarge(53, 4) <= 0; angryBirdLarge(53, 5) <= 0; angryBirdLarge(53, 6) <= 0; angryBirdLarge(53, 7) <= 0; angryBirdLarge(53, 8) <= 0; angryBirdLarge(53, 9) <= 0; angryBirdLarge(53, 10) <= 0; angryBirdLarge(53, 11) <= 0; angryBirdLarge(53, 12) <= 0; angryBirdLarge(53, 13) <= 0; angryBirdLarge(53, 14) <= 0; angryBirdLarge(53, 15) <= 0; angryBirdLarge(53, 16) <= 0; angryBirdLarge(53, 17) <= 0; angryBirdLarge(53, 18) <= 0; angryBirdLarge(53, 19) <= 0; angryBirdLarge(53, 20) <= 0; angryBirdLarge(53, 21) <= 0; angryBirdLarge(53, 22) <= 0; angryBirdLarge(53, 23) <= 0; angryBirdLarge(53, 24) <= 0; angryBirdLarge(53, 25) <= 0; angryBirdLarge(53, 26) <= 0; angryBirdLarge(53, 27) <= 0; angryBirdLarge(53, 28) <= 0; angryBirdLarge(53, 29) <= 0; angryBirdLarge(53, 30) <= 0; angryBirdLarge(53, 31) <= 0; angryBirdLarge(53, 32) <= 0; angryBirdLarge(53, 33) <= 0; angryBirdLarge(53, 34) <= 0; angryBirdLarge(53, 35) <= 0; angryBirdLarge(53, 36) <= 5; angryBirdLarge(53, 37) <= 5; angryBirdLarge(53, 38) <= 5; angryBirdLarge(53, 39) <= 5; angryBirdLarge(53, 40) <= 5; angryBirdLarge(53, 41) <= 5; angryBirdLarge(53, 42) <= 4; angryBirdLarge(53, 43) <= 4; angryBirdLarge(53, 44) <= 4; angryBirdLarge(53, 45) <= 4; angryBirdLarge(53, 46) <= 4; angryBirdLarge(53, 47) <= 4; angryBirdLarge(53, 48) <= 4; angryBirdLarge(53, 49) <= 4; angryBirdLarge(53, 50) <= 4; angryBirdLarge(53, 51) <= 4; angryBirdLarge(53, 52) <= 4; angryBirdLarge(53, 53) <= 4; angryBirdLarge(53, 54) <= 4; angryBirdLarge(53, 55) <= 4; angryBirdLarge(53, 56) <= 4; angryBirdLarge(53, 57) <= 4; angryBirdLarge(53, 58) <= 4; angryBirdLarge(53, 59) <= 4; angryBirdLarge(53, 60) <= 4; angryBirdLarge(53, 61) <= 4; angryBirdLarge(53, 62) <= 4; angryBirdLarge(53, 63) <= 4; angryBirdLarge(53, 64) <= 4; angryBirdLarge(53, 65) <= 4; angryBirdLarge(53, 66) <= 4; angryBirdLarge(53, 67) <= 4; angryBirdLarge(53, 68) <= 4; angryBirdLarge(53, 69) <= 4; angryBirdLarge(53, 70) <= 4; angryBirdLarge(53, 71) <= 4; angryBirdLarge(53, 72) <= 4; angryBirdLarge(53, 73) <= 4; angryBirdLarge(53, 74) <= 4; angryBirdLarge(53, 75) <= 4; angryBirdLarge(53, 76) <= 4; angryBirdLarge(53, 77) <= 4; angryBirdLarge(53, 78) <= 4; angryBirdLarge(53, 79) <= 4; angryBirdLarge(53, 80) <= 4; angryBirdLarge(53, 81) <= 4; angryBirdLarge(53, 82) <= 4; angryBirdLarge(53, 83) <= 4; angryBirdLarge(53, 84) <= 4; angryBirdLarge(53, 85) <= 4; angryBirdLarge(53, 86) <= 4; angryBirdLarge(53, 87) <= 4; angryBirdLarge(53, 88) <= 4; angryBirdLarge(53, 89) <= 4; angryBirdLarge(53, 90) <= 4; angryBirdLarge(53, 91) <= 4; angryBirdLarge(53, 92) <= 4; angryBirdLarge(53, 93) <= 4; angryBirdLarge(53, 94) <= 4; angryBirdLarge(53, 95) <= 4; angryBirdLarge(53, 96) <= 4; angryBirdLarge(53, 97) <= 4; angryBirdLarge(53, 98) <= 4; angryBirdLarge(53, 99) <= 4; angryBirdLarge(53, 100) <= 4; angryBirdLarge(53, 101) <= 4; angryBirdLarge(53, 102) <= 4; angryBirdLarge(53, 103) <= 4; angryBirdLarge(53, 104) <= 4; angryBirdLarge(53, 105) <= 4; angryBirdLarge(53, 106) <= 4; angryBirdLarge(53, 107) <= 4; angryBirdLarge(53, 108) <= 4; angryBirdLarge(53, 109) <= 4; angryBirdLarge(53, 110) <= 4; angryBirdLarge(53, 111) <= 4; angryBirdLarge(53, 112) <= 4; angryBirdLarge(53, 113) <= 4; angryBirdLarge(53, 114) <= 4; angryBirdLarge(53, 115) <= 4; angryBirdLarge(53, 116) <= 4; angryBirdLarge(53, 117) <= 4; angryBirdLarge(53, 118) <= 4; angryBirdLarge(53, 119) <= 4; angryBirdLarge(53, 120) <= 4; angryBirdLarge(53, 121) <= 4; angryBirdLarge(53, 122) <= 4; angryBirdLarge(53, 123) <= 4; angryBirdLarge(53, 124) <= 4; angryBirdLarge(53, 125) <= 4; angryBirdLarge(53, 126) <= 4; angryBirdLarge(53, 127) <= 4; angryBirdLarge(53, 128) <= 4; angryBirdLarge(53, 129) <= 4; angryBirdLarge(53, 130) <= 4; angryBirdLarge(53, 131) <= 4; angryBirdLarge(53, 132) <= 5; angryBirdLarge(53, 133) <= 5; angryBirdLarge(53, 134) <= 5; angryBirdLarge(53, 135) <= 5; angryBirdLarge(53, 136) <= 5; angryBirdLarge(53, 137) <= 5; angryBirdLarge(53, 138) <= 0; angryBirdLarge(53, 139) <= 0; angryBirdLarge(53, 140) <= 0; angryBirdLarge(53, 141) <= 0; angryBirdLarge(53, 142) <= 0; angryBirdLarge(53, 143) <= 0; angryBirdLarge(53, 144) <= 0; angryBirdLarge(53, 145) <= 0; angryBirdLarge(53, 146) <= 0; angryBirdLarge(53, 147) <= 0; angryBirdLarge(53, 148) <= 0; angryBirdLarge(53, 149) <= 0; 
angryBirdLarge(54, 0) <= 0; angryBirdLarge(54, 1) <= 0; angryBirdLarge(54, 2) <= 0; angryBirdLarge(54, 3) <= 0; angryBirdLarge(54, 4) <= 0; angryBirdLarge(54, 5) <= 0; angryBirdLarge(54, 6) <= 0; angryBirdLarge(54, 7) <= 0; angryBirdLarge(54, 8) <= 0; angryBirdLarge(54, 9) <= 0; angryBirdLarge(54, 10) <= 0; angryBirdLarge(54, 11) <= 0; angryBirdLarge(54, 12) <= 0; angryBirdLarge(54, 13) <= 0; angryBirdLarge(54, 14) <= 0; angryBirdLarge(54, 15) <= 0; angryBirdLarge(54, 16) <= 0; angryBirdLarge(54, 17) <= 0; angryBirdLarge(54, 18) <= 0; angryBirdLarge(54, 19) <= 0; angryBirdLarge(54, 20) <= 0; angryBirdLarge(54, 21) <= 0; angryBirdLarge(54, 22) <= 0; angryBirdLarge(54, 23) <= 0; angryBirdLarge(54, 24) <= 0; angryBirdLarge(54, 25) <= 0; angryBirdLarge(54, 26) <= 0; angryBirdLarge(54, 27) <= 0; angryBirdLarge(54, 28) <= 0; angryBirdLarge(54, 29) <= 0; angryBirdLarge(54, 30) <= 0; angryBirdLarge(54, 31) <= 0; angryBirdLarge(54, 32) <= 0; angryBirdLarge(54, 33) <= 0; angryBirdLarge(54, 34) <= 0; angryBirdLarge(54, 35) <= 0; angryBirdLarge(54, 36) <= 5; angryBirdLarge(54, 37) <= 5; angryBirdLarge(54, 38) <= 5; angryBirdLarge(54, 39) <= 5; angryBirdLarge(54, 40) <= 5; angryBirdLarge(54, 41) <= 5; angryBirdLarge(54, 42) <= 4; angryBirdLarge(54, 43) <= 4; angryBirdLarge(54, 44) <= 4; angryBirdLarge(54, 45) <= 4; angryBirdLarge(54, 46) <= 4; angryBirdLarge(54, 47) <= 4; angryBirdLarge(54, 48) <= 4; angryBirdLarge(54, 49) <= 4; angryBirdLarge(54, 50) <= 4; angryBirdLarge(54, 51) <= 4; angryBirdLarge(54, 52) <= 4; angryBirdLarge(54, 53) <= 4; angryBirdLarge(54, 54) <= 4; angryBirdLarge(54, 55) <= 4; angryBirdLarge(54, 56) <= 4; angryBirdLarge(54, 57) <= 4; angryBirdLarge(54, 58) <= 4; angryBirdLarge(54, 59) <= 4; angryBirdLarge(54, 60) <= 4; angryBirdLarge(54, 61) <= 4; angryBirdLarge(54, 62) <= 4; angryBirdLarge(54, 63) <= 4; angryBirdLarge(54, 64) <= 4; angryBirdLarge(54, 65) <= 4; angryBirdLarge(54, 66) <= 4; angryBirdLarge(54, 67) <= 4; angryBirdLarge(54, 68) <= 4; angryBirdLarge(54, 69) <= 4; angryBirdLarge(54, 70) <= 4; angryBirdLarge(54, 71) <= 4; angryBirdLarge(54, 72) <= 4; angryBirdLarge(54, 73) <= 4; angryBirdLarge(54, 74) <= 4; angryBirdLarge(54, 75) <= 4; angryBirdLarge(54, 76) <= 4; angryBirdLarge(54, 77) <= 4; angryBirdLarge(54, 78) <= 4; angryBirdLarge(54, 79) <= 4; angryBirdLarge(54, 80) <= 4; angryBirdLarge(54, 81) <= 4; angryBirdLarge(54, 82) <= 4; angryBirdLarge(54, 83) <= 4; angryBirdLarge(54, 84) <= 4; angryBirdLarge(54, 85) <= 4; angryBirdLarge(54, 86) <= 4; angryBirdLarge(54, 87) <= 4; angryBirdLarge(54, 88) <= 4; angryBirdLarge(54, 89) <= 4; angryBirdLarge(54, 90) <= 4; angryBirdLarge(54, 91) <= 4; angryBirdLarge(54, 92) <= 4; angryBirdLarge(54, 93) <= 4; angryBirdLarge(54, 94) <= 4; angryBirdLarge(54, 95) <= 4; angryBirdLarge(54, 96) <= 4; angryBirdLarge(54, 97) <= 4; angryBirdLarge(54, 98) <= 4; angryBirdLarge(54, 99) <= 4; angryBirdLarge(54, 100) <= 4; angryBirdLarge(54, 101) <= 4; angryBirdLarge(54, 102) <= 4; angryBirdLarge(54, 103) <= 4; angryBirdLarge(54, 104) <= 4; angryBirdLarge(54, 105) <= 4; angryBirdLarge(54, 106) <= 4; angryBirdLarge(54, 107) <= 4; angryBirdLarge(54, 108) <= 4; angryBirdLarge(54, 109) <= 4; angryBirdLarge(54, 110) <= 4; angryBirdLarge(54, 111) <= 4; angryBirdLarge(54, 112) <= 4; angryBirdLarge(54, 113) <= 4; angryBirdLarge(54, 114) <= 4; angryBirdLarge(54, 115) <= 4; angryBirdLarge(54, 116) <= 4; angryBirdLarge(54, 117) <= 4; angryBirdLarge(54, 118) <= 4; angryBirdLarge(54, 119) <= 4; angryBirdLarge(54, 120) <= 4; angryBirdLarge(54, 121) <= 4; angryBirdLarge(54, 122) <= 4; angryBirdLarge(54, 123) <= 4; angryBirdLarge(54, 124) <= 4; angryBirdLarge(54, 125) <= 4; angryBirdLarge(54, 126) <= 4; angryBirdLarge(54, 127) <= 4; angryBirdLarge(54, 128) <= 4; angryBirdLarge(54, 129) <= 4; angryBirdLarge(54, 130) <= 4; angryBirdLarge(54, 131) <= 4; angryBirdLarge(54, 132) <= 4; angryBirdLarge(54, 133) <= 4; angryBirdLarge(54, 134) <= 4; angryBirdLarge(54, 135) <= 4; angryBirdLarge(54, 136) <= 4; angryBirdLarge(54, 137) <= 4; angryBirdLarge(54, 138) <= 5; angryBirdLarge(54, 139) <= 5; angryBirdLarge(54, 140) <= 5; angryBirdLarge(54, 141) <= 5; angryBirdLarge(54, 142) <= 5; angryBirdLarge(54, 143) <= 5; angryBirdLarge(54, 144) <= 0; angryBirdLarge(54, 145) <= 0; angryBirdLarge(54, 146) <= 0; angryBirdLarge(54, 147) <= 0; angryBirdLarge(54, 148) <= 0; angryBirdLarge(54, 149) <= 0; 
angryBirdLarge(55, 0) <= 0; angryBirdLarge(55, 1) <= 0; angryBirdLarge(55, 2) <= 0; angryBirdLarge(55, 3) <= 0; angryBirdLarge(55, 4) <= 0; angryBirdLarge(55, 5) <= 0; angryBirdLarge(55, 6) <= 0; angryBirdLarge(55, 7) <= 0; angryBirdLarge(55, 8) <= 0; angryBirdLarge(55, 9) <= 0; angryBirdLarge(55, 10) <= 0; angryBirdLarge(55, 11) <= 0; angryBirdLarge(55, 12) <= 0; angryBirdLarge(55, 13) <= 0; angryBirdLarge(55, 14) <= 0; angryBirdLarge(55, 15) <= 0; angryBirdLarge(55, 16) <= 0; angryBirdLarge(55, 17) <= 0; angryBirdLarge(55, 18) <= 0; angryBirdLarge(55, 19) <= 0; angryBirdLarge(55, 20) <= 0; angryBirdLarge(55, 21) <= 0; angryBirdLarge(55, 22) <= 0; angryBirdLarge(55, 23) <= 0; angryBirdLarge(55, 24) <= 0; angryBirdLarge(55, 25) <= 0; angryBirdLarge(55, 26) <= 0; angryBirdLarge(55, 27) <= 0; angryBirdLarge(55, 28) <= 0; angryBirdLarge(55, 29) <= 0; angryBirdLarge(55, 30) <= 0; angryBirdLarge(55, 31) <= 0; angryBirdLarge(55, 32) <= 0; angryBirdLarge(55, 33) <= 0; angryBirdLarge(55, 34) <= 0; angryBirdLarge(55, 35) <= 0; angryBirdLarge(55, 36) <= 5; angryBirdLarge(55, 37) <= 5; angryBirdLarge(55, 38) <= 5; angryBirdLarge(55, 39) <= 5; angryBirdLarge(55, 40) <= 5; angryBirdLarge(55, 41) <= 5; angryBirdLarge(55, 42) <= 4; angryBirdLarge(55, 43) <= 4; angryBirdLarge(55, 44) <= 4; angryBirdLarge(55, 45) <= 4; angryBirdLarge(55, 46) <= 4; angryBirdLarge(55, 47) <= 4; angryBirdLarge(55, 48) <= 4; angryBirdLarge(55, 49) <= 4; angryBirdLarge(55, 50) <= 4; angryBirdLarge(55, 51) <= 4; angryBirdLarge(55, 52) <= 4; angryBirdLarge(55, 53) <= 4; angryBirdLarge(55, 54) <= 4; angryBirdLarge(55, 55) <= 4; angryBirdLarge(55, 56) <= 4; angryBirdLarge(55, 57) <= 4; angryBirdLarge(55, 58) <= 4; angryBirdLarge(55, 59) <= 4; angryBirdLarge(55, 60) <= 4; angryBirdLarge(55, 61) <= 4; angryBirdLarge(55, 62) <= 4; angryBirdLarge(55, 63) <= 4; angryBirdLarge(55, 64) <= 4; angryBirdLarge(55, 65) <= 4; angryBirdLarge(55, 66) <= 4; angryBirdLarge(55, 67) <= 4; angryBirdLarge(55, 68) <= 4; angryBirdLarge(55, 69) <= 4; angryBirdLarge(55, 70) <= 4; angryBirdLarge(55, 71) <= 4; angryBirdLarge(55, 72) <= 4; angryBirdLarge(55, 73) <= 4; angryBirdLarge(55, 74) <= 4; angryBirdLarge(55, 75) <= 4; angryBirdLarge(55, 76) <= 4; angryBirdLarge(55, 77) <= 4; angryBirdLarge(55, 78) <= 4; angryBirdLarge(55, 79) <= 4; angryBirdLarge(55, 80) <= 4; angryBirdLarge(55, 81) <= 4; angryBirdLarge(55, 82) <= 4; angryBirdLarge(55, 83) <= 4; angryBirdLarge(55, 84) <= 4; angryBirdLarge(55, 85) <= 4; angryBirdLarge(55, 86) <= 4; angryBirdLarge(55, 87) <= 4; angryBirdLarge(55, 88) <= 4; angryBirdLarge(55, 89) <= 4; angryBirdLarge(55, 90) <= 4; angryBirdLarge(55, 91) <= 4; angryBirdLarge(55, 92) <= 4; angryBirdLarge(55, 93) <= 4; angryBirdLarge(55, 94) <= 4; angryBirdLarge(55, 95) <= 4; angryBirdLarge(55, 96) <= 4; angryBirdLarge(55, 97) <= 4; angryBirdLarge(55, 98) <= 4; angryBirdLarge(55, 99) <= 4; angryBirdLarge(55, 100) <= 4; angryBirdLarge(55, 101) <= 4; angryBirdLarge(55, 102) <= 4; angryBirdLarge(55, 103) <= 4; angryBirdLarge(55, 104) <= 4; angryBirdLarge(55, 105) <= 4; angryBirdLarge(55, 106) <= 4; angryBirdLarge(55, 107) <= 4; angryBirdLarge(55, 108) <= 4; angryBirdLarge(55, 109) <= 4; angryBirdLarge(55, 110) <= 4; angryBirdLarge(55, 111) <= 4; angryBirdLarge(55, 112) <= 4; angryBirdLarge(55, 113) <= 4; angryBirdLarge(55, 114) <= 4; angryBirdLarge(55, 115) <= 4; angryBirdLarge(55, 116) <= 4; angryBirdLarge(55, 117) <= 4; angryBirdLarge(55, 118) <= 4; angryBirdLarge(55, 119) <= 4; angryBirdLarge(55, 120) <= 4; angryBirdLarge(55, 121) <= 4; angryBirdLarge(55, 122) <= 4; angryBirdLarge(55, 123) <= 4; angryBirdLarge(55, 124) <= 4; angryBirdLarge(55, 125) <= 4; angryBirdLarge(55, 126) <= 4; angryBirdLarge(55, 127) <= 4; angryBirdLarge(55, 128) <= 4; angryBirdLarge(55, 129) <= 4; angryBirdLarge(55, 130) <= 4; angryBirdLarge(55, 131) <= 4; angryBirdLarge(55, 132) <= 4; angryBirdLarge(55, 133) <= 4; angryBirdLarge(55, 134) <= 4; angryBirdLarge(55, 135) <= 4; angryBirdLarge(55, 136) <= 4; angryBirdLarge(55, 137) <= 4; angryBirdLarge(55, 138) <= 5; angryBirdLarge(55, 139) <= 5; angryBirdLarge(55, 140) <= 5; angryBirdLarge(55, 141) <= 5; angryBirdLarge(55, 142) <= 5; angryBirdLarge(55, 143) <= 5; angryBirdLarge(55, 144) <= 0; angryBirdLarge(55, 145) <= 0; angryBirdLarge(55, 146) <= 0; angryBirdLarge(55, 147) <= 0; angryBirdLarge(55, 148) <= 0; angryBirdLarge(55, 149) <= 0; 
angryBirdLarge(56, 0) <= 0; angryBirdLarge(56, 1) <= 0; angryBirdLarge(56, 2) <= 0; angryBirdLarge(56, 3) <= 0; angryBirdLarge(56, 4) <= 0; angryBirdLarge(56, 5) <= 0; angryBirdLarge(56, 6) <= 0; angryBirdLarge(56, 7) <= 0; angryBirdLarge(56, 8) <= 0; angryBirdLarge(56, 9) <= 0; angryBirdLarge(56, 10) <= 0; angryBirdLarge(56, 11) <= 0; angryBirdLarge(56, 12) <= 0; angryBirdLarge(56, 13) <= 0; angryBirdLarge(56, 14) <= 0; angryBirdLarge(56, 15) <= 0; angryBirdLarge(56, 16) <= 0; angryBirdLarge(56, 17) <= 0; angryBirdLarge(56, 18) <= 0; angryBirdLarge(56, 19) <= 0; angryBirdLarge(56, 20) <= 0; angryBirdLarge(56, 21) <= 0; angryBirdLarge(56, 22) <= 0; angryBirdLarge(56, 23) <= 0; angryBirdLarge(56, 24) <= 0; angryBirdLarge(56, 25) <= 0; angryBirdLarge(56, 26) <= 0; angryBirdLarge(56, 27) <= 0; angryBirdLarge(56, 28) <= 0; angryBirdLarge(56, 29) <= 0; angryBirdLarge(56, 30) <= 0; angryBirdLarge(56, 31) <= 0; angryBirdLarge(56, 32) <= 0; angryBirdLarge(56, 33) <= 0; angryBirdLarge(56, 34) <= 0; angryBirdLarge(56, 35) <= 0; angryBirdLarge(56, 36) <= 5; angryBirdLarge(56, 37) <= 5; angryBirdLarge(56, 38) <= 5; angryBirdLarge(56, 39) <= 5; angryBirdLarge(56, 40) <= 5; angryBirdLarge(56, 41) <= 5; angryBirdLarge(56, 42) <= 4; angryBirdLarge(56, 43) <= 4; angryBirdLarge(56, 44) <= 4; angryBirdLarge(56, 45) <= 4; angryBirdLarge(56, 46) <= 4; angryBirdLarge(56, 47) <= 4; angryBirdLarge(56, 48) <= 4; angryBirdLarge(56, 49) <= 4; angryBirdLarge(56, 50) <= 4; angryBirdLarge(56, 51) <= 4; angryBirdLarge(56, 52) <= 4; angryBirdLarge(56, 53) <= 4; angryBirdLarge(56, 54) <= 4; angryBirdLarge(56, 55) <= 4; angryBirdLarge(56, 56) <= 4; angryBirdLarge(56, 57) <= 4; angryBirdLarge(56, 58) <= 4; angryBirdLarge(56, 59) <= 4; angryBirdLarge(56, 60) <= 4; angryBirdLarge(56, 61) <= 4; angryBirdLarge(56, 62) <= 4; angryBirdLarge(56, 63) <= 4; angryBirdLarge(56, 64) <= 4; angryBirdLarge(56, 65) <= 4; angryBirdLarge(56, 66) <= 4; angryBirdLarge(56, 67) <= 4; angryBirdLarge(56, 68) <= 4; angryBirdLarge(56, 69) <= 4; angryBirdLarge(56, 70) <= 4; angryBirdLarge(56, 71) <= 4; angryBirdLarge(56, 72) <= 4; angryBirdLarge(56, 73) <= 4; angryBirdLarge(56, 74) <= 4; angryBirdLarge(56, 75) <= 4; angryBirdLarge(56, 76) <= 4; angryBirdLarge(56, 77) <= 4; angryBirdLarge(56, 78) <= 4; angryBirdLarge(56, 79) <= 4; angryBirdLarge(56, 80) <= 4; angryBirdLarge(56, 81) <= 4; angryBirdLarge(56, 82) <= 4; angryBirdLarge(56, 83) <= 4; angryBirdLarge(56, 84) <= 4; angryBirdLarge(56, 85) <= 4; angryBirdLarge(56, 86) <= 4; angryBirdLarge(56, 87) <= 4; angryBirdLarge(56, 88) <= 4; angryBirdLarge(56, 89) <= 4; angryBirdLarge(56, 90) <= 4; angryBirdLarge(56, 91) <= 4; angryBirdLarge(56, 92) <= 4; angryBirdLarge(56, 93) <= 4; angryBirdLarge(56, 94) <= 4; angryBirdLarge(56, 95) <= 4; angryBirdLarge(56, 96) <= 4; angryBirdLarge(56, 97) <= 4; angryBirdLarge(56, 98) <= 4; angryBirdLarge(56, 99) <= 4; angryBirdLarge(56, 100) <= 4; angryBirdLarge(56, 101) <= 4; angryBirdLarge(56, 102) <= 4; angryBirdLarge(56, 103) <= 4; angryBirdLarge(56, 104) <= 4; angryBirdLarge(56, 105) <= 4; angryBirdLarge(56, 106) <= 4; angryBirdLarge(56, 107) <= 4; angryBirdLarge(56, 108) <= 4; angryBirdLarge(56, 109) <= 4; angryBirdLarge(56, 110) <= 4; angryBirdLarge(56, 111) <= 4; angryBirdLarge(56, 112) <= 4; angryBirdLarge(56, 113) <= 4; angryBirdLarge(56, 114) <= 4; angryBirdLarge(56, 115) <= 4; angryBirdLarge(56, 116) <= 4; angryBirdLarge(56, 117) <= 4; angryBirdLarge(56, 118) <= 4; angryBirdLarge(56, 119) <= 4; angryBirdLarge(56, 120) <= 4; angryBirdLarge(56, 121) <= 4; angryBirdLarge(56, 122) <= 4; angryBirdLarge(56, 123) <= 4; angryBirdLarge(56, 124) <= 4; angryBirdLarge(56, 125) <= 4; angryBirdLarge(56, 126) <= 4; angryBirdLarge(56, 127) <= 4; angryBirdLarge(56, 128) <= 4; angryBirdLarge(56, 129) <= 4; angryBirdLarge(56, 130) <= 4; angryBirdLarge(56, 131) <= 4; angryBirdLarge(56, 132) <= 4; angryBirdLarge(56, 133) <= 4; angryBirdLarge(56, 134) <= 4; angryBirdLarge(56, 135) <= 4; angryBirdLarge(56, 136) <= 4; angryBirdLarge(56, 137) <= 4; angryBirdLarge(56, 138) <= 5; angryBirdLarge(56, 139) <= 5; angryBirdLarge(56, 140) <= 5; angryBirdLarge(56, 141) <= 5; angryBirdLarge(56, 142) <= 5; angryBirdLarge(56, 143) <= 5; angryBirdLarge(56, 144) <= 0; angryBirdLarge(56, 145) <= 0; angryBirdLarge(56, 146) <= 0; angryBirdLarge(56, 147) <= 0; angryBirdLarge(56, 148) <= 0; angryBirdLarge(56, 149) <= 0; 
angryBirdLarge(57, 0) <= 0; angryBirdLarge(57, 1) <= 0; angryBirdLarge(57, 2) <= 0; angryBirdLarge(57, 3) <= 0; angryBirdLarge(57, 4) <= 0; angryBirdLarge(57, 5) <= 0; angryBirdLarge(57, 6) <= 0; angryBirdLarge(57, 7) <= 0; angryBirdLarge(57, 8) <= 0; angryBirdLarge(57, 9) <= 0; angryBirdLarge(57, 10) <= 0; angryBirdLarge(57, 11) <= 0; angryBirdLarge(57, 12) <= 0; angryBirdLarge(57, 13) <= 0; angryBirdLarge(57, 14) <= 0; angryBirdLarge(57, 15) <= 0; angryBirdLarge(57, 16) <= 0; angryBirdLarge(57, 17) <= 0; angryBirdLarge(57, 18) <= 0; angryBirdLarge(57, 19) <= 0; angryBirdLarge(57, 20) <= 0; angryBirdLarge(57, 21) <= 0; angryBirdLarge(57, 22) <= 0; angryBirdLarge(57, 23) <= 0; angryBirdLarge(57, 24) <= 0; angryBirdLarge(57, 25) <= 0; angryBirdLarge(57, 26) <= 0; angryBirdLarge(57, 27) <= 0; angryBirdLarge(57, 28) <= 0; angryBirdLarge(57, 29) <= 0; angryBirdLarge(57, 30) <= 0; angryBirdLarge(57, 31) <= 0; angryBirdLarge(57, 32) <= 0; angryBirdLarge(57, 33) <= 0; angryBirdLarge(57, 34) <= 0; angryBirdLarge(57, 35) <= 0; angryBirdLarge(57, 36) <= 5; angryBirdLarge(57, 37) <= 5; angryBirdLarge(57, 38) <= 5; angryBirdLarge(57, 39) <= 5; angryBirdLarge(57, 40) <= 5; angryBirdLarge(57, 41) <= 5; angryBirdLarge(57, 42) <= 4; angryBirdLarge(57, 43) <= 4; angryBirdLarge(57, 44) <= 4; angryBirdLarge(57, 45) <= 4; angryBirdLarge(57, 46) <= 4; angryBirdLarge(57, 47) <= 4; angryBirdLarge(57, 48) <= 4; angryBirdLarge(57, 49) <= 4; angryBirdLarge(57, 50) <= 4; angryBirdLarge(57, 51) <= 4; angryBirdLarge(57, 52) <= 4; angryBirdLarge(57, 53) <= 4; angryBirdLarge(57, 54) <= 4; angryBirdLarge(57, 55) <= 4; angryBirdLarge(57, 56) <= 4; angryBirdLarge(57, 57) <= 4; angryBirdLarge(57, 58) <= 4; angryBirdLarge(57, 59) <= 4; angryBirdLarge(57, 60) <= 4; angryBirdLarge(57, 61) <= 4; angryBirdLarge(57, 62) <= 4; angryBirdLarge(57, 63) <= 4; angryBirdLarge(57, 64) <= 4; angryBirdLarge(57, 65) <= 4; angryBirdLarge(57, 66) <= 4; angryBirdLarge(57, 67) <= 4; angryBirdLarge(57, 68) <= 4; angryBirdLarge(57, 69) <= 4; angryBirdLarge(57, 70) <= 4; angryBirdLarge(57, 71) <= 4; angryBirdLarge(57, 72) <= 4; angryBirdLarge(57, 73) <= 4; angryBirdLarge(57, 74) <= 4; angryBirdLarge(57, 75) <= 4; angryBirdLarge(57, 76) <= 4; angryBirdLarge(57, 77) <= 4; angryBirdLarge(57, 78) <= 4; angryBirdLarge(57, 79) <= 4; angryBirdLarge(57, 80) <= 4; angryBirdLarge(57, 81) <= 4; angryBirdLarge(57, 82) <= 4; angryBirdLarge(57, 83) <= 4; angryBirdLarge(57, 84) <= 4; angryBirdLarge(57, 85) <= 4; angryBirdLarge(57, 86) <= 4; angryBirdLarge(57, 87) <= 4; angryBirdLarge(57, 88) <= 4; angryBirdLarge(57, 89) <= 4; angryBirdLarge(57, 90) <= 4; angryBirdLarge(57, 91) <= 4; angryBirdLarge(57, 92) <= 4; angryBirdLarge(57, 93) <= 4; angryBirdLarge(57, 94) <= 4; angryBirdLarge(57, 95) <= 4; angryBirdLarge(57, 96) <= 4; angryBirdLarge(57, 97) <= 4; angryBirdLarge(57, 98) <= 4; angryBirdLarge(57, 99) <= 4; angryBirdLarge(57, 100) <= 4; angryBirdLarge(57, 101) <= 4; angryBirdLarge(57, 102) <= 4; angryBirdLarge(57, 103) <= 4; angryBirdLarge(57, 104) <= 4; angryBirdLarge(57, 105) <= 4; angryBirdLarge(57, 106) <= 4; angryBirdLarge(57, 107) <= 4; angryBirdLarge(57, 108) <= 4; angryBirdLarge(57, 109) <= 4; angryBirdLarge(57, 110) <= 4; angryBirdLarge(57, 111) <= 4; angryBirdLarge(57, 112) <= 4; angryBirdLarge(57, 113) <= 4; angryBirdLarge(57, 114) <= 4; angryBirdLarge(57, 115) <= 4; angryBirdLarge(57, 116) <= 4; angryBirdLarge(57, 117) <= 4; angryBirdLarge(57, 118) <= 4; angryBirdLarge(57, 119) <= 4; angryBirdLarge(57, 120) <= 4; angryBirdLarge(57, 121) <= 4; angryBirdLarge(57, 122) <= 4; angryBirdLarge(57, 123) <= 4; angryBirdLarge(57, 124) <= 4; angryBirdLarge(57, 125) <= 4; angryBirdLarge(57, 126) <= 4; angryBirdLarge(57, 127) <= 4; angryBirdLarge(57, 128) <= 4; angryBirdLarge(57, 129) <= 4; angryBirdLarge(57, 130) <= 4; angryBirdLarge(57, 131) <= 4; angryBirdLarge(57, 132) <= 4; angryBirdLarge(57, 133) <= 4; angryBirdLarge(57, 134) <= 4; angryBirdLarge(57, 135) <= 4; angryBirdLarge(57, 136) <= 4; angryBirdLarge(57, 137) <= 4; angryBirdLarge(57, 138) <= 5; angryBirdLarge(57, 139) <= 5; angryBirdLarge(57, 140) <= 5; angryBirdLarge(57, 141) <= 5; angryBirdLarge(57, 142) <= 5; angryBirdLarge(57, 143) <= 5; angryBirdLarge(57, 144) <= 0; angryBirdLarge(57, 145) <= 0; angryBirdLarge(57, 146) <= 0; angryBirdLarge(57, 147) <= 0; angryBirdLarge(57, 148) <= 0; angryBirdLarge(57, 149) <= 0; 
angryBirdLarge(58, 0) <= 0; angryBirdLarge(58, 1) <= 0; angryBirdLarge(58, 2) <= 0; angryBirdLarge(58, 3) <= 0; angryBirdLarge(58, 4) <= 0; angryBirdLarge(58, 5) <= 0; angryBirdLarge(58, 6) <= 0; angryBirdLarge(58, 7) <= 0; angryBirdLarge(58, 8) <= 0; angryBirdLarge(58, 9) <= 0; angryBirdLarge(58, 10) <= 0; angryBirdLarge(58, 11) <= 0; angryBirdLarge(58, 12) <= 0; angryBirdLarge(58, 13) <= 0; angryBirdLarge(58, 14) <= 0; angryBirdLarge(58, 15) <= 0; angryBirdLarge(58, 16) <= 0; angryBirdLarge(58, 17) <= 0; angryBirdLarge(58, 18) <= 0; angryBirdLarge(58, 19) <= 0; angryBirdLarge(58, 20) <= 0; angryBirdLarge(58, 21) <= 0; angryBirdLarge(58, 22) <= 0; angryBirdLarge(58, 23) <= 0; angryBirdLarge(58, 24) <= 0; angryBirdLarge(58, 25) <= 0; angryBirdLarge(58, 26) <= 0; angryBirdLarge(58, 27) <= 0; angryBirdLarge(58, 28) <= 0; angryBirdLarge(58, 29) <= 0; angryBirdLarge(58, 30) <= 0; angryBirdLarge(58, 31) <= 0; angryBirdLarge(58, 32) <= 0; angryBirdLarge(58, 33) <= 0; angryBirdLarge(58, 34) <= 0; angryBirdLarge(58, 35) <= 0; angryBirdLarge(58, 36) <= 5; angryBirdLarge(58, 37) <= 5; angryBirdLarge(58, 38) <= 5; angryBirdLarge(58, 39) <= 5; angryBirdLarge(58, 40) <= 5; angryBirdLarge(58, 41) <= 5; angryBirdLarge(58, 42) <= 4; angryBirdLarge(58, 43) <= 4; angryBirdLarge(58, 44) <= 4; angryBirdLarge(58, 45) <= 4; angryBirdLarge(58, 46) <= 4; angryBirdLarge(58, 47) <= 4; angryBirdLarge(58, 48) <= 4; angryBirdLarge(58, 49) <= 4; angryBirdLarge(58, 50) <= 4; angryBirdLarge(58, 51) <= 4; angryBirdLarge(58, 52) <= 4; angryBirdLarge(58, 53) <= 4; angryBirdLarge(58, 54) <= 4; angryBirdLarge(58, 55) <= 4; angryBirdLarge(58, 56) <= 4; angryBirdLarge(58, 57) <= 4; angryBirdLarge(58, 58) <= 4; angryBirdLarge(58, 59) <= 4; angryBirdLarge(58, 60) <= 4; angryBirdLarge(58, 61) <= 4; angryBirdLarge(58, 62) <= 4; angryBirdLarge(58, 63) <= 4; angryBirdLarge(58, 64) <= 4; angryBirdLarge(58, 65) <= 4; angryBirdLarge(58, 66) <= 4; angryBirdLarge(58, 67) <= 4; angryBirdLarge(58, 68) <= 4; angryBirdLarge(58, 69) <= 4; angryBirdLarge(58, 70) <= 4; angryBirdLarge(58, 71) <= 4; angryBirdLarge(58, 72) <= 4; angryBirdLarge(58, 73) <= 4; angryBirdLarge(58, 74) <= 4; angryBirdLarge(58, 75) <= 4; angryBirdLarge(58, 76) <= 4; angryBirdLarge(58, 77) <= 4; angryBirdLarge(58, 78) <= 4; angryBirdLarge(58, 79) <= 4; angryBirdLarge(58, 80) <= 4; angryBirdLarge(58, 81) <= 4; angryBirdLarge(58, 82) <= 4; angryBirdLarge(58, 83) <= 4; angryBirdLarge(58, 84) <= 4; angryBirdLarge(58, 85) <= 4; angryBirdLarge(58, 86) <= 4; angryBirdLarge(58, 87) <= 4; angryBirdLarge(58, 88) <= 4; angryBirdLarge(58, 89) <= 4; angryBirdLarge(58, 90) <= 4; angryBirdLarge(58, 91) <= 4; angryBirdLarge(58, 92) <= 4; angryBirdLarge(58, 93) <= 4; angryBirdLarge(58, 94) <= 4; angryBirdLarge(58, 95) <= 4; angryBirdLarge(58, 96) <= 4; angryBirdLarge(58, 97) <= 4; angryBirdLarge(58, 98) <= 4; angryBirdLarge(58, 99) <= 4; angryBirdLarge(58, 100) <= 4; angryBirdLarge(58, 101) <= 4; angryBirdLarge(58, 102) <= 4; angryBirdLarge(58, 103) <= 4; angryBirdLarge(58, 104) <= 4; angryBirdLarge(58, 105) <= 4; angryBirdLarge(58, 106) <= 4; angryBirdLarge(58, 107) <= 4; angryBirdLarge(58, 108) <= 4; angryBirdLarge(58, 109) <= 4; angryBirdLarge(58, 110) <= 4; angryBirdLarge(58, 111) <= 4; angryBirdLarge(58, 112) <= 4; angryBirdLarge(58, 113) <= 4; angryBirdLarge(58, 114) <= 4; angryBirdLarge(58, 115) <= 4; angryBirdLarge(58, 116) <= 4; angryBirdLarge(58, 117) <= 4; angryBirdLarge(58, 118) <= 4; angryBirdLarge(58, 119) <= 4; angryBirdLarge(58, 120) <= 4; angryBirdLarge(58, 121) <= 4; angryBirdLarge(58, 122) <= 4; angryBirdLarge(58, 123) <= 4; angryBirdLarge(58, 124) <= 4; angryBirdLarge(58, 125) <= 4; angryBirdLarge(58, 126) <= 4; angryBirdLarge(58, 127) <= 4; angryBirdLarge(58, 128) <= 4; angryBirdLarge(58, 129) <= 4; angryBirdLarge(58, 130) <= 4; angryBirdLarge(58, 131) <= 4; angryBirdLarge(58, 132) <= 4; angryBirdLarge(58, 133) <= 4; angryBirdLarge(58, 134) <= 4; angryBirdLarge(58, 135) <= 4; angryBirdLarge(58, 136) <= 4; angryBirdLarge(58, 137) <= 4; angryBirdLarge(58, 138) <= 5; angryBirdLarge(58, 139) <= 5; angryBirdLarge(58, 140) <= 5; angryBirdLarge(58, 141) <= 5; angryBirdLarge(58, 142) <= 5; angryBirdLarge(58, 143) <= 5; angryBirdLarge(58, 144) <= 0; angryBirdLarge(58, 145) <= 0; angryBirdLarge(58, 146) <= 0; angryBirdLarge(58, 147) <= 0; angryBirdLarge(58, 148) <= 0; angryBirdLarge(58, 149) <= 0; 
angryBirdLarge(59, 0) <= 0; angryBirdLarge(59, 1) <= 0; angryBirdLarge(59, 2) <= 0; angryBirdLarge(59, 3) <= 0; angryBirdLarge(59, 4) <= 0; angryBirdLarge(59, 5) <= 0; angryBirdLarge(59, 6) <= 0; angryBirdLarge(59, 7) <= 0; angryBirdLarge(59, 8) <= 0; angryBirdLarge(59, 9) <= 0; angryBirdLarge(59, 10) <= 0; angryBirdLarge(59, 11) <= 0; angryBirdLarge(59, 12) <= 0; angryBirdLarge(59, 13) <= 0; angryBirdLarge(59, 14) <= 0; angryBirdLarge(59, 15) <= 0; angryBirdLarge(59, 16) <= 0; angryBirdLarge(59, 17) <= 0; angryBirdLarge(59, 18) <= 0; angryBirdLarge(59, 19) <= 0; angryBirdLarge(59, 20) <= 0; angryBirdLarge(59, 21) <= 0; angryBirdLarge(59, 22) <= 0; angryBirdLarge(59, 23) <= 0; angryBirdLarge(59, 24) <= 0; angryBirdLarge(59, 25) <= 0; angryBirdLarge(59, 26) <= 0; angryBirdLarge(59, 27) <= 0; angryBirdLarge(59, 28) <= 0; angryBirdLarge(59, 29) <= 0; angryBirdLarge(59, 30) <= 0; angryBirdLarge(59, 31) <= 0; angryBirdLarge(59, 32) <= 0; angryBirdLarge(59, 33) <= 0; angryBirdLarge(59, 34) <= 0; angryBirdLarge(59, 35) <= 0; angryBirdLarge(59, 36) <= 5; angryBirdLarge(59, 37) <= 5; angryBirdLarge(59, 38) <= 5; angryBirdLarge(59, 39) <= 5; angryBirdLarge(59, 40) <= 5; angryBirdLarge(59, 41) <= 5; angryBirdLarge(59, 42) <= 4; angryBirdLarge(59, 43) <= 4; angryBirdLarge(59, 44) <= 4; angryBirdLarge(59, 45) <= 4; angryBirdLarge(59, 46) <= 4; angryBirdLarge(59, 47) <= 4; angryBirdLarge(59, 48) <= 4; angryBirdLarge(59, 49) <= 4; angryBirdLarge(59, 50) <= 4; angryBirdLarge(59, 51) <= 4; angryBirdLarge(59, 52) <= 4; angryBirdLarge(59, 53) <= 4; angryBirdLarge(59, 54) <= 4; angryBirdLarge(59, 55) <= 4; angryBirdLarge(59, 56) <= 4; angryBirdLarge(59, 57) <= 4; angryBirdLarge(59, 58) <= 4; angryBirdLarge(59, 59) <= 4; angryBirdLarge(59, 60) <= 4; angryBirdLarge(59, 61) <= 4; angryBirdLarge(59, 62) <= 4; angryBirdLarge(59, 63) <= 4; angryBirdLarge(59, 64) <= 4; angryBirdLarge(59, 65) <= 4; angryBirdLarge(59, 66) <= 4; angryBirdLarge(59, 67) <= 4; angryBirdLarge(59, 68) <= 4; angryBirdLarge(59, 69) <= 4; angryBirdLarge(59, 70) <= 4; angryBirdLarge(59, 71) <= 4; angryBirdLarge(59, 72) <= 4; angryBirdLarge(59, 73) <= 4; angryBirdLarge(59, 74) <= 4; angryBirdLarge(59, 75) <= 4; angryBirdLarge(59, 76) <= 4; angryBirdLarge(59, 77) <= 4; angryBirdLarge(59, 78) <= 4; angryBirdLarge(59, 79) <= 4; angryBirdLarge(59, 80) <= 4; angryBirdLarge(59, 81) <= 4; angryBirdLarge(59, 82) <= 4; angryBirdLarge(59, 83) <= 4; angryBirdLarge(59, 84) <= 4; angryBirdLarge(59, 85) <= 4; angryBirdLarge(59, 86) <= 4; angryBirdLarge(59, 87) <= 4; angryBirdLarge(59, 88) <= 4; angryBirdLarge(59, 89) <= 4; angryBirdLarge(59, 90) <= 4; angryBirdLarge(59, 91) <= 4; angryBirdLarge(59, 92) <= 4; angryBirdLarge(59, 93) <= 4; angryBirdLarge(59, 94) <= 4; angryBirdLarge(59, 95) <= 4; angryBirdLarge(59, 96) <= 4; angryBirdLarge(59, 97) <= 4; angryBirdLarge(59, 98) <= 4; angryBirdLarge(59, 99) <= 4; angryBirdLarge(59, 100) <= 4; angryBirdLarge(59, 101) <= 4; angryBirdLarge(59, 102) <= 4; angryBirdLarge(59, 103) <= 4; angryBirdLarge(59, 104) <= 4; angryBirdLarge(59, 105) <= 4; angryBirdLarge(59, 106) <= 4; angryBirdLarge(59, 107) <= 4; angryBirdLarge(59, 108) <= 4; angryBirdLarge(59, 109) <= 4; angryBirdLarge(59, 110) <= 4; angryBirdLarge(59, 111) <= 4; angryBirdLarge(59, 112) <= 4; angryBirdLarge(59, 113) <= 4; angryBirdLarge(59, 114) <= 4; angryBirdLarge(59, 115) <= 4; angryBirdLarge(59, 116) <= 4; angryBirdLarge(59, 117) <= 4; angryBirdLarge(59, 118) <= 4; angryBirdLarge(59, 119) <= 4; angryBirdLarge(59, 120) <= 4; angryBirdLarge(59, 121) <= 4; angryBirdLarge(59, 122) <= 4; angryBirdLarge(59, 123) <= 4; angryBirdLarge(59, 124) <= 4; angryBirdLarge(59, 125) <= 4; angryBirdLarge(59, 126) <= 4; angryBirdLarge(59, 127) <= 4; angryBirdLarge(59, 128) <= 4; angryBirdLarge(59, 129) <= 4; angryBirdLarge(59, 130) <= 4; angryBirdLarge(59, 131) <= 4; angryBirdLarge(59, 132) <= 4; angryBirdLarge(59, 133) <= 4; angryBirdLarge(59, 134) <= 4; angryBirdLarge(59, 135) <= 4; angryBirdLarge(59, 136) <= 4; angryBirdLarge(59, 137) <= 4; angryBirdLarge(59, 138) <= 5; angryBirdLarge(59, 139) <= 5; angryBirdLarge(59, 140) <= 5; angryBirdLarge(59, 141) <= 5; angryBirdLarge(59, 142) <= 5; angryBirdLarge(59, 143) <= 5; angryBirdLarge(59, 144) <= 0; angryBirdLarge(59, 145) <= 0; angryBirdLarge(59, 146) <= 0; angryBirdLarge(59, 147) <= 0; angryBirdLarge(59, 148) <= 0; angryBirdLarge(59, 149) <= 0; 
angryBirdLarge(60, 0) <= 0; angryBirdLarge(60, 1) <= 0; angryBirdLarge(60, 2) <= 0; angryBirdLarge(60, 3) <= 0; angryBirdLarge(60, 4) <= 0; angryBirdLarge(60, 5) <= 0; angryBirdLarge(60, 6) <= 0; angryBirdLarge(60, 7) <= 0; angryBirdLarge(60, 8) <= 0; angryBirdLarge(60, 9) <= 0; angryBirdLarge(60, 10) <= 0; angryBirdLarge(60, 11) <= 0; angryBirdLarge(60, 12) <= 0; angryBirdLarge(60, 13) <= 0; angryBirdLarge(60, 14) <= 0; angryBirdLarge(60, 15) <= 0; angryBirdLarge(60, 16) <= 0; angryBirdLarge(60, 17) <= 0; angryBirdLarge(60, 18) <= 0; angryBirdLarge(60, 19) <= 0; angryBirdLarge(60, 20) <= 0; angryBirdLarge(60, 21) <= 0; angryBirdLarge(60, 22) <= 0; angryBirdLarge(60, 23) <= 0; angryBirdLarge(60, 24) <= 0; angryBirdLarge(60, 25) <= 0; angryBirdLarge(60, 26) <= 0; angryBirdLarge(60, 27) <= 0; angryBirdLarge(60, 28) <= 0; angryBirdLarge(60, 29) <= 0; angryBirdLarge(60, 30) <= 5; angryBirdLarge(60, 31) <= 5; angryBirdLarge(60, 32) <= 5; angryBirdLarge(60, 33) <= 5; angryBirdLarge(60, 34) <= 5; angryBirdLarge(60, 35) <= 5; angryBirdLarge(60, 36) <= 4; angryBirdLarge(60, 37) <= 4; angryBirdLarge(60, 38) <= 4; angryBirdLarge(60, 39) <= 4; angryBirdLarge(60, 40) <= 4; angryBirdLarge(60, 41) <= 4; angryBirdLarge(60, 42) <= 4; angryBirdLarge(60, 43) <= 4; angryBirdLarge(60, 44) <= 4; angryBirdLarge(60, 45) <= 4; angryBirdLarge(60, 46) <= 4; angryBirdLarge(60, 47) <= 4; angryBirdLarge(60, 48) <= 4; angryBirdLarge(60, 49) <= 4; angryBirdLarge(60, 50) <= 4; angryBirdLarge(60, 51) <= 4; angryBirdLarge(60, 52) <= 4; angryBirdLarge(60, 53) <= 4; angryBirdLarge(60, 54) <= 4; angryBirdLarge(60, 55) <= 4; angryBirdLarge(60, 56) <= 4; angryBirdLarge(60, 57) <= 4; angryBirdLarge(60, 58) <= 4; angryBirdLarge(60, 59) <= 4; angryBirdLarge(60, 60) <= 4; angryBirdLarge(60, 61) <= 4; angryBirdLarge(60, 62) <= 4; angryBirdLarge(60, 63) <= 4; angryBirdLarge(60, 64) <= 4; angryBirdLarge(60, 65) <= 4; angryBirdLarge(60, 66) <= 4; angryBirdLarge(60, 67) <= 4; angryBirdLarge(60, 68) <= 4; angryBirdLarge(60, 69) <= 4; angryBirdLarge(60, 70) <= 4; angryBirdLarge(60, 71) <= 4; angryBirdLarge(60, 72) <= 5; angryBirdLarge(60, 73) <= 5; angryBirdLarge(60, 74) <= 5; angryBirdLarge(60, 75) <= 5; angryBirdLarge(60, 76) <= 5; angryBirdLarge(60, 77) <= 5; angryBirdLarge(60, 78) <= 5; angryBirdLarge(60, 79) <= 5; angryBirdLarge(60, 80) <= 5; angryBirdLarge(60, 81) <= 5; angryBirdLarge(60, 82) <= 5; angryBirdLarge(60, 83) <= 5; angryBirdLarge(60, 84) <= 5; angryBirdLarge(60, 85) <= 5; angryBirdLarge(60, 86) <= 5; angryBirdLarge(60, 87) <= 5; angryBirdLarge(60, 88) <= 5; angryBirdLarge(60, 89) <= 5; angryBirdLarge(60, 90) <= 5; angryBirdLarge(60, 91) <= 5; angryBirdLarge(60, 92) <= 5; angryBirdLarge(60, 93) <= 5; angryBirdLarge(60, 94) <= 5; angryBirdLarge(60, 95) <= 5; angryBirdLarge(60, 96) <= 4; angryBirdLarge(60, 97) <= 4; angryBirdLarge(60, 98) <= 4; angryBirdLarge(60, 99) <= 4; angryBirdLarge(60, 100) <= 4; angryBirdLarge(60, 101) <= 4; angryBirdLarge(60, 102) <= 4; angryBirdLarge(60, 103) <= 4; angryBirdLarge(60, 104) <= 4; angryBirdLarge(60, 105) <= 4; angryBirdLarge(60, 106) <= 4; angryBirdLarge(60, 107) <= 4; angryBirdLarge(60, 108) <= 4; angryBirdLarge(60, 109) <= 4; angryBirdLarge(60, 110) <= 4; angryBirdLarge(60, 111) <= 4; angryBirdLarge(60, 112) <= 4; angryBirdLarge(60, 113) <= 4; angryBirdLarge(60, 114) <= 4; angryBirdLarge(60, 115) <= 4; angryBirdLarge(60, 116) <= 4; angryBirdLarge(60, 117) <= 4; angryBirdLarge(60, 118) <= 4; angryBirdLarge(60, 119) <= 4; angryBirdLarge(60, 120) <= 4; angryBirdLarge(60, 121) <= 4; angryBirdLarge(60, 122) <= 4; angryBirdLarge(60, 123) <= 4; angryBirdLarge(60, 124) <= 4; angryBirdLarge(60, 125) <= 4; angryBirdLarge(60, 126) <= 5; angryBirdLarge(60, 127) <= 5; angryBirdLarge(60, 128) <= 5; angryBirdLarge(60, 129) <= 5; angryBirdLarge(60, 130) <= 5; angryBirdLarge(60, 131) <= 5; angryBirdLarge(60, 132) <= 5; angryBirdLarge(60, 133) <= 5; angryBirdLarge(60, 134) <= 5; angryBirdLarge(60, 135) <= 5; angryBirdLarge(60, 136) <= 5; angryBirdLarge(60, 137) <= 5; angryBirdLarge(60, 138) <= 5; angryBirdLarge(60, 139) <= 5; angryBirdLarge(60, 140) <= 5; angryBirdLarge(60, 141) <= 5; angryBirdLarge(60, 142) <= 5; angryBirdLarge(60, 143) <= 5; angryBirdLarge(60, 144) <= 0; angryBirdLarge(60, 145) <= 0; angryBirdLarge(60, 146) <= 0; angryBirdLarge(60, 147) <= 0; angryBirdLarge(60, 148) <= 0; angryBirdLarge(60, 149) <= 0; 
angryBirdLarge(61, 0) <= 0; angryBirdLarge(61, 1) <= 0; angryBirdLarge(61, 2) <= 0; angryBirdLarge(61, 3) <= 0; angryBirdLarge(61, 4) <= 0; angryBirdLarge(61, 5) <= 0; angryBirdLarge(61, 6) <= 0; angryBirdLarge(61, 7) <= 0; angryBirdLarge(61, 8) <= 0; angryBirdLarge(61, 9) <= 0; angryBirdLarge(61, 10) <= 0; angryBirdLarge(61, 11) <= 0; angryBirdLarge(61, 12) <= 0; angryBirdLarge(61, 13) <= 0; angryBirdLarge(61, 14) <= 0; angryBirdLarge(61, 15) <= 0; angryBirdLarge(61, 16) <= 0; angryBirdLarge(61, 17) <= 0; angryBirdLarge(61, 18) <= 0; angryBirdLarge(61, 19) <= 0; angryBirdLarge(61, 20) <= 0; angryBirdLarge(61, 21) <= 0; angryBirdLarge(61, 22) <= 0; angryBirdLarge(61, 23) <= 0; angryBirdLarge(61, 24) <= 0; angryBirdLarge(61, 25) <= 0; angryBirdLarge(61, 26) <= 0; angryBirdLarge(61, 27) <= 0; angryBirdLarge(61, 28) <= 0; angryBirdLarge(61, 29) <= 0; angryBirdLarge(61, 30) <= 5; angryBirdLarge(61, 31) <= 5; angryBirdLarge(61, 32) <= 5; angryBirdLarge(61, 33) <= 5; angryBirdLarge(61, 34) <= 5; angryBirdLarge(61, 35) <= 5; angryBirdLarge(61, 36) <= 4; angryBirdLarge(61, 37) <= 4; angryBirdLarge(61, 38) <= 4; angryBirdLarge(61, 39) <= 4; angryBirdLarge(61, 40) <= 4; angryBirdLarge(61, 41) <= 4; angryBirdLarge(61, 42) <= 4; angryBirdLarge(61, 43) <= 4; angryBirdLarge(61, 44) <= 4; angryBirdLarge(61, 45) <= 4; angryBirdLarge(61, 46) <= 4; angryBirdLarge(61, 47) <= 4; angryBirdLarge(61, 48) <= 4; angryBirdLarge(61, 49) <= 4; angryBirdLarge(61, 50) <= 4; angryBirdLarge(61, 51) <= 4; angryBirdLarge(61, 52) <= 4; angryBirdLarge(61, 53) <= 4; angryBirdLarge(61, 54) <= 4; angryBirdLarge(61, 55) <= 4; angryBirdLarge(61, 56) <= 4; angryBirdLarge(61, 57) <= 4; angryBirdLarge(61, 58) <= 4; angryBirdLarge(61, 59) <= 4; angryBirdLarge(61, 60) <= 4; angryBirdLarge(61, 61) <= 4; angryBirdLarge(61, 62) <= 4; angryBirdLarge(61, 63) <= 4; angryBirdLarge(61, 64) <= 4; angryBirdLarge(61, 65) <= 4; angryBirdLarge(61, 66) <= 4; angryBirdLarge(61, 67) <= 4; angryBirdLarge(61, 68) <= 4; angryBirdLarge(61, 69) <= 4; angryBirdLarge(61, 70) <= 4; angryBirdLarge(61, 71) <= 4; angryBirdLarge(61, 72) <= 5; angryBirdLarge(61, 73) <= 5; angryBirdLarge(61, 74) <= 5; angryBirdLarge(61, 75) <= 5; angryBirdLarge(61, 76) <= 5; angryBirdLarge(61, 77) <= 5; angryBirdLarge(61, 78) <= 5; angryBirdLarge(61, 79) <= 5; angryBirdLarge(61, 80) <= 5; angryBirdLarge(61, 81) <= 5; angryBirdLarge(61, 82) <= 5; angryBirdLarge(61, 83) <= 5; angryBirdLarge(61, 84) <= 5; angryBirdLarge(61, 85) <= 5; angryBirdLarge(61, 86) <= 5; angryBirdLarge(61, 87) <= 5; angryBirdLarge(61, 88) <= 5; angryBirdLarge(61, 89) <= 5; angryBirdLarge(61, 90) <= 5; angryBirdLarge(61, 91) <= 5; angryBirdLarge(61, 92) <= 5; angryBirdLarge(61, 93) <= 5; angryBirdLarge(61, 94) <= 5; angryBirdLarge(61, 95) <= 5; angryBirdLarge(61, 96) <= 4; angryBirdLarge(61, 97) <= 4; angryBirdLarge(61, 98) <= 4; angryBirdLarge(61, 99) <= 4; angryBirdLarge(61, 100) <= 4; angryBirdLarge(61, 101) <= 4; angryBirdLarge(61, 102) <= 4; angryBirdLarge(61, 103) <= 4; angryBirdLarge(61, 104) <= 4; angryBirdLarge(61, 105) <= 4; angryBirdLarge(61, 106) <= 4; angryBirdLarge(61, 107) <= 4; angryBirdLarge(61, 108) <= 4; angryBirdLarge(61, 109) <= 4; angryBirdLarge(61, 110) <= 4; angryBirdLarge(61, 111) <= 4; angryBirdLarge(61, 112) <= 4; angryBirdLarge(61, 113) <= 4; angryBirdLarge(61, 114) <= 4; angryBirdLarge(61, 115) <= 4; angryBirdLarge(61, 116) <= 4; angryBirdLarge(61, 117) <= 4; angryBirdLarge(61, 118) <= 4; angryBirdLarge(61, 119) <= 4; angryBirdLarge(61, 120) <= 4; angryBirdLarge(61, 121) <= 4; angryBirdLarge(61, 122) <= 4; angryBirdLarge(61, 123) <= 4; angryBirdLarge(61, 124) <= 4; angryBirdLarge(61, 125) <= 4; angryBirdLarge(61, 126) <= 5; angryBirdLarge(61, 127) <= 5; angryBirdLarge(61, 128) <= 5; angryBirdLarge(61, 129) <= 5; angryBirdLarge(61, 130) <= 5; angryBirdLarge(61, 131) <= 5; angryBirdLarge(61, 132) <= 5; angryBirdLarge(61, 133) <= 5; angryBirdLarge(61, 134) <= 5; angryBirdLarge(61, 135) <= 5; angryBirdLarge(61, 136) <= 5; angryBirdLarge(61, 137) <= 5; angryBirdLarge(61, 138) <= 5; angryBirdLarge(61, 139) <= 5; angryBirdLarge(61, 140) <= 5; angryBirdLarge(61, 141) <= 5; angryBirdLarge(61, 142) <= 5; angryBirdLarge(61, 143) <= 5; angryBirdLarge(61, 144) <= 0; angryBirdLarge(61, 145) <= 0; angryBirdLarge(61, 146) <= 0; angryBirdLarge(61, 147) <= 0; angryBirdLarge(61, 148) <= 0; angryBirdLarge(61, 149) <= 0; 
angryBirdLarge(62, 0) <= 0; angryBirdLarge(62, 1) <= 0; angryBirdLarge(62, 2) <= 0; angryBirdLarge(62, 3) <= 0; angryBirdLarge(62, 4) <= 0; angryBirdLarge(62, 5) <= 0; angryBirdLarge(62, 6) <= 0; angryBirdLarge(62, 7) <= 0; angryBirdLarge(62, 8) <= 0; angryBirdLarge(62, 9) <= 0; angryBirdLarge(62, 10) <= 0; angryBirdLarge(62, 11) <= 0; angryBirdLarge(62, 12) <= 0; angryBirdLarge(62, 13) <= 0; angryBirdLarge(62, 14) <= 0; angryBirdLarge(62, 15) <= 0; angryBirdLarge(62, 16) <= 0; angryBirdLarge(62, 17) <= 0; angryBirdLarge(62, 18) <= 0; angryBirdLarge(62, 19) <= 0; angryBirdLarge(62, 20) <= 0; angryBirdLarge(62, 21) <= 0; angryBirdLarge(62, 22) <= 0; angryBirdLarge(62, 23) <= 0; angryBirdLarge(62, 24) <= 0; angryBirdLarge(62, 25) <= 0; angryBirdLarge(62, 26) <= 0; angryBirdLarge(62, 27) <= 0; angryBirdLarge(62, 28) <= 0; angryBirdLarge(62, 29) <= 0; angryBirdLarge(62, 30) <= 5; angryBirdLarge(62, 31) <= 5; angryBirdLarge(62, 32) <= 5; angryBirdLarge(62, 33) <= 5; angryBirdLarge(62, 34) <= 5; angryBirdLarge(62, 35) <= 5; angryBirdLarge(62, 36) <= 4; angryBirdLarge(62, 37) <= 4; angryBirdLarge(62, 38) <= 4; angryBirdLarge(62, 39) <= 4; angryBirdLarge(62, 40) <= 4; angryBirdLarge(62, 41) <= 4; angryBirdLarge(62, 42) <= 4; angryBirdLarge(62, 43) <= 4; angryBirdLarge(62, 44) <= 4; angryBirdLarge(62, 45) <= 4; angryBirdLarge(62, 46) <= 4; angryBirdLarge(62, 47) <= 4; angryBirdLarge(62, 48) <= 4; angryBirdLarge(62, 49) <= 4; angryBirdLarge(62, 50) <= 4; angryBirdLarge(62, 51) <= 4; angryBirdLarge(62, 52) <= 4; angryBirdLarge(62, 53) <= 4; angryBirdLarge(62, 54) <= 4; angryBirdLarge(62, 55) <= 4; angryBirdLarge(62, 56) <= 4; angryBirdLarge(62, 57) <= 4; angryBirdLarge(62, 58) <= 4; angryBirdLarge(62, 59) <= 4; angryBirdLarge(62, 60) <= 4; angryBirdLarge(62, 61) <= 4; angryBirdLarge(62, 62) <= 4; angryBirdLarge(62, 63) <= 4; angryBirdLarge(62, 64) <= 4; angryBirdLarge(62, 65) <= 4; angryBirdLarge(62, 66) <= 4; angryBirdLarge(62, 67) <= 4; angryBirdLarge(62, 68) <= 4; angryBirdLarge(62, 69) <= 4; angryBirdLarge(62, 70) <= 4; angryBirdLarge(62, 71) <= 4; angryBirdLarge(62, 72) <= 5; angryBirdLarge(62, 73) <= 5; angryBirdLarge(62, 74) <= 5; angryBirdLarge(62, 75) <= 5; angryBirdLarge(62, 76) <= 5; angryBirdLarge(62, 77) <= 5; angryBirdLarge(62, 78) <= 5; angryBirdLarge(62, 79) <= 5; angryBirdLarge(62, 80) <= 5; angryBirdLarge(62, 81) <= 5; angryBirdLarge(62, 82) <= 5; angryBirdLarge(62, 83) <= 5; angryBirdLarge(62, 84) <= 5; angryBirdLarge(62, 85) <= 5; angryBirdLarge(62, 86) <= 5; angryBirdLarge(62, 87) <= 5; angryBirdLarge(62, 88) <= 5; angryBirdLarge(62, 89) <= 5; angryBirdLarge(62, 90) <= 5; angryBirdLarge(62, 91) <= 5; angryBirdLarge(62, 92) <= 5; angryBirdLarge(62, 93) <= 5; angryBirdLarge(62, 94) <= 5; angryBirdLarge(62, 95) <= 5; angryBirdLarge(62, 96) <= 4; angryBirdLarge(62, 97) <= 4; angryBirdLarge(62, 98) <= 4; angryBirdLarge(62, 99) <= 4; angryBirdLarge(62, 100) <= 4; angryBirdLarge(62, 101) <= 4; angryBirdLarge(62, 102) <= 4; angryBirdLarge(62, 103) <= 4; angryBirdLarge(62, 104) <= 4; angryBirdLarge(62, 105) <= 4; angryBirdLarge(62, 106) <= 4; angryBirdLarge(62, 107) <= 4; angryBirdLarge(62, 108) <= 4; angryBirdLarge(62, 109) <= 4; angryBirdLarge(62, 110) <= 4; angryBirdLarge(62, 111) <= 4; angryBirdLarge(62, 112) <= 4; angryBirdLarge(62, 113) <= 4; angryBirdLarge(62, 114) <= 4; angryBirdLarge(62, 115) <= 4; angryBirdLarge(62, 116) <= 4; angryBirdLarge(62, 117) <= 4; angryBirdLarge(62, 118) <= 4; angryBirdLarge(62, 119) <= 4; angryBirdLarge(62, 120) <= 4; angryBirdLarge(62, 121) <= 4; angryBirdLarge(62, 122) <= 4; angryBirdLarge(62, 123) <= 4; angryBirdLarge(62, 124) <= 4; angryBirdLarge(62, 125) <= 4; angryBirdLarge(62, 126) <= 5; angryBirdLarge(62, 127) <= 5; angryBirdLarge(62, 128) <= 5; angryBirdLarge(62, 129) <= 5; angryBirdLarge(62, 130) <= 5; angryBirdLarge(62, 131) <= 5; angryBirdLarge(62, 132) <= 5; angryBirdLarge(62, 133) <= 5; angryBirdLarge(62, 134) <= 5; angryBirdLarge(62, 135) <= 5; angryBirdLarge(62, 136) <= 5; angryBirdLarge(62, 137) <= 5; angryBirdLarge(62, 138) <= 5; angryBirdLarge(62, 139) <= 5; angryBirdLarge(62, 140) <= 5; angryBirdLarge(62, 141) <= 5; angryBirdLarge(62, 142) <= 5; angryBirdLarge(62, 143) <= 5; angryBirdLarge(62, 144) <= 0; angryBirdLarge(62, 145) <= 0; angryBirdLarge(62, 146) <= 0; angryBirdLarge(62, 147) <= 0; angryBirdLarge(62, 148) <= 0; angryBirdLarge(62, 149) <= 0; 
angryBirdLarge(63, 0) <= 0; angryBirdLarge(63, 1) <= 0; angryBirdLarge(63, 2) <= 0; angryBirdLarge(63, 3) <= 0; angryBirdLarge(63, 4) <= 0; angryBirdLarge(63, 5) <= 0; angryBirdLarge(63, 6) <= 0; angryBirdLarge(63, 7) <= 0; angryBirdLarge(63, 8) <= 0; angryBirdLarge(63, 9) <= 0; angryBirdLarge(63, 10) <= 0; angryBirdLarge(63, 11) <= 0; angryBirdLarge(63, 12) <= 0; angryBirdLarge(63, 13) <= 0; angryBirdLarge(63, 14) <= 0; angryBirdLarge(63, 15) <= 0; angryBirdLarge(63, 16) <= 0; angryBirdLarge(63, 17) <= 0; angryBirdLarge(63, 18) <= 0; angryBirdLarge(63, 19) <= 0; angryBirdLarge(63, 20) <= 0; angryBirdLarge(63, 21) <= 0; angryBirdLarge(63, 22) <= 0; angryBirdLarge(63, 23) <= 0; angryBirdLarge(63, 24) <= 0; angryBirdLarge(63, 25) <= 0; angryBirdLarge(63, 26) <= 0; angryBirdLarge(63, 27) <= 0; angryBirdLarge(63, 28) <= 0; angryBirdLarge(63, 29) <= 0; angryBirdLarge(63, 30) <= 5; angryBirdLarge(63, 31) <= 5; angryBirdLarge(63, 32) <= 5; angryBirdLarge(63, 33) <= 5; angryBirdLarge(63, 34) <= 5; angryBirdLarge(63, 35) <= 5; angryBirdLarge(63, 36) <= 4; angryBirdLarge(63, 37) <= 4; angryBirdLarge(63, 38) <= 4; angryBirdLarge(63, 39) <= 4; angryBirdLarge(63, 40) <= 4; angryBirdLarge(63, 41) <= 4; angryBirdLarge(63, 42) <= 4; angryBirdLarge(63, 43) <= 4; angryBirdLarge(63, 44) <= 4; angryBirdLarge(63, 45) <= 4; angryBirdLarge(63, 46) <= 4; angryBirdLarge(63, 47) <= 4; angryBirdLarge(63, 48) <= 4; angryBirdLarge(63, 49) <= 4; angryBirdLarge(63, 50) <= 4; angryBirdLarge(63, 51) <= 4; angryBirdLarge(63, 52) <= 4; angryBirdLarge(63, 53) <= 4; angryBirdLarge(63, 54) <= 4; angryBirdLarge(63, 55) <= 4; angryBirdLarge(63, 56) <= 4; angryBirdLarge(63, 57) <= 4; angryBirdLarge(63, 58) <= 4; angryBirdLarge(63, 59) <= 4; angryBirdLarge(63, 60) <= 4; angryBirdLarge(63, 61) <= 4; angryBirdLarge(63, 62) <= 4; angryBirdLarge(63, 63) <= 4; angryBirdLarge(63, 64) <= 4; angryBirdLarge(63, 65) <= 4; angryBirdLarge(63, 66) <= 4; angryBirdLarge(63, 67) <= 4; angryBirdLarge(63, 68) <= 4; angryBirdLarge(63, 69) <= 4; angryBirdLarge(63, 70) <= 4; angryBirdLarge(63, 71) <= 4; angryBirdLarge(63, 72) <= 5; angryBirdLarge(63, 73) <= 5; angryBirdLarge(63, 74) <= 5; angryBirdLarge(63, 75) <= 5; angryBirdLarge(63, 76) <= 5; angryBirdLarge(63, 77) <= 5; angryBirdLarge(63, 78) <= 5; angryBirdLarge(63, 79) <= 5; angryBirdLarge(63, 80) <= 5; angryBirdLarge(63, 81) <= 5; angryBirdLarge(63, 82) <= 5; angryBirdLarge(63, 83) <= 5; angryBirdLarge(63, 84) <= 5; angryBirdLarge(63, 85) <= 5; angryBirdLarge(63, 86) <= 5; angryBirdLarge(63, 87) <= 5; angryBirdLarge(63, 88) <= 5; angryBirdLarge(63, 89) <= 5; angryBirdLarge(63, 90) <= 5; angryBirdLarge(63, 91) <= 5; angryBirdLarge(63, 92) <= 5; angryBirdLarge(63, 93) <= 5; angryBirdLarge(63, 94) <= 5; angryBirdLarge(63, 95) <= 5; angryBirdLarge(63, 96) <= 4; angryBirdLarge(63, 97) <= 4; angryBirdLarge(63, 98) <= 4; angryBirdLarge(63, 99) <= 4; angryBirdLarge(63, 100) <= 4; angryBirdLarge(63, 101) <= 4; angryBirdLarge(63, 102) <= 4; angryBirdLarge(63, 103) <= 4; angryBirdLarge(63, 104) <= 4; angryBirdLarge(63, 105) <= 4; angryBirdLarge(63, 106) <= 4; angryBirdLarge(63, 107) <= 4; angryBirdLarge(63, 108) <= 4; angryBirdLarge(63, 109) <= 4; angryBirdLarge(63, 110) <= 4; angryBirdLarge(63, 111) <= 4; angryBirdLarge(63, 112) <= 4; angryBirdLarge(63, 113) <= 4; angryBirdLarge(63, 114) <= 4; angryBirdLarge(63, 115) <= 4; angryBirdLarge(63, 116) <= 4; angryBirdLarge(63, 117) <= 4; angryBirdLarge(63, 118) <= 4; angryBirdLarge(63, 119) <= 4; angryBirdLarge(63, 120) <= 4; angryBirdLarge(63, 121) <= 4; angryBirdLarge(63, 122) <= 4; angryBirdLarge(63, 123) <= 4; angryBirdLarge(63, 124) <= 4; angryBirdLarge(63, 125) <= 4; angryBirdLarge(63, 126) <= 5; angryBirdLarge(63, 127) <= 5; angryBirdLarge(63, 128) <= 5; angryBirdLarge(63, 129) <= 5; angryBirdLarge(63, 130) <= 5; angryBirdLarge(63, 131) <= 5; angryBirdLarge(63, 132) <= 5; angryBirdLarge(63, 133) <= 5; angryBirdLarge(63, 134) <= 5; angryBirdLarge(63, 135) <= 5; angryBirdLarge(63, 136) <= 5; angryBirdLarge(63, 137) <= 5; angryBirdLarge(63, 138) <= 5; angryBirdLarge(63, 139) <= 5; angryBirdLarge(63, 140) <= 5; angryBirdLarge(63, 141) <= 5; angryBirdLarge(63, 142) <= 5; angryBirdLarge(63, 143) <= 5; angryBirdLarge(63, 144) <= 0; angryBirdLarge(63, 145) <= 0; angryBirdLarge(63, 146) <= 0; angryBirdLarge(63, 147) <= 0; angryBirdLarge(63, 148) <= 0; angryBirdLarge(63, 149) <= 0; 
angryBirdLarge(64, 0) <= 0; angryBirdLarge(64, 1) <= 0; angryBirdLarge(64, 2) <= 0; angryBirdLarge(64, 3) <= 0; angryBirdLarge(64, 4) <= 0; angryBirdLarge(64, 5) <= 0; angryBirdLarge(64, 6) <= 0; angryBirdLarge(64, 7) <= 0; angryBirdLarge(64, 8) <= 0; angryBirdLarge(64, 9) <= 0; angryBirdLarge(64, 10) <= 0; angryBirdLarge(64, 11) <= 0; angryBirdLarge(64, 12) <= 0; angryBirdLarge(64, 13) <= 0; angryBirdLarge(64, 14) <= 0; angryBirdLarge(64, 15) <= 0; angryBirdLarge(64, 16) <= 0; angryBirdLarge(64, 17) <= 0; angryBirdLarge(64, 18) <= 0; angryBirdLarge(64, 19) <= 0; angryBirdLarge(64, 20) <= 0; angryBirdLarge(64, 21) <= 0; angryBirdLarge(64, 22) <= 0; angryBirdLarge(64, 23) <= 0; angryBirdLarge(64, 24) <= 0; angryBirdLarge(64, 25) <= 0; angryBirdLarge(64, 26) <= 0; angryBirdLarge(64, 27) <= 0; angryBirdLarge(64, 28) <= 0; angryBirdLarge(64, 29) <= 0; angryBirdLarge(64, 30) <= 5; angryBirdLarge(64, 31) <= 5; angryBirdLarge(64, 32) <= 5; angryBirdLarge(64, 33) <= 5; angryBirdLarge(64, 34) <= 5; angryBirdLarge(64, 35) <= 5; angryBirdLarge(64, 36) <= 4; angryBirdLarge(64, 37) <= 4; angryBirdLarge(64, 38) <= 4; angryBirdLarge(64, 39) <= 4; angryBirdLarge(64, 40) <= 4; angryBirdLarge(64, 41) <= 4; angryBirdLarge(64, 42) <= 4; angryBirdLarge(64, 43) <= 4; angryBirdLarge(64, 44) <= 4; angryBirdLarge(64, 45) <= 4; angryBirdLarge(64, 46) <= 4; angryBirdLarge(64, 47) <= 4; angryBirdLarge(64, 48) <= 4; angryBirdLarge(64, 49) <= 4; angryBirdLarge(64, 50) <= 4; angryBirdLarge(64, 51) <= 4; angryBirdLarge(64, 52) <= 4; angryBirdLarge(64, 53) <= 4; angryBirdLarge(64, 54) <= 4; angryBirdLarge(64, 55) <= 4; angryBirdLarge(64, 56) <= 4; angryBirdLarge(64, 57) <= 4; angryBirdLarge(64, 58) <= 4; angryBirdLarge(64, 59) <= 4; angryBirdLarge(64, 60) <= 4; angryBirdLarge(64, 61) <= 4; angryBirdLarge(64, 62) <= 4; angryBirdLarge(64, 63) <= 4; angryBirdLarge(64, 64) <= 4; angryBirdLarge(64, 65) <= 4; angryBirdLarge(64, 66) <= 4; angryBirdLarge(64, 67) <= 4; angryBirdLarge(64, 68) <= 4; angryBirdLarge(64, 69) <= 4; angryBirdLarge(64, 70) <= 4; angryBirdLarge(64, 71) <= 4; angryBirdLarge(64, 72) <= 5; angryBirdLarge(64, 73) <= 5; angryBirdLarge(64, 74) <= 5; angryBirdLarge(64, 75) <= 5; angryBirdLarge(64, 76) <= 5; angryBirdLarge(64, 77) <= 5; angryBirdLarge(64, 78) <= 5; angryBirdLarge(64, 79) <= 5; angryBirdLarge(64, 80) <= 5; angryBirdLarge(64, 81) <= 5; angryBirdLarge(64, 82) <= 5; angryBirdLarge(64, 83) <= 5; angryBirdLarge(64, 84) <= 5; angryBirdLarge(64, 85) <= 5; angryBirdLarge(64, 86) <= 5; angryBirdLarge(64, 87) <= 5; angryBirdLarge(64, 88) <= 5; angryBirdLarge(64, 89) <= 5; angryBirdLarge(64, 90) <= 5; angryBirdLarge(64, 91) <= 5; angryBirdLarge(64, 92) <= 5; angryBirdLarge(64, 93) <= 5; angryBirdLarge(64, 94) <= 5; angryBirdLarge(64, 95) <= 5; angryBirdLarge(64, 96) <= 4; angryBirdLarge(64, 97) <= 4; angryBirdLarge(64, 98) <= 4; angryBirdLarge(64, 99) <= 4; angryBirdLarge(64, 100) <= 4; angryBirdLarge(64, 101) <= 4; angryBirdLarge(64, 102) <= 4; angryBirdLarge(64, 103) <= 4; angryBirdLarge(64, 104) <= 4; angryBirdLarge(64, 105) <= 4; angryBirdLarge(64, 106) <= 4; angryBirdLarge(64, 107) <= 4; angryBirdLarge(64, 108) <= 4; angryBirdLarge(64, 109) <= 4; angryBirdLarge(64, 110) <= 4; angryBirdLarge(64, 111) <= 4; angryBirdLarge(64, 112) <= 4; angryBirdLarge(64, 113) <= 4; angryBirdLarge(64, 114) <= 4; angryBirdLarge(64, 115) <= 4; angryBirdLarge(64, 116) <= 4; angryBirdLarge(64, 117) <= 4; angryBirdLarge(64, 118) <= 4; angryBirdLarge(64, 119) <= 4; angryBirdLarge(64, 120) <= 4; angryBirdLarge(64, 121) <= 4; angryBirdLarge(64, 122) <= 4; angryBirdLarge(64, 123) <= 4; angryBirdLarge(64, 124) <= 4; angryBirdLarge(64, 125) <= 4; angryBirdLarge(64, 126) <= 5; angryBirdLarge(64, 127) <= 5; angryBirdLarge(64, 128) <= 5; angryBirdLarge(64, 129) <= 5; angryBirdLarge(64, 130) <= 5; angryBirdLarge(64, 131) <= 5; angryBirdLarge(64, 132) <= 5; angryBirdLarge(64, 133) <= 5; angryBirdLarge(64, 134) <= 5; angryBirdLarge(64, 135) <= 5; angryBirdLarge(64, 136) <= 5; angryBirdLarge(64, 137) <= 5; angryBirdLarge(64, 138) <= 5; angryBirdLarge(64, 139) <= 5; angryBirdLarge(64, 140) <= 5; angryBirdLarge(64, 141) <= 5; angryBirdLarge(64, 142) <= 5; angryBirdLarge(64, 143) <= 5; angryBirdLarge(64, 144) <= 0; angryBirdLarge(64, 145) <= 0; angryBirdLarge(64, 146) <= 0; angryBirdLarge(64, 147) <= 0; angryBirdLarge(64, 148) <= 0; angryBirdLarge(64, 149) <= 0; 
angryBirdLarge(65, 0) <= 0; angryBirdLarge(65, 1) <= 0; angryBirdLarge(65, 2) <= 0; angryBirdLarge(65, 3) <= 0; angryBirdLarge(65, 4) <= 0; angryBirdLarge(65, 5) <= 0; angryBirdLarge(65, 6) <= 0; angryBirdLarge(65, 7) <= 0; angryBirdLarge(65, 8) <= 0; angryBirdLarge(65, 9) <= 0; angryBirdLarge(65, 10) <= 0; angryBirdLarge(65, 11) <= 0; angryBirdLarge(65, 12) <= 0; angryBirdLarge(65, 13) <= 0; angryBirdLarge(65, 14) <= 0; angryBirdLarge(65, 15) <= 0; angryBirdLarge(65, 16) <= 0; angryBirdLarge(65, 17) <= 0; angryBirdLarge(65, 18) <= 0; angryBirdLarge(65, 19) <= 0; angryBirdLarge(65, 20) <= 0; angryBirdLarge(65, 21) <= 0; angryBirdLarge(65, 22) <= 0; angryBirdLarge(65, 23) <= 0; angryBirdLarge(65, 24) <= 0; angryBirdLarge(65, 25) <= 0; angryBirdLarge(65, 26) <= 0; angryBirdLarge(65, 27) <= 0; angryBirdLarge(65, 28) <= 0; angryBirdLarge(65, 29) <= 0; angryBirdLarge(65, 30) <= 5; angryBirdLarge(65, 31) <= 5; angryBirdLarge(65, 32) <= 5; angryBirdLarge(65, 33) <= 5; angryBirdLarge(65, 34) <= 5; angryBirdLarge(65, 35) <= 5; angryBirdLarge(65, 36) <= 4; angryBirdLarge(65, 37) <= 4; angryBirdLarge(65, 38) <= 4; angryBirdLarge(65, 39) <= 4; angryBirdLarge(65, 40) <= 4; angryBirdLarge(65, 41) <= 4; angryBirdLarge(65, 42) <= 4; angryBirdLarge(65, 43) <= 4; angryBirdLarge(65, 44) <= 4; angryBirdLarge(65, 45) <= 4; angryBirdLarge(65, 46) <= 4; angryBirdLarge(65, 47) <= 4; angryBirdLarge(65, 48) <= 4; angryBirdLarge(65, 49) <= 4; angryBirdLarge(65, 50) <= 4; angryBirdLarge(65, 51) <= 4; angryBirdLarge(65, 52) <= 4; angryBirdLarge(65, 53) <= 4; angryBirdLarge(65, 54) <= 4; angryBirdLarge(65, 55) <= 4; angryBirdLarge(65, 56) <= 4; angryBirdLarge(65, 57) <= 4; angryBirdLarge(65, 58) <= 4; angryBirdLarge(65, 59) <= 4; angryBirdLarge(65, 60) <= 4; angryBirdLarge(65, 61) <= 4; angryBirdLarge(65, 62) <= 4; angryBirdLarge(65, 63) <= 4; angryBirdLarge(65, 64) <= 4; angryBirdLarge(65, 65) <= 4; angryBirdLarge(65, 66) <= 4; angryBirdLarge(65, 67) <= 4; angryBirdLarge(65, 68) <= 4; angryBirdLarge(65, 69) <= 4; angryBirdLarge(65, 70) <= 4; angryBirdLarge(65, 71) <= 4; angryBirdLarge(65, 72) <= 5; angryBirdLarge(65, 73) <= 5; angryBirdLarge(65, 74) <= 5; angryBirdLarge(65, 75) <= 5; angryBirdLarge(65, 76) <= 5; angryBirdLarge(65, 77) <= 5; angryBirdLarge(65, 78) <= 5; angryBirdLarge(65, 79) <= 5; angryBirdLarge(65, 80) <= 5; angryBirdLarge(65, 81) <= 5; angryBirdLarge(65, 82) <= 5; angryBirdLarge(65, 83) <= 5; angryBirdLarge(65, 84) <= 5; angryBirdLarge(65, 85) <= 5; angryBirdLarge(65, 86) <= 5; angryBirdLarge(65, 87) <= 5; angryBirdLarge(65, 88) <= 5; angryBirdLarge(65, 89) <= 5; angryBirdLarge(65, 90) <= 5; angryBirdLarge(65, 91) <= 5; angryBirdLarge(65, 92) <= 5; angryBirdLarge(65, 93) <= 5; angryBirdLarge(65, 94) <= 5; angryBirdLarge(65, 95) <= 5; angryBirdLarge(65, 96) <= 4; angryBirdLarge(65, 97) <= 4; angryBirdLarge(65, 98) <= 4; angryBirdLarge(65, 99) <= 4; angryBirdLarge(65, 100) <= 4; angryBirdLarge(65, 101) <= 4; angryBirdLarge(65, 102) <= 4; angryBirdLarge(65, 103) <= 4; angryBirdLarge(65, 104) <= 4; angryBirdLarge(65, 105) <= 4; angryBirdLarge(65, 106) <= 4; angryBirdLarge(65, 107) <= 4; angryBirdLarge(65, 108) <= 4; angryBirdLarge(65, 109) <= 4; angryBirdLarge(65, 110) <= 4; angryBirdLarge(65, 111) <= 4; angryBirdLarge(65, 112) <= 4; angryBirdLarge(65, 113) <= 4; angryBirdLarge(65, 114) <= 4; angryBirdLarge(65, 115) <= 4; angryBirdLarge(65, 116) <= 4; angryBirdLarge(65, 117) <= 4; angryBirdLarge(65, 118) <= 4; angryBirdLarge(65, 119) <= 4; angryBirdLarge(65, 120) <= 4; angryBirdLarge(65, 121) <= 4; angryBirdLarge(65, 122) <= 4; angryBirdLarge(65, 123) <= 4; angryBirdLarge(65, 124) <= 4; angryBirdLarge(65, 125) <= 4; angryBirdLarge(65, 126) <= 5; angryBirdLarge(65, 127) <= 5; angryBirdLarge(65, 128) <= 5; angryBirdLarge(65, 129) <= 5; angryBirdLarge(65, 130) <= 5; angryBirdLarge(65, 131) <= 5; angryBirdLarge(65, 132) <= 5; angryBirdLarge(65, 133) <= 5; angryBirdLarge(65, 134) <= 5; angryBirdLarge(65, 135) <= 5; angryBirdLarge(65, 136) <= 5; angryBirdLarge(65, 137) <= 5; angryBirdLarge(65, 138) <= 5; angryBirdLarge(65, 139) <= 5; angryBirdLarge(65, 140) <= 5; angryBirdLarge(65, 141) <= 5; angryBirdLarge(65, 142) <= 5; angryBirdLarge(65, 143) <= 5; angryBirdLarge(65, 144) <= 0; angryBirdLarge(65, 145) <= 0; angryBirdLarge(65, 146) <= 0; angryBirdLarge(65, 147) <= 0; angryBirdLarge(65, 148) <= 0; angryBirdLarge(65, 149) <= 0; 
angryBirdLarge(66, 0) <= 5; angryBirdLarge(66, 1) <= 5; angryBirdLarge(66, 2) <= 5; angryBirdLarge(66, 3) <= 5; angryBirdLarge(66, 4) <= 5; angryBirdLarge(66, 5) <= 5; angryBirdLarge(66, 6) <= 5; angryBirdLarge(66, 7) <= 5; angryBirdLarge(66, 8) <= 5; angryBirdLarge(66, 9) <= 5; angryBirdLarge(66, 10) <= 5; angryBirdLarge(66, 11) <= 5; angryBirdLarge(66, 12) <= 5; angryBirdLarge(66, 13) <= 5; angryBirdLarge(66, 14) <= 5; angryBirdLarge(66, 15) <= 5; angryBirdLarge(66, 16) <= 5; angryBirdLarge(66, 17) <= 5; angryBirdLarge(66, 18) <= 0; angryBirdLarge(66, 19) <= 0; angryBirdLarge(66, 20) <= 0; angryBirdLarge(66, 21) <= 0; angryBirdLarge(66, 22) <= 0; angryBirdLarge(66, 23) <= 0; angryBirdLarge(66, 24) <= 5; angryBirdLarge(66, 25) <= 5; angryBirdLarge(66, 26) <= 5; angryBirdLarge(66, 27) <= 5; angryBirdLarge(66, 28) <= 5; angryBirdLarge(66, 29) <= 5; angryBirdLarge(66, 30) <= 4; angryBirdLarge(66, 31) <= 4; angryBirdLarge(66, 32) <= 4; angryBirdLarge(66, 33) <= 4; angryBirdLarge(66, 34) <= 4; angryBirdLarge(66, 35) <= 4; angryBirdLarge(66, 36) <= 4; angryBirdLarge(66, 37) <= 4; angryBirdLarge(66, 38) <= 4; angryBirdLarge(66, 39) <= 4; angryBirdLarge(66, 40) <= 4; angryBirdLarge(66, 41) <= 4; angryBirdLarge(66, 42) <= 4; angryBirdLarge(66, 43) <= 4; angryBirdLarge(66, 44) <= 4; angryBirdLarge(66, 45) <= 4; angryBirdLarge(66, 46) <= 4; angryBirdLarge(66, 47) <= 4; angryBirdLarge(66, 48) <= 4; angryBirdLarge(66, 49) <= 4; angryBirdLarge(66, 50) <= 4; angryBirdLarge(66, 51) <= 4; angryBirdLarge(66, 52) <= 4; angryBirdLarge(66, 53) <= 4; angryBirdLarge(66, 54) <= 4; angryBirdLarge(66, 55) <= 4; angryBirdLarge(66, 56) <= 4; angryBirdLarge(66, 57) <= 4; angryBirdLarge(66, 58) <= 4; angryBirdLarge(66, 59) <= 4; angryBirdLarge(66, 60) <= 4; angryBirdLarge(66, 61) <= 4; angryBirdLarge(66, 62) <= 4; angryBirdLarge(66, 63) <= 4; angryBirdLarge(66, 64) <= 4; angryBirdLarge(66, 65) <= 4; angryBirdLarge(66, 66) <= 4; angryBirdLarge(66, 67) <= 4; angryBirdLarge(66, 68) <= 4; angryBirdLarge(66, 69) <= 4; angryBirdLarge(66, 70) <= 4; angryBirdLarge(66, 71) <= 4; angryBirdLarge(66, 72) <= 4; angryBirdLarge(66, 73) <= 4; angryBirdLarge(66, 74) <= 4; angryBirdLarge(66, 75) <= 4; angryBirdLarge(66, 76) <= 4; angryBirdLarge(66, 77) <= 4; angryBirdLarge(66, 78) <= 5; angryBirdLarge(66, 79) <= 5; angryBirdLarge(66, 80) <= 5; angryBirdLarge(66, 81) <= 5; angryBirdLarge(66, 82) <= 5; angryBirdLarge(66, 83) <= 5; angryBirdLarge(66, 84) <= 5; angryBirdLarge(66, 85) <= 5; angryBirdLarge(66, 86) <= 5; angryBirdLarge(66, 87) <= 5; angryBirdLarge(66, 88) <= 5; angryBirdLarge(66, 89) <= 5; angryBirdLarge(66, 90) <= 5; angryBirdLarge(66, 91) <= 5; angryBirdLarge(66, 92) <= 5; angryBirdLarge(66, 93) <= 5; angryBirdLarge(66, 94) <= 5; angryBirdLarge(66, 95) <= 5; angryBirdLarge(66, 96) <= 5; angryBirdLarge(66, 97) <= 5; angryBirdLarge(66, 98) <= 5; angryBirdLarge(66, 99) <= 5; angryBirdLarge(66, 100) <= 5; angryBirdLarge(66, 101) <= 5; angryBirdLarge(66, 102) <= 5; angryBirdLarge(66, 103) <= 5; angryBirdLarge(66, 104) <= 5; angryBirdLarge(66, 105) <= 5; angryBirdLarge(66, 106) <= 5; angryBirdLarge(66, 107) <= 5; angryBirdLarge(66, 108) <= 4; angryBirdLarge(66, 109) <= 4; angryBirdLarge(66, 110) <= 4; angryBirdLarge(66, 111) <= 4; angryBirdLarge(66, 112) <= 4; angryBirdLarge(66, 113) <= 4; angryBirdLarge(66, 114) <= 4; angryBirdLarge(66, 115) <= 4; angryBirdLarge(66, 116) <= 4; angryBirdLarge(66, 117) <= 4; angryBirdLarge(66, 118) <= 4; angryBirdLarge(66, 119) <= 4; angryBirdLarge(66, 120) <= 5; angryBirdLarge(66, 121) <= 5; angryBirdLarge(66, 122) <= 5; angryBirdLarge(66, 123) <= 5; angryBirdLarge(66, 124) <= 5; angryBirdLarge(66, 125) <= 5; angryBirdLarge(66, 126) <= 5; angryBirdLarge(66, 127) <= 5; angryBirdLarge(66, 128) <= 5; angryBirdLarge(66, 129) <= 5; angryBirdLarge(66, 130) <= 5; angryBirdLarge(66, 131) <= 5; angryBirdLarge(66, 132) <= 5; angryBirdLarge(66, 133) <= 5; angryBirdLarge(66, 134) <= 5; angryBirdLarge(66, 135) <= 5; angryBirdLarge(66, 136) <= 5; angryBirdLarge(66, 137) <= 5; angryBirdLarge(66, 138) <= 5; angryBirdLarge(66, 139) <= 5; angryBirdLarge(66, 140) <= 5; angryBirdLarge(66, 141) <= 5; angryBirdLarge(66, 142) <= 5; angryBirdLarge(66, 143) <= 5; angryBirdLarge(66, 144) <= 5; angryBirdLarge(66, 145) <= 5; angryBirdLarge(66, 146) <= 5; angryBirdLarge(66, 147) <= 5; angryBirdLarge(66, 148) <= 5; angryBirdLarge(66, 149) <= 5; 
angryBirdLarge(67, 0) <= 5; angryBirdLarge(67, 1) <= 5; angryBirdLarge(67, 2) <= 5; angryBirdLarge(67, 3) <= 5; angryBirdLarge(67, 4) <= 5; angryBirdLarge(67, 5) <= 5; angryBirdLarge(67, 6) <= 5; angryBirdLarge(67, 7) <= 5; angryBirdLarge(67, 8) <= 5; angryBirdLarge(67, 9) <= 5; angryBirdLarge(67, 10) <= 5; angryBirdLarge(67, 11) <= 5; angryBirdLarge(67, 12) <= 5; angryBirdLarge(67, 13) <= 5; angryBirdLarge(67, 14) <= 5; angryBirdLarge(67, 15) <= 5; angryBirdLarge(67, 16) <= 5; angryBirdLarge(67, 17) <= 5; angryBirdLarge(67, 18) <= 0; angryBirdLarge(67, 19) <= 0; angryBirdLarge(67, 20) <= 0; angryBirdLarge(67, 21) <= 0; angryBirdLarge(67, 22) <= 0; angryBirdLarge(67, 23) <= 0; angryBirdLarge(67, 24) <= 5; angryBirdLarge(67, 25) <= 5; angryBirdLarge(67, 26) <= 5; angryBirdLarge(67, 27) <= 5; angryBirdLarge(67, 28) <= 5; angryBirdLarge(67, 29) <= 5; angryBirdLarge(67, 30) <= 4; angryBirdLarge(67, 31) <= 4; angryBirdLarge(67, 32) <= 4; angryBirdLarge(67, 33) <= 4; angryBirdLarge(67, 34) <= 4; angryBirdLarge(67, 35) <= 4; angryBirdLarge(67, 36) <= 4; angryBirdLarge(67, 37) <= 4; angryBirdLarge(67, 38) <= 4; angryBirdLarge(67, 39) <= 4; angryBirdLarge(67, 40) <= 4; angryBirdLarge(67, 41) <= 4; angryBirdLarge(67, 42) <= 4; angryBirdLarge(67, 43) <= 4; angryBirdLarge(67, 44) <= 4; angryBirdLarge(67, 45) <= 4; angryBirdLarge(67, 46) <= 4; angryBirdLarge(67, 47) <= 4; angryBirdLarge(67, 48) <= 4; angryBirdLarge(67, 49) <= 4; angryBirdLarge(67, 50) <= 4; angryBirdLarge(67, 51) <= 4; angryBirdLarge(67, 52) <= 4; angryBirdLarge(67, 53) <= 4; angryBirdLarge(67, 54) <= 4; angryBirdLarge(67, 55) <= 4; angryBirdLarge(67, 56) <= 4; angryBirdLarge(67, 57) <= 4; angryBirdLarge(67, 58) <= 4; angryBirdLarge(67, 59) <= 4; angryBirdLarge(67, 60) <= 4; angryBirdLarge(67, 61) <= 4; angryBirdLarge(67, 62) <= 4; angryBirdLarge(67, 63) <= 4; angryBirdLarge(67, 64) <= 4; angryBirdLarge(67, 65) <= 4; angryBirdLarge(67, 66) <= 4; angryBirdLarge(67, 67) <= 4; angryBirdLarge(67, 68) <= 4; angryBirdLarge(67, 69) <= 4; angryBirdLarge(67, 70) <= 4; angryBirdLarge(67, 71) <= 4; angryBirdLarge(67, 72) <= 4; angryBirdLarge(67, 73) <= 4; angryBirdLarge(67, 74) <= 4; angryBirdLarge(67, 75) <= 4; angryBirdLarge(67, 76) <= 4; angryBirdLarge(67, 77) <= 4; angryBirdLarge(67, 78) <= 5; angryBirdLarge(67, 79) <= 5; angryBirdLarge(67, 80) <= 5; angryBirdLarge(67, 81) <= 5; angryBirdLarge(67, 82) <= 5; angryBirdLarge(67, 83) <= 5; angryBirdLarge(67, 84) <= 5; angryBirdLarge(67, 85) <= 5; angryBirdLarge(67, 86) <= 5; angryBirdLarge(67, 87) <= 5; angryBirdLarge(67, 88) <= 5; angryBirdLarge(67, 89) <= 5; angryBirdLarge(67, 90) <= 5; angryBirdLarge(67, 91) <= 5; angryBirdLarge(67, 92) <= 5; angryBirdLarge(67, 93) <= 5; angryBirdLarge(67, 94) <= 5; angryBirdLarge(67, 95) <= 5; angryBirdLarge(67, 96) <= 5; angryBirdLarge(67, 97) <= 5; angryBirdLarge(67, 98) <= 5; angryBirdLarge(67, 99) <= 5; angryBirdLarge(67, 100) <= 5; angryBirdLarge(67, 101) <= 5; angryBirdLarge(67, 102) <= 5; angryBirdLarge(67, 103) <= 5; angryBirdLarge(67, 104) <= 5; angryBirdLarge(67, 105) <= 5; angryBirdLarge(67, 106) <= 5; angryBirdLarge(67, 107) <= 5; angryBirdLarge(67, 108) <= 4; angryBirdLarge(67, 109) <= 4; angryBirdLarge(67, 110) <= 4; angryBirdLarge(67, 111) <= 4; angryBirdLarge(67, 112) <= 4; angryBirdLarge(67, 113) <= 4; angryBirdLarge(67, 114) <= 4; angryBirdLarge(67, 115) <= 4; angryBirdLarge(67, 116) <= 4; angryBirdLarge(67, 117) <= 4; angryBirdLarge(67, 118) <= 4; angryBirdLarge(67, 119) <= 4; angryBirdLarge(67, 120) <= 5; angryBirdLarge(67, 121) <= 5; angryBirdLarge(67, 122) <= 5; angryBirdLarge(67, 123) <= 5; angryBirdLarge(67, 124) <= 5; angryBirdLarge(67, 125) <= 5; angryBirdLarge(67, 126) <= 5; angryBirdLarge(67, 127) <= 5; angryBirdLarge(67, 128) <= 5; angryBirdLarge(67, 129) <= 5; angryBirdLarge(67, 130) <= 5; angryBirdLarge(67, 131) <= 5; angryBirdLarge(67, 132) <= 5; angryBirdLarge(67, 133) <= 5; angryBirdLarge(67, 134) <= 5; angryBirdLarge(67, 135) <= 5; angryBirdLarge(67, 136) <= 5; angryBirdLarge(67, 137) <= 5; angryBirdLarge(67, 138) <= 5; angryBirdLarge(67, 139) <= 5; angryBirdLarge(67, 140) <= 5; angryBirdLarge(67, 141) <= 5; angryBirdLarge(67, 142) <= 5; angryBirdLarge(67, 143) <= 5; angryBirdLarge(67, 144) <= 5; angryBirdLarge(67, 145) <= 5; angryBirdLarge(67, 146) <= 5; angryBirdLarge(67, 147) <= 5; angryBirdLarge(67, 148) <= 5; angryBirdLarge(67, 149) <= 5; 
angryBirdLarge(68, 0) <= 5; angryBirdLarge(68, 1) <= 5; angryBirdLarge(68, 2) <= 5; angryBirdLarge(68, 3) <= 5; angryBirdLarge(68, 4) <= 5; angryBirdLarge(68, 5) <= 5; angryBirdLarge(68, 6) <= 5; angryBirdLarge(68, 7) <= 5; angryBirdLarge(68, 8) <= 5; angryBirdLarge(68, 9) <= 5; angryBirdLarge(68, 10) <= 5; angryBirdLarge(68, 11) <= 5; angryBirdLarge(68, 12) <= 5; angryBirdLarge(68, 13) <= 5; angryBirdLarge(68, 14) <= 5; angryBirdLarge(68, 15) <= 5; angryBirdLarge(68, 16) <= 5; angryBirdLarge(68, 17) <= 5; angryBirdLarge(68, 18) <= 0; angryBirdLarge(68, 19) <= 0; angryBirdLarge(68, 20) <= 0; angryBirdLarge(68, 21) <= 0; angryBirdLarge(68, 22) <= 0; angryBirdLarge(68, 23) <= 0; angryBirdLarge(68, 24) <= 5; angryBirdLarge(68, 25) <= 5; angryBirdLarge(68, 26) <= 5; angryBirdLarge(68, 27) <= 5; angryBirdLarge(68, 28) <= 5; angryBirdLarge(68, 29) <= 5; angryBirdLarge(68, 30) <= 4; angryBirdLarge(68, 31) <= 4; angryBirdLarge(68, 32) <= 4; angryBirdLarge(68, 33) <= 4; angryBirdLarge(68, 34) <= 4; angryBirdLarge(68, 35) <= 4; angryBirdLarge(68, 36) <= 4; angryBirdLarge(68, 37) <= 4; angryBirdLarge(68, 38) <= 4; angryBirdLarge(68, 39) <= 4; angryBirdLarge(68, 40) <= 4; angryBirdLarge(68, 41) <= 4; angryBirdLarge(68, 42) <= 4; angryBirdLarge(68, 43) <= 4; angryBirdLarge(68, 44) <= 4; angryBirdLarge(68, 45) <= 4; angryBirdLarge(68, 46) <= 4; angryBirdLarge(68, 47) <= 4; angryBirdLarge(68, 48) <= 4; angryBirdLarge(68, 49) <= 4; angryBirdLarge(68, 50) <= 4; angryBirdLarge(68, 51) <= 4; angryBirdLarge(68, 52) <= 4; angryBirdLarge(68, 53) <= 4; angryBirdLarge(68, 54) <= 4; angryBirdLarge(68, 55) <= 4; angryBirdLarge(68, 56) <= 4; angryBirdLarge(68, 57) <= 4; angryBirdLarge(68, 58) <= 4; angryBirdLarge(68, 59) <= 4; angryBirdLarge(68, 60) <= 4; angryBirdLarge(68, 61) <= 4; angryBirdLarge(68, 62) <= 4; angryBirdLarge(68, 63) <= 4; angryBirdLarge(68, 64) <= 4; angryBirdLarge(68, 65) <= 4; angryBirdLarge(68, 66) <= 4; angryBirdLarge(68, 67) <= 4; angryBirdLarge(68, 68) <= 4; angryBirdLarge(68, 69) <= 4; angryBirdLarge(68, 70) <= 4; angryBirdLarge(68, 71) <= 4; angryBirdLarge(68, 72) <= 4; angryBirdLarge(68, 73) <= 4; angryBirdLarge(68, 74) <= 4; angryBirdLarge(68, 75) <= 4; angryBirdLarge(68, 76) <= 4; angryBirdLarge(68, 77) <= 4; angryBirdLarge(68, 78) <= 5; angryBirdLarge(68, 79) <= 5; angryBirdLarge(68, 80) <= 5; angryBirdLarge(68, 81) <= 5; angryBirdLarge(68, 82) <= 5; angryBirdLarge(68, 83) <= 5; angryBirdLarge(68, 84) <= 5; angryBirdLarge(68, 85) <= 5; angryBirdLarge(68, 86) <= 5; angryBirdLarge(68, 87) <= 5; angryBirdLarge(68, 88) <= 5; angryBirdLarge(68, 89) <= 5; angryBirdLarge(68, 90) <= 5; angryBirdLarge(68, 91) <= 5; angryBirdLarge(68, 92) <= 5; angryBirdLarge(68, 93) <= 5; angryBirdLarge(68, 94) <= 5; angryBirdLarge(68, 95) <= 5; angryBirdLarge(68, 96) <= 5; angryBirdLarge(68, 97) <= 5; angryBirdLarge(68, 98) <= 5; angryBirdLarge(68, 99) <= 5; angryBirdLarge(68, 100) <= 5; angryBirdLarge(68, 101) <= 5; angryBirdLarge(68, 102) <= 5; angryBirdLarge(68, 103) <= 5; angryBirdLarge(68, 104) <= 5; angryBirdLarge(68, 105) <= 5; angryBirdLarge(68, 106) <= 5; angryBirdLarge(68, 107) <= 5; angryBirdLarge(68, 108) <= 4; angryBirdLarge(68, 109) <= 4; angryBirdLarge(68, 110) <= 4; angryBirdLarge(68, 111) <= 4; angryBirdLarge(68, 112) <= 4; angryBirdLarge(68, 113) <= 4; angryBirdLarge(68, 114) <= 4; angryBirdLarge(68, 115) <= 4; angryBirdLarge(68, 116) <= 4; angryBirdLarge(68, 117) <= 4; angryBirdLarge(68, 118) <= 4; angryBirdLarge(68, 119) <= 4; angryBirdLarge(68, 120) <= 5; angryBirdLarge(68, 121) <= 5; angryBirdLarge(68, 122) <= 5; angryBirdLarge(68, 123) <= 5; angryBirdLarge(68, 124) <= 5; angryBirdLarge(68, 125) <= 5; angryBirdLarge(68, 126) <= 5; angryBirdLarge(68, 127) <= 5; angryBirdLarge(68, 128) <= 5; angryBirdLarge(68, 129) <= 5; angryBirdLarge(68, 130) <= 5; angryBirdLarge(68, 131) <= 5; angryBirdLarge(68, 132) <= 5; angryBirdLarge(68, 133) <= 5; angryBirdLarge(68, 134) <= 5; angryBirdLarge(68, 135) <= 5; angryBirdLarge(68, 136) <= 5; angryBirdLarge(68, 137) <= 5; angryBirdLarge(68, 138) <= 5; angryBirdLarge(68, 139) <= 5; angryBirdLarge(68, 140) <= 5; angryBirdLarge(68, 141) <= 5; angryBirdLarge(68, 142) <= 5; angryBirdLarge(68, 143) <= 5; angryBirdLarge(68, 144) <= 5; angryBirdLarge(68, 145) <= 5; angryBirdLarge(68, 146) <= 5; angryBirdLarge(68, 147) <= 5; angryBirdLarge(68, 148) <= 5; angryBirdLarge(68, 149) <= 5; 
angryBirdLarge(69, 0) <= 5; angryBirdLarge(69, 1) <= 5; angryBirdLarge(69, 2) <= 5; angryBirdLarge(69, 3) <= 5; angryBirdLarge(69, 4) <= 5; angryBirdLarge(69, 5) <= 5; angryBirdLarge(69, 6) <= 5; angryBirdLarge(69, 7) <= 5; angryBirdLarge(69, 8) <= 5; angryBirdLarge(69, 9) <= 5; angryBirdLarge(69, 10) <= 5; angryBirdLarge(69, 11) <= 5; angryBirdLarge(69, 12) <= 5; angryBirdLarge(69, 13) <= 5; angryBirdLarge(69, 14) <= 5; angryBirdLarge(69, 15) <= 5; angryBirdLarge(69, 16) <= 5; angryBirdLarge(69, 17) <= 5; angryBirdLarge(69, 18) <= 0; angryBirdLarge(69, 19) <= 0; angryBirdLarge(69, 20) <= 0; angryBirdLarge(69, 21) <= 0; angryBirdLarge(69, 22) <= 0; angryBirdLarge(69, 23) <= 0; angryBirdLarge(69, 24) <= 5; angryBirdLarge(69, 25) <= 5; angryBirdLarge(69, 26) <= 5; angryBirdLarge(69, 27) <= 5; angryBirdLarge(69, 28) <= 5; angryBirdLarge(69, 29) <= 5; angryBirdLarge(69, 30) <= 4; angryBirdLarge(69, 31) <= 4; angryBirdLarge(69, 32) <= 4; angryBirdLarge(69, 33) <= 4; angryBirdLarge(69, 34) <= 4; angryBirdLarge(69, 35) <= 4; angryBirdLarge(69, 36) <= 4; angryBirdLarge(69, 37) <= 4; angryBirdLarge(69, 38) <= 4; angryBirdLarge(69, 39) <= 4; angryBirdLarge(69, 40) <= 4; angryBirdLarge(69, 41) <= 4; angryBirdLarge(69, 42) <= 4; angryBirdLarge(69, 43) <= 4; angryBirdLarge(69, 44) <= 4; angryBirdLarge(69, 45) <= 4; angryBirdLarge(69, 46) <= 4; angryBirdLarge(69, 47) <= 4; angryBirdLarge(69, 48) <= 4; angryBirdLarge(69, 49) <= 4; angryBirdLarge(69, 50) <= 4; angryBirdLarge(69, 51) <= 4; angryBirdLarge(69, 52) <= 4; angryBirdLarge(69, 53) <= 4; angryBirdLarge(69, 54) <= 4; angryBirdLarge(69, 55) <= 4; angryBirdLarge(69, 56) <= 4; angryBirdLarge(69, 57) <= 4; angryBirdLarge(69, 58) <= 4; angryBirdLarge(69, 59) <= 4; angryBirdLarge(69, 60) <= 4; angryBirdLarge(69, 61) <= 4; angryBirdLarge(69, 62) <= 4; angryBirdLarge(69, 63) <= 4; angryBirdLarge(69, 64) <= 4; angryBirdLarge(69, 65) <= 4; angryBirdLarge(69, 66) <= 4; angryBirdLarge(69, 67) <= 4; angryBirdLarge(69, 68) <= 4; angryBirdLarge(69, 69) <= 4; angryBirdLarge(69, 70) <= 4; angryBirdLarge(69, 71) <= 4; angryBirdLarge(69, 72) <= 4; angryBirdLarge(69, 73) <= 4; angryBirdLarge(69, 74) <= 4; angryBirdLarge(69, 75) <= 4; angryBirdLarge(69, 76) <= 4; angryBirdLarge(69, 77) <= 4; angryBirdLarge(69, 78) <= 5; angryBirdLarge(69, 79) <= 5; angryBirdLarge(69, 80) <= 5; angryBirdLarge(69, 81) <= 5; angryBirdLarge(69, 82) <= 5; angryBirdLarge(69, 83) <= 5; angryBirdLarge(69, 84) <= 5; angryBirdLarge(69, 85) <= 5; angryBirdLarge(69, 86) <= 5; angryBirdLarge(69, 87) <= 5; angryBirdLarge(69, 88) <= 5; angryBirdLarge(69, 89) <= 5; angryBirdLarge(69, 90) <= 5; angryBirdLarge(69, 91) <= 5; angryBirdLarge(69, 92) <= 5; angryBirdLarge(69, 93) <= 5; angryBirdLarge(69, 94) <= 5; angryBirdLarge(69, 95) <= 5; angryBirdLarge(69, 96) <= 5; angryBirdLarge(69, 97) <= 5; angryBirdLarge(69, 98) <= 5; angryBirdLarge(69, 99) <= 5; angryBirdLarge(69, 100) <= 5; angryBirdLarge(69, 101) <= 5; angryBirdLarge(69, 102) <= 5; angryBirdLarge(69, 103) <= 5; angryBirdLarge(69, 104) <= 5; angryBirdLarge(69, 105) <= 5; angryBirdLarge(69, 106) <= 5; angryBirdLarge(69, 107) <= 5; angryBirdLarge(69, 108) <= 4; angryBirdLarge(69, 109) <= 4; angryBirdLarge(69, 110) <= 4; angryBirdLarge(69, 111) <= 4; angryBirdLarge(69, 112) <= 4; angryBirdLarge(69, 113) <= 4; angryBirdLarge(69, 114) <= 4; angryBirdLarge(69, 115) <= 4; angryBirdLarge(69, 116) <= 4; angryBirdLarge(69, 117) <= 4; angryBirdLarge(69, 118) <= 4; angryBirdLarge(69, 119) <= 4; angryBirdLarge(69, 120) <= 5; angryBirdLarge(69, 121) <= 5; angryBirdLarge(69, 122) <= 5; angryBirdLarge(69, 123) <= 5; angryBirdLarge(69, 124) <= 5; angryBirdLarge(69, 125) <= 5; angryBirdLarge(69, 126) <= 5; angryBirdLarge(69, 127) <= 5; angryBirdLarge(69, 128) <= 5; angryBirdLarge(69, 129) <= 5; angryBirdLarge(69, 130) <= 5; angryBirdLarge(69, 131) <= 5; angryBirdLarge(69, 132) <= 5; angryBirdLarge(69, 133) <= 5; angryBirdLarge(69, 134) <= 5; angryBirdLarge(69, 135) <= 5; angryBirdLarge(69, 136) <= 5; angryBirdLarge(69, 137) <= 5; angryBirdLarge(69, 138) <= 5; angryBirdLarge(69, 139) <= 5; angryBirdLarge(69, 140) <= 5; angryBirdLarge(69, 141) <= 5; angryBirdLarge(69, 142) <= 5; angryBirdLarge(69, 143) <= 5; angryBirdLarge(69, 144) <= 5; angryBirdLarge(69, 145) <= 5; angryBirdLarge(69, 146) <= 5; angryBirdLarge(69, 147) <= 5; angryBirdLarge(69, 148) <= 5; angryBirdLarge(69, 149) <= 5; 
angryBirdLarge(70, 0) <= 5; angryBirdLarge(70, 1) <= 5; angryBirdLarge(70, 2) <= 5; angryBirdLarge(70, 3) <= 5; angryBirdLarge(70, 4) <= 5; angryBirdLarge(70, 5) <= 5; angryBirdLarge(70, 6) <= 5; angryBirdLarge(70, 7) <= 5; angryBirdLarge(70, 8) <= 5; angryBirdLarge(70, 9) <= 5; angryBirdLarge(70, 10) <= 5; angryBirdLarge(70, 11) <= 5; angryBirdLarge(70, 12) <= 5; angryBirdLarge(70, 13) <= 5; angryBirdLarge(70, 14) <= 5; angryBirdLarge(70, 15) <= 5; angryBirdLarge(70, 16) <= 5; angryBirdLarge(70, 17) <= 5; angryBirdLarge(70, 18) <= 0; angryBirdLarge(70, 19) <= 0; angryBirdLarge(70, 20) <= 0; angryBirdLarge(70, 21) <= 0; angryBirdLarge(70, 22) <= 0; angryBirdLarge(70, 23) <= 0; angryBirdLarge(70, 24) <= 5; angryBirdLarge(70, 25) <= 5; angryBirdLarge(70, 26) <= 5; angryBirdLarge(70, 27) <= 5; angryBirdLarge(70, 28) <= 5; angryBirdLarge(70, 29) <= 5; angryBirdLarge(70, 30) <= 4; angryBirdLarge(70, 31) <= 4; angryBirdLarge(70, 32) <= 4; angryBirdLarge(70, 33) <= 4; angryBirdLarge(70, 34) <= 4; angryBirdLarge(70, 35) <= 4; angryBirdLarge(70, 36) <= 4; angryBirdLarge(70, 37) <= 4; angryBirdLarge(70, 38) <= 4; angryBirdLarge(70, 39) <= 4; angryBirdLarge(70, 40) <= 4; angryBirdLarge(70, 41) <= 4; angryBirdLarge(70, 42) <= 4; angryBirdLarge(70, 43) <= 4; angryBirdLarge(70, 44) <= 4; angryBirdLarge(70, 45) <= 4; angryBirdLarge(70, 46) <= 4; angryBirdLarge(70, 47) <= 4; angryBirdLarge(70, 48) <= 4; angryBirdLarge(70, 49) <= 4; angryBirdLarge(70, 50) <= 4; angryBirdLarge(70, 51) <= 4; angryBirdLarge(70, 52) <= 4; angryBirdLarge(70, 53) <= 4; angryBirdLarge(70, 54) <= 4; angryBirdLarge(70, 55) <= 4; angryBirdLarge(70, 56) <= 4; angryBirdLarge(70, 57) <= 4; angryBirdLarge(70, 58) <= 4; angryBirdLarge(70, 59) <= 4; angryBirdLarge(70, 60) <= 4; angryBirdLarge(70, 61) <= 4; angryBirdLarge(70, 62) <= 4; angryBirdLarge(70, 63) <= 4; angryBirdLarge(70, 64) <= 4; angryBirdLarge(70, 65) <= 4; angryBirdLarge(70, 66) <= 4; angryBirdLarge(70, 67) <= 4; angryBirdLarge(70, 68) <= 4; angryBirdLarge(70, 69) <= 4; angryBirdLarge(70, 70) <= 4; angryBirdLarge(70, 71) <= 4; angryBirdLarge(70, 72) <= 4; angryBirdLarge(70, 73) <= 4; angryBirdLarge(70, 74) <= 4; angryBirdLarge(70, 75) <= 4; angryBirdLarge(70, 76) <= 4; angryBirdLarge(70, 77) <= 4; angryBirdLarge(70, 78) <= 5; angryBirdLarge(70, 79) <= 5; angryBirdLarge(70, 80) <= 5; angryBirdLarge(70, 81) <= 5; angryBirdLarge(70, 82) <= 5; angryBirdLarge(70, 83) <= 5; angryBirdLarge(70, 84) <= 5; angryBirdLarge(70, 85) <= 5; angryBirdLarge(70, 86) <= 5; angryBirdLarge(70, 87) <= 5; angryBirdLarge(70, 88) <= 5; angryBirdLarge(70, 89) <= 5; angryBirdLarge(70, 90) <= 5; angryBirdLarge(70, 91) <= 5; angryBirdLarge(70, 92) <= 5; angryBirdLarge(70, 93) <= 5; angryBirdLarge(70, 94) <= 5; angryBirdLarge(70, 95) <= 5; angryBirdLarge(70, 96) <= 5; angryBirdLarge(70, 97) <= 5; angryBirdLarge(70, 98) <= 5; angryBirdLarge(70, 99) <= 5; angryBirdLarge(70, 100) <= 5; angryBirdLarge(70, 101) <= 5; angryBirdLarge(70, 102) <= 5; angryBirdLarge(70, 103) <= 5; angryBirdLarge(70, 104) <= 5; angryBirdLarge(70, 105) <= 5; angryBirdLarge(70, 106) <= 5; angryBirdLarge(70, 107) <= 5; angryBirdLarge(70, 108) <= 4; angryBirdLarge(70, 109) <= 4; angryBirdLarge(70, 110) <= 4; angryBirdLarge(70, 111) <= 4; angryBirdLarge(70, 112) <= 4; angryBirdLarge(70, 113) <= 4; angryBirdLarge(70, 114) <= 4; angryBirdLarge(70, 115) <= 4; angryBirdLarge(70, 116) <= 4; angryBirdLarge(70, 117) <= 4; angryBirdLarge(70, 118) <= 4; angryBirdLarge(70, 119) <= 4; angryBirdLarge(70, 120) <= 5; angryBirdLarge(70, 121) <= 5; angryBirdLarge(70, 122) <= 5; angryBirdLarge(70, 123) <= 5; angryBirdLarge(70, 124) <= 5; angryBirdLarge(70, 125) <= 5; angryBirdLarge(70, 126) <= 5; angryBirdLarge(70, 127) <= 5; angryBirdLarge(70, 128) <= 5; angryBirdLarge(70, 129) <= 5; angryBirdLarge(70, 130) <= 5; angryBirdLarge(70, 131) <= 5; angryBirdLarge(70, 132) <= 5; angryBirdLarge(70, 133) <= 5; angryBirdLarge(70, 134) <= 5; angryBirdLarge(70, 135) <= 5; angryBirdLarge(70, 136) <= 5; angryBirdLarge(70, 137) <= 5; angryBirdLarge(70, 138) <= 5; angryBirdLarge(70, 139) <= 5; angryBirdLarge(70, 140) <= 5; angryBirdLarge(70, 141) <= 5; angryBirdLarge(70, 142) <= 5; angryBirdLarge(70, 143) <= 5; angryBirdLarge(70, 144) <= 5; angryBirdLarge(70, 145) <= 5; angryBirdLarge(70, 146) <= 5; angryBirdLarge(70, 147) <= 5; angryBirdLarge(70, 148) <= 5; angryBirdLarge(70, 149) <= 5; 
angryBirdLarge(71, 0) <= 5; angryBirdLarge(71, 1) <= 5; angryBirdLarge(71, 2) <= 5; angryBirdLarge(71, 3) <= 5; angryBirdLarge(71, 4) <= 5; angryBirdLarge(71, 5) <= 5; angryBirdLarge(71, 6) <= 5; angryBirdLarge(71, 7) <= 5; angryBirdLarge(71, 8) <= 5; angryBirdLarge(71, 9) <= 5; angryBirdLarge(71, 10) <= 5; angryBirdLarge(71, 11) <= 5; angryBirdLarge(71, 12) <= 5; angryBirdLarge(71, 13) <= 5; angryBirdLarge(71, 14) <= 5; angryBirdLarge(71, 15) <= 5; angryBirdLarge(71, 16) <= 5; angryBirdLarge(71, 17) <= 5; angryBirdLarge(71, 18) <= 0; angryBirdLarge(71, 19) <= 0; angryBirdLarge(71, 20) <= 0; angryBirdLarge(71, 21) <= 0; angryBirdLarge(71, 22) <= 0; angryBirdLarge(71, 23) <= 0; angryBirdLarge(71, 24) <= 5; angryBirdLarge(71, 25) <= 5; angryBirdLarge(71, 26) <= 5; angryBirdLarge(71, 27) <= 5; angryBirdLarge(71, 28) <= 5; angryBirdLarge(71, 29) <= 5; angryBirdLarge(71, 30) <= 4; angryBirdLarge(71, 31) <= 4; angryBirdLarge(71, 32) <= 4; angryBirdLarge(71, 33) <= 4; angryBirdLarge(71, 34) <= 4; angryBirdLarge(71, 35) <= 4; angryBirdLarge(71, 36) <= 4; angryBirdLarge(71, 37) <= 4; angryBirdLarge(71, 38) <= 4; angryBirdLarge(71, 39) <= 4; angryBirdLarge(71, 40) <= 4; angryBirdLarge(71, 41) <= 4; angryBirdLarge(71, 42) <= 4; angryBirdLarge(71, 43) <= 4; angryBirdLarge(71, 44) <= 4; angryBirdLarge(71, 45) <= 4; angryBirdLarge(71, 46) <= 4; angryBirdLarge(71, 47) <= 4; angryBirdLarge(71, 48) <= 4; angryBirdLarge(71, 49) <= 4; angryBirdLarge(71, 50) <= 4; angryBirdLarge(71, 51) <= 4; angryBirdLarge(71, 52) <= 4; angryBirdLarge(71, 53) <= 4; angryBirdLarge(71, 54) <= 4; angryBirdLarge(71, 55) <= 4; angryBirdLarge(71, 56) <= 4; angryBirdLarge(71, 57) <= 4; angryBirdLarge(71, 58) <= 4; angryBirdLarge(71, 59) <= 4; angryBirdLarge(71, 60) <= 4; angryBirdLarge(71, 61) <= 4; angryBirdLarge(71, 62) <= 4; angryBirdLarge(71, 63) <= 4; angryBirdLarge(71, 64) <= 4; angryBirdLarge(71, 65) <= 4; angryBirdLarge(71, 66) <= 4; angryBirdLarge(71, 67) <= 4; angryBirdLarge(71, 68) <= 4; angryBirdLarge(71, 69) <= 4; angryBirdLarge(71, 70) <= 4; angryBirdLarge(71, 71) <= 4; angryBirdLarge(71, 72) <= 4; angryBirdLarge(71, 73) <= 4; angryBirdLarge(71, 74) <= 4; angryBirdLarge(71, 75) <= 4; angryBirdLarge(71, 76) <= 4; angryBirdLarge(71, 77) <= 4; angryBirdLarge(71, 78) <= 5; angryBirdLarge(71, 79) <= 5; angryBirdLarge(71, 80) <= 5; angryBirdLarge(71, 81) <= 5; angryBirdLarge(71, 82) <= 5; angryBirdLarge(71, 83) <= 5; angryBirdLarge(71, 84) <= 5; angryBirdLarge(71, 85) <= 5; angryBirdLarge(71, 86) <= 5; angryBirdLarge(71, 87) <= 5; angryBirdLarge(71, 88) <= 5; angryBirdLarge(71, 89) <= 5; angryBirdLarge(71, 90) <= 5; angryBirdLarge(71, 91) <= 5; angryBirdLarge(71, 92) <= 5; angryBirdLarge(71, 93) <= 5; angryBirdLarge(71, 94) <= 5; angryBirdLarge(71, 95) <= 5; angryBirdLarge(71, 96) <= 5; angryBirdLarge(71, 97) <= 5; angryBirdLarge(71, 98) <= 5; angryBirdLarge(71, 99) <= 5; angryBirdLarge(71, 100) <= 5; angryBirdLarge(71, 101) <= 5; angryBirdLarge(71, 102) <= 5; angryBirdLarge(71, 103) <= 5; angryBirdLarge(71, 104) <= 5; angryBirdLarge(71, 105) <= 5; angryBirdLarge(71, 106) <= 5; angryBirdLarge(71, 107) <= 5; angryBirdLarge(71, 108) <= 4; angryBirdLarge(71, 109) <= 4; angryBirdLarge(71, 110) <= 4; angryBirdLarge(71, 111) <= 4; angryBirdLarge(71, 112) <= 4; angryBirdLarge(71, 113) <= 4; angryBirdLarge(71, 114) <= 4; angryBirdLarge(71, 115) <= 4; angryBirdLarge(71, 116) <= 4; angryBirdLarge(71, 117) <= 4; angryBirdLarge(71, 118) <= 4; angryBirdLarge(71, 119) <= 4; angryBirdLarge(71, 120) <= 5; angryBirdLarge(71, 121) <= 5; angryBirdLarge(71, 122) <= 5; angryBirdLarge(71, 123) <= 5; angryBirdLarge(71, 124) <= 5; angryBirdLarge(71, 125) <= 5; angryBirdLarge(71, 126) <= 5; angryBirdLarge(71, 127) <= 5; angryBirdLarge(71, 128) <= 5; angryBirdLarge(71, 129) <= 5; angryBirdLarge(71, 130) <= 5; angryBirdLarge(71, 131) <= 5; angryBirdLarge(71, 132) <= 5; angryBirdLarge(71, 133) <= 5; angryBirdLarge(71, 134) <= 5; angryBirdLarge(71, 135) <= 5; angryBirdLarge(71, 136) <= 5; angryBirdLarge(71, 137) <= 5; angryBirdLarge(71, 138) <= 5; angryBirdLarge(71, 139) <= 5; angryBirdLarge(71, 140) <= 5; angryBirdLarge(71, 141) <= 5; angryBirdLarge(71, 142) <= 5; angryBirdLarge(71, 143) <= 5; angryBirdLarge(71, 144) <= 5; angryBirdLarge(71, 145) <= 5; angryBirdLarge(71, 146) <= 5; angryBirdLarge(71, 147) <= 5; angryBirdLarge(71, 148) <= 5; angryBirdLarge(71, 149) <= 5; 
angryBirdLarge(72, 0) <= 0; angryBirdLarge(72, 1) <= 0; angryBirdLarge(72, 2) <= 0; angryBirdLarge(72, 3) <= 0; angryBirdLarge(72, 4) <= 0; angryBirdLarge(72, 5) <= 0; angryBirdLarge(72, 6) <= 5; angryBirdLarge(72, 7) <= 5; angryBirdLarge(72, 8) <= 5; angryBirdLarge(72, 9) <= 5; angryBirdLarge(72, 10) <= 5; angryBirdLarge(72, 11) <= 5; angryBirdLarge(72, 12) <= 5; angryBirdLarge(72, 13) <= 5; angryBirdLarge(72, 14) <= 5; angryBirdLarge(72, 15) <= 5; angryBirdLarge(72, 16) <= 5; angryBirdLarge(72, 17) <= 5; angryBirdLarge(72, 18) <= 5; angryBirdLarge(72, 19) <= 5; angryBirdLarge(72, 20) <= 5; angryBirdLarge(72, 21) <= 5; angryBirdLarge(72, 22) <= 5; angryBirdLarge(72, 23) <= 5; angryBirdLarge(72, 24) <= 5; angryBirdLarge(72, 25) <= 5; angryBirdLarge(72, 26) <= 5; angryBirdLarge(72, 27) <= 5; angryBirdLarge(72, 28) <= 5; angryBirdLarge(72, 29) <= 5; angryBirdLarge(72, 30) <= 4; angryBirdLarge(72, 31) <= 4; angryBirdLarge(72, 32) <= 4; angryBirdLarge(72, 33) <= 4; angryBirdLarge(72, 34) <= 4; angryBirdLarge(72, 35) <= 4; angryBirdLarge(72, 36) <= 4; angryBirdLarge(72, 37) <= 4; angryBirdLarge(72, 38) <= 4; angryBirdLarge(72, 39) <= 4; angryBirdLarge(72, 40) <= 4; angryBirdLarge(72, 41) <= 4; angryBirdLarge(72, 42) <= 4; angryBirdLarge(72, 43) <= 4; angryBirdLarge(72, 44) <= 4; angryBirdLarge(72, 45) <= 4; angryBirdLarge(72, 46) <= 4; angryBirdLarge(72, 47) <= 4; angryBirdLarge(72, 48) <= 4; angryBirdLarge(72, 49) <= 4; angryBirdLarge(72, 50) <= 4; angryBirdLarge(72, 51) <= 4; angryBirdLarge(72, 52) <= 4; angryBirdLarge(72, 53) <= 4; angryBirdLarge(72, 54) <= 4; angryBirdLarge(72, 55) <= 4; angryBirdLarge(72, 56) <= 4; angryBirdLarge(72, 57) <= 4; angryBirdLarge(72, 58) <= 4; angryBirdLarge(72, 59) <= 4; angryBirdLarge(72, 60) <= 4; angryBirdLarge(72, 61) <= 4; angryBirdLarge(72, 62) <= 4; angryBirdLarge(72, 63) <= 4; angryBirdLarge(72, 64) <= 4; angryBirdLarge(72, 65) <= 4; angryBirdLarge(72, 66) <= 4; angryBirdLarge(72, 67) <= 4; angryBirdLarge(72, 68) <= 4; angryBirdLarge(72, 69) <= 4; angryBirdLarge(72, 70) <= 4; angryBirdLarge(72, 71) <= 4; angryBirdLarge(72, 72) <= 4; angryBirdLarge(72, 73) <= 4; angryBirdLarge(72, 74) <= 4; angryBirdLarge(72, 75) <= 4; angryBirdLarge(72, 76) <= 4; angryBirdLarge(72, 77) <= 4; angryBirdLarge(72, 78) <= 5; angryBirdLarge(72, 79) <= 5; angryBirdLarge(72, 80) <= 5; angryBirdLarge(72, 81) <= 5; angryBirdLarge(72, 82) <= 5; angryBirdLarge(72, 83) <= 5; angryBirdLarge(72, 84) <= 2; angryBirdLarge(72, 85) <= 2; angryBirdLarge(72, 86) <= 2; angryBirdLarge(72, 87) <= 2; angryBirdLarge(72, 88) <= 2; angryBirdLarge(72, 89) <= 2; angryBirdLarge(72, 90) <= 2; angryBirdLarge(72, 91) <= 2; angryBirdLarge(72, 92) <= 2; angryBirdLarge(72, 93) <= 2; angryBirdLarge(72, 94) <= 2; angryBirdLarge(72, 95) <= 2; angryBirdLarge(72, 96) <= 5; angryBirdLarge(72, 97) <= 5; angryBirdLarge(72, 98) <= 5; angryBirdLarge(72, 99) <= 5; angryBirdLarge(72, 100) <= 5; angryBirdLarge(72, 101) <= 5; angryBirdLarge(72, 102) <= 5; angryBirdLarge(72, 103) <= 5; angryBirdLarge(72, 104) <= 5; angryBirdLarge(72, 105) <= 5; angryBirdLarge(72, 106) <= 5; angryBirdLarge(72, 107) <= 5; angryBirdLarge(72, 108) <= 5; angryBirdLarge(72, 109) <= 5; angryBirdLarge(72, 110) <= 5; angryBirdLarge(72, 111) <= 5; angryBirdLarge(72, 112) <= 5; angryBirdLarge(72, 113) <= 5; angryBirdLarge(72, 114) <= 5; angryBirdLarge(72, 115) <= 5; angryBirdLarge(72, 116) <= 5; angryBirdLarge(72, 117) <= 5; angryBirdLarge(72, 118) <= 5; angryBirdLarge(72, 119) <= 5; angryBirdLarge(72, 120) <= 5; angryBirdLarge(72, 121) <= 5; angryBirdLarge(72, 122) <= 5; angryBirdLarge(72, 123) <= 5; angryBirdLarge(72, 124) <= 5; angryBirdLarge(72, 125) <= 5; angryBirdLarge(72, 126) <= 5; angryBirdLarge(72, 127) <= 5; angryBirdLarge(72, 128) <= 5; angryBirdLarge(72, 129) <= 5; angryBirdLarge(72, 130) <= 5; angryBirdLarge(72, 131) <= 5; angryBirdLarge(72, 132) <= 5; angryBirdLarge(72, 133) <= 5; angryBirdLarge(72, 134) <= 5; angryBirdLarge(72, 135) <= 5; angryBirdLarge(72, 136) <= 5; angryBirdLarge(72, 137) <= 5; angryBirdLarge(72, 138) <= 4; angryBirdLarge(72, 139) <= 4; angryBirdLarge(72, 140) <= 4; angryBirdLarge(72, 141) <= 4; angryBirdLarge(72, 142) <= 4; angryBirdLarge(72, 143) <= 4; angryBirdLarge(72, 144) <= 5; angryBirdLarge(72, 145) <= 5; angryBirdLarge(72, 146) <= 5; angryBirdLarge(72, 147) <= 5; angryBirdLarge(72, 148) <= 5; angryBirdLarge(72, 149) <= 5; 
angryBirdLarge(73, 0) <= 0; angryBirdLarge(73, 1) <= 0; angryBirdLarge(73, 2) <= 0; angryBirdLarge(73, 3) <= 0; angryBirdLarge(73, 4) <= 0; angryBirdLarge(73, 5) <= 0; angryBirdLarge(73, 6) <= 5; angryBirdLarge(73, 7) <= 5; angryBirdLarge(73, 8) <= 5; angryBirdLarge(73, 9) <= 5; angryBirdLarge(73, 10) <= 5; angryBirdLarge(73, 11) <= 5; angryBirdLarge(73, 12) <= 5; angryBirdLarge(73, 13) <= 5; angryBirdLarge(73, 14) <= 5; angryBirdLarge(73, 15) <= 5; angryBirdLarge(73, 16) <= 5; angryBirdLarge(73, 17) <= 5; angryBirdLarge(73, 18) <= 5; angryBirdLarge(73, 19) <= 5; angryBirdLarge(73, 20) <= 5; angryBirdLarge(73, 21) <= 5; angryBirdLarge(73, 22) <= 5; angryBirdLarge(73, 23) <= 5; angryBirdLarge(73, 24) <= 5; angryBirdLarge(73, 25) <= 5; angryBirdLarge(73, 26) <= 5; angryBirdLarge(73, 27) <= 5; angryBirdLarge(73, 28) <= 5; angryBirdLarge(73, 29) <= 5; angryBirdLarge(73, 30) <= 4; angryBirdLarge(73, 31) <= 4; angryBirdLarge(73, 32) <= 4; angryBirdLarge(73, 33) <= 4; angryBirdLarge(73, 34) <= 4; angryBirdLarge(73, 35) <= 4; angryBirdLarge(73, 36) <= 4; angryBirdLarge(73, 37) <= 4; angryBirdLarge(73, 38) <= 4; angryBirdLarge(73, 39) <= 4; angryBirdLarge(73, 40) <= 4; angryBirdLarge(73, 41) <= 4; angryBirdLarge(73, 42) <= 4; angryBirdLarge(73, 43) <= 4; angryBirdLarge(73, 44) <= 4; angryBirdLarge(73, 45) <= 4; angryBirdLarge(73, 46) <= 4; angryBirdLarge(73, 47) <= 4; angryBirdLarge(73, 48) <= 4; angryBirdLarge(73, 49) <= 4; angryBirdLarge(73, 50) <= 4; angryBirdLarge(73, 51) <= 4; angryBirdLarge(73, 52) <= 4; angryBirdLarge(73, 53) <= 4; angryBirdLarge(73, 54) <= 4; angryBirdLarge(73, 55) <= 4; angryBirdLarge(73, 56) <= 4; angryBirdLarge(73, 57) <= 4; angryBirdLarge(73, 58) <= 4; angryBirdLarge(73, 59) <= 4; angryBirdLarge(73, 60) <= 4; angryBirdLarge(73, 61) <= 4; angryBirdLarge(73, 62) <= 4; angryBirdLarge(73, 63) <= 4; angryBirdLarge(73, 64) <= 4; angryBirdLarge(73, 65) <= 4; angryBirdLarge(73, 66) <= 4; angryBirdLarge(73, 67) <= 4; angryBirdLarge(73, 68) <= 4; angryBirdLarge(73, 69) <= 4; angryBirdLarge(73, 70) <= 4; angryBirdLarge(73, 71) <= 4; angryBirdLarge(73, 72) <= 4; angryBirdLarge(73, 73) <= 4; angryBirdLarge(73, 74) <= 4; angryBirdLarge(73, 75) <= 4; angryBirdLarge(73, 76) <= 4; angryBirdLarge(73, 77) <= 4; angryBirdLarge(73, 78) <= 5; angryBirdLarge(73, 79) <= 5; angryBirdLarge(73, 80) <= 5; angryBirdLarge(73, 81) <= 5; angryBirdLarge(73, 82) <= 5; angryBirdLarge(73, 83) <= 5; angryBirdLarge(73, 84) <= 2; angryBirdLarge(73, 85) <= 2; angryBirdLarge(73, 86) <= 2; angryBirdLarge(73, 87) <= 2; angryBirdLarge(73, 88) <= 2; angryBirdLarge(73, 89) <= 2; angryBirdLarge(73, 90) <= 2; angryBirdLarge(73, 91) <= 2; angryBirdLarge(73, 92) <= 2; angryBirdLarge(73, 93) <= 2; angryBirdLarge(73, 94) <= 2; angryBirdLarge(73, 95) <= 2; angryBirdLarge(73, 96) <= 5; angryBirdLarge(73, 97) <= 5; angryBirdLarge(73, 98) <= 5; angryBirdLarge(73, 99) <= 5; angryBirdLarge(73, 100) <= 5; angryBirdLarge(73, 101) <= 5; angryBirdLarge(73, 102) <= 5; angryBirdLarge(73, 103) <= 5; angryBirdLarge(73, 104) <= 5; angryBirdLarge(73, 105) <= 5; angryBirdLarge(73, 106) <= 5; angryBirdLarge(73, 107) <= 5; angryBirdLarge(73, 108) <= 5; angryBirdLarge(73, 109) <= 5; angryBirdLarge(73, 110) <= 5; angryBirdLarge(73, 111) <= 5; angryBirdLarge(73, 112) <= 5; angryBirdLarge(73, 113) <= 5; angryBirdLarge(73, 114) <= 5; angryBirdLarge(73, 115) <= 5; angryBirdLarge(73, 116) <= 5; angryBirdLarge(73, 117) <= 5; angryBirdLarge(73, 118) <= 5; angryBirdLarge(73, 119) <= 5; angryBirdLarge(73, 120) <= 5; angryBirdLarge(73, 121) <= 5; angryBirdLarge(73, 122) <= 5; angryBirdLarge(73, 123) <= 5; angryBirdLarge(73, 124) <= 5; angryBirdLarge(73, 125) <= 5; angryBirdLarge(73, 126) <= 5; angryBirdLarge(73, 127) <= 5; angryBirdLarge(73, 128) <= 5; angryBirdLarge(73, 129) <= 5; angryBirdLarge(73, 130) <= 5; angryBirdLarge(73, 131) <= 5; angryBirdLarge(73, 132) <= 5; angryBirdLarge(73, 133) <= 5; angryBirdLarge(73, 134) <= 5; angryBirdLarge(73, 135) <= 5; angryBirdLarge(73, 136) <= 5; angryBirdLarge(73, 137) <= 5; angryBirdLarge(73, 138) <= 4; angryBirdLarge(73, 139) <= 4; angryBirdLarge(73, 140) <= 4; angryBirdLarge(73, 141) <= 4; angryBirdLarge(73, 142) <= 4; angryBirdLarge(73, 143) <= 4; angryBirdLarge(73, 144) <= 5; angryBirdLarge(73, 145) <= 5; angryBirdLarge(73, 146) <= 5; angryBirdLarge(73, 147) <= 5; angryBirdLarge(73, 148) <= 5; angryBirdLarge(73, 149) <= 5; 
angryBirdLarge(74, 0) <= 0; angryBirdLarge(74, 1) <= 0; angryBirdLarge(74, 2) <= 0; angryBirdLarge(74, 3) <= 0; angryBirdLarge(74, 4) <= 0; angryBirdLarge(74, 5) <= 0; angryBirdLarge(74, 6) <= 5; angryBirdLarge(74, 7) <= 5; angryBirdLarge(74, 8) <= 5; angryBirdLarge(74, 9) <= 5; angryBirdLarge(74, 10) <= 5; angryBirdLarge(74, 11) <= 5; angryBirdLarge(74, 12) <= 5; angryBirdLarge(74, 13) <= 5; angryBirdLarge(74, 14) <= 5; angryBirdLarge(74, 15) <= 5; angryBirdLarge(74, 16) <= 5; angryBirdLarge(74, 17) <= 5; angryBirdLarge(74, 18) <= 5; angryBirdLarge(74, 19) <= 5; angryBirdLarge(74, 20) <= 5; angryBirdLarge(74, 21) <= 5; angryBirdLarge(74, 22) <= 5; angryBirdLarge(74, 23) <= 5; angryBirdLarge(74, 24) <= 5; angryBirdLarge(74, 25) <= 5; angryBirdLarge(74, 26) <= 5; angryBirdLarge(74, 27) <= 5; angryBirdLarge(74, 28) <= 5; angryBirdLarge(74, 29) <= 5; angryBirdLarge(74, 30) <= 4; angryBirdLarge(74, 31) <= 4; angryBirdLarge(74, 32) <= 4; angryBirdLarge(74, 33) <= 4; angryBirdLarge(74, 34) <= 4; angryBirdLarge(74, 35) <= 4; angryBirdLarge(74, 36) <= 4; angryBirdLarge(74, 37) <= 4; angryBirdLarge(74, 38) <= 4; angryBirdLarge(74, 39) <= 4; angryBirdLarge(74, 40) <= 4; angryBirdLarge(74, 41) <= 4; angryBirdLarge(74, 42) <= 4; angryBirdLarge(74, 43) <= 4; angryBirdLarge(74, 44) <= 4; angryBirdLarge(74, 45) <= 4; angryBirdLarge(74, 46) <= 4; angryBirdLarge(74, 47) <= 4; angryBirdLarge(74, 48) <= 4; angryBirdLarge(74, 49) <= 4; angryBirdLarge(74, 50) <= 4; angryBirdLarge(74, 51) <= 4; angryBirdLarge(74, 52) <= 4; angryBirdLarge(74, 53) <= 4; angryBirdLarge(74, 54) <= 4; angryBirdLarge(74, 55) <= 4; angryBirdLarge(74, 56) <= 4; angryBirdLarge(74, 57) <= 4; angryBirdLarge(74, 58) <= 4; angryBirdLarge(74, 59) <= 4; angryBirdLarge(74, 60) <= 4; angryBirdLarge(74, 61) <= 4; angryBirdLarge(74, 62) <= 4; angryBirdLarge(74, 63) <= 4; angryBirdLarge(74, 64) <= 4; angryBirdLarge(74, 65) <= 4; angryBirdLarge(74, 66) <= 4; angryBirdLarge(74, 67) <= 4; angryBirdLarge(74, 68) <= 4; angryBirdLarge(74, 69) <= 4; angryBirdLarge(74, 70) <= 4; angryBirdLarge(74, 71) <= 4; angryBirdLarge(74, 72) <= 4; angryBirdLarge(74, 73) <= 4; angryBirdLarge(74, 74) <= 4; angryBirdLarge(74, 75) <= 4; angryBirdLarge(74, 76) <= 4; angryBirdLarge(74, 77) <= 4; angryBirdLarge(74, 78) <= 5; angryBirdLarge(74, 79) <= 5; angryBirdLarge(74, 80) <= 5; angryBirdLarge(74, 81) <= 5; angryBirdLarge(74, 82) <= 5; angryBirdLarge(74, 83) <= 5; angryBirdLarge(74, 84) <= 2; angryBirdLarge(74, 85) <= 2; angryBirdLarge(74, 86) <= 2; angryBirdLarge(74, 87) <= 2; angryBirdLarge(74, 88) <= 2; angryBirdLarge(74, 89) <= 2; angryBirdLarge(74, 90) <= 2; angryBirdLarge(74, 91) <= 2; angryBirdLarge(74, 92) <= 2; angryBirdLarge(74, 93) <= 2; angryBirdLarge(74, 94) <= 2; angryBirdLarge(74, 95) <= 2; angryBirdLarge(74, 96) <= 5; angryBirdLarge(74, 97) <= 5; angryBirdLarge(74, 98) <= 5; angryBirdLarge(74, 99) <= 5; angryBirdLarge(74, 100) <= 5; angryBirdLarge(74, 101) <= 5; angryBirdLarge(74, 102) <= 5; angryBirdLarge(74, 103) <= 5; angryBirdLarge(74, 104) <= 5; angryBirdLarge(74, 105) <= 5; angryBirdLarge(74, 106) <= 5; angryBirdLarge(74, 107) <= 5; angryBirdLarge(74, 108) <= 5; angryBirdLarge(74, 109) <= 5; angryBirdLarge(74, 110) <= 5; angryBirdLarge(74, 111) <= 5; angryBirdLarge(74, 112) <= 5; angryBirdLarge(74, 113) <= 5; angryBirdLarge(74, 114) <= 5; angryBirdLarge(74, 115) <= 5; angryBirdLarge(74, 116) <= 5; angryBirdLarge(74, 117) <= 5; angryBirdLarge(74, 118) <= 5; angryBirdLarge(74, 119) <= 5; angryBirdLarge(74, 120) <= 5; angryBirdLarge(74, 121) <= 5; angryBirdLarge(74, 122) <= 5; angryBirdLarge(74, 123) <= 5; angryBirdLarge(74, 124) <= 5; angryBirdLarge(74, 125) <= 5; angryBirdLarge(74, 126) <= 5; angryBirdLarge(74, 127) <= 5; angryBirdLarge(74, 128) <= 5; angryBirdLarge(74, 129) <= 5; angryBirdLarge(74, 130) <= 5; angryBirdLarge(74, 131) <= 5; angryBirdLarge(74, 132) <= 5; angryBirdLarge(74, 133) <= 5; angryBirdLarge(74, 134) <= 5; angryBirdLarge(74, 135) <= 5; angryBirdLarge(74, 136) <= 5; angryBirdLarge(74, 137) <= 5; angryBirdLarge(74, 138) <= 4; angryBirdLarge(74, 139) <= 4; angryBirdLarge(74, 140) <= 4; angryBirdLarge(74, 141) <= 4; angryBirdLarge(74, 142) <= 4; angryBirdLarge(74, 143) <= 4; angryBirdLarge(74, 144) <= 5; angryBirdLarge(74, 145) <= 5; angryBirdLarge(74, 146) <= 5; angryBirdLarge(74, 147) <= 5; angryBirdLarge(74, 148) <= 5; angryBirdLarge(74, 149) <= 5; 
angryBirdLarge(75, 0) <= 0; angryBirdLarge(75, 1) <= 0; angryBirdLarge(75, 2) <= 0; angryBirdLarge(75, 3) <= 0; angryBirdLarge(75, 4) <= 0; angryBirdLarge(75, 5) <= 0; angryBirdLarge(75, 6) <= 5; angryBirdLarge(75, 7) <= 5; angryBirdLarge(75, 8) <= 5; angryBirdLarge(75, 9) <= 5; angryBirdLarge(75, 10) <= 5; angryBirdLarge(75, 11) <= 5; angryBirdLarge(75, 12) <= 5; angryBirdLarge(75, 13) <= 5; angryBirdLarge(75, 14) <= 5; angryBirdLarge(75, 15) <= 5; angryBirdLarge(75, 16) <= 5; angryBirdLarge(75, 17) <= 5; angryBirdLarge(75, 18) <= 5; angryBirdLarge(75, 19) <= 5; angryBirdLarge(75, 20) <= 5; angryBirdLarge(75, 21) <= 5; angryBirdLarge(75, 22) <= 5; angryBirdLarge(75, 23) <= 5; angryBirdLarge(75, 24) <= 5; angryBirdLarge(75, 25) <= 5; angryBirdLarge(75, 26) <= 5; angryBirdLarge(75, 27) <= 5; angryBirdLarge(75, 28) <= 5; angryBirdLarge(75, 29) <= 5; angryBirdLarge(75, 30) <= 4; angryBirdLarge(75, 31) <= 4; angryBirdLarge(75, 32) <= 4; angryBirdLarge(75, 33) <= 4; angryBirdLarge(75, 34) <= 4; angryBirdLarge(75, 35) <= 4; angryBirdLarge(75, 36) <= 4; angryBirdLarge(75, 37) <= 4; angryBirdLarge(75, 38) <= 4; angryBirdLarge(75, 39) <= 4; angryBirdLarge(75, 40) <= 4; angryBirdLarge(75, 41) <= 4; angryBirdLarge(75, 42) <= 4; angryBirdLarge(75, 43) <= 4; angryBirdLarge(75, 44) <= 4; angryBirdLarge(75, 45) <= 4; angryBirdLarge(75, 46) <= 4; angryBirdLarge(75, 47) <= 4; angryBirdLarge(75, 48) <= 4; angryBirdLarge(75, 49) <= 4; angryBirdLarge(75, 50) <= 4; angryBirdLarge(75, 51) <= 4; angryBirdLarge(75, 52) <= 4; angryBirdLarge(75, 53) <= 4; angryBirdLarge(75, 54) <= 4; angryBirdLarge(75, 55) <= 4; angryBirdLarge(75, 56) <= 4; angryBirdLarge(75, 57) <= 4; angryBirdLarge(75, 58) <= 4; angryBirdLarge(75, 59) <= 4; angryBirdLarge(75, 60) <= 4; angryBirdLarge(75, 61) <= 4; angryBirdLarge(75, 62) <= 4; angryBirdLarge(75, 63) <= 4; angryBirdLarge(75, 64) <= 4; angryBirdLarge(75, 65) <= 4; angryBirdLarge(75, 66) <= 4; angryBirdLarge(75, 67) <= 4; angryBirdLarge(75, 68) <= 4; angryBirdLarge(75, 69) <= 4; angryBirdLarge(75, 70) <= 4; angryBirdLarge(75, 71) <= 4; angryBirdLarge(75, 72) <= 4; angryBirdLarge(75, 73) <= 4; angryBirdLarge(75, 74) <= 4; angryBirdLarge(75, 75) <= 4; angryBirdLarge(75, 76) <= 4; angryBirdLarge(75, 77) <= 4; angryBirdLarge(75, 78) <= 5; angryBirdLarge(75, 79) <= 5; angryBirdLarge(75, 80) <= 5; angryBirdLarge(75, 81) <= 5; angryBirdLarge(75, 82) <= 5; angryBirdLarge(75, 83) <= 5; angryBirdLarge(75, 84) <= 2; angryBirdLarge(75, 85) <= 2; angryBirdLarge(75, 86) <= 2; angryBirdLarge(75, 87) <= 2; angryBirdLarge(75, 88) <= 2; angryBirdLarge(75, 89) <= 2; angryBirdLarge(75, 90) <= 2; angryBirdLarge(75, 91) <= 2; angryBirdLarge(75, 92) <= 2; angryBirdLarge(75, 93) <= 2; angryBirdLarge(75, 94) <= 2; angryBirdLarge(75, 95) <= 2; angryBirdLarge(75, 96) <= 5; angryBirdLarge(75, 97) <= 5; angryBirdLarge(75, 98) <= 5; angryBirdLarge(75, 99) <= 5; angryBirdLarge(75, 100) <= 5; angryBirdLarge(75, 101) <= 5; angryBirdLarge(75, 102) <= 5; angryBirdLarge(75, 103) <= 5; angryBirdLarge(75, 104) <= 5; angryBirdLarge(75, 105) <= 5; angryBirdLarge(75, 106) <= 5; angryBirdLarge(75, 107) <= 5; angryBirdLarge(75, 108) <= 5; angryBirdLarge(75, 109) <= 5; angryBirdLarge(75, 110) <= 5; angryBirdLarge(75, 111) <= 5; angryBirdLarge(75, 112) <= 5; angryBirdLarge(75, 113) <= 5; angryBirdLarge(75, 114) <= 5; angryBirdLarge(75, 115) <= 5; angryBirdLarge(75, 116) <= 5; angryBirdLarge(75, 117) <= 5; angryBirdLarge(75, 118) <= 5; angryBirdLarge(75, 119) <= 5; angryBirdLarge(75, 120) <= 5; angryBirdLarge(75, 121) <= 5; angryBirdLarge(75, 122) <= 5; angryBirdLarge(75, 123) <= 5; angryBirdLarge(75, 124) <= 5; angryBirdLarge(75, 125) <= 5; angryBirdLarge(75, 126) <= 5; angryBirdLarge(75, 127) <= 5; angryBirdLarge(75, 128) <= 5; angryBirdLarge(75, 129) <= 5; angryBirdLarge(75, 130) <= 5; angryBirdLarge(75, 131) <= 5; angryBirdLarge(75, 132) <= 5; angryBirdLarge(75, 133) <= 5; angryBirdLarge(75, 134) <= 5; angryBirdLarge(75, 135) <= 5; angryBirdLarge(75, 136) <= 5; angryBirdLarge(75, 137) <= 5; angryBirdLarge(75, 138) <= 4; angryBirdLarge(75, 139) <= 4; angryBirdLarge(75, 140) <= 4; angryBirdLarge(75, 141) <= 4; angryBirdLarge(75, 142) <= 4; angryBirdLarge(75, 143) <= 4; angryBirdLarge(75, 144) <= 5; angryBirdLarge(75, 145) <= 5; angryBirdLarge(75, 146) <= 5; angryBirdLarge(75, 147) <= 5; angryBirdLarge(75, 148) <= 5; angryBirdLarge(75, 149) <= 5; 
angryBirdLarge(76, 0) <= 0; angryBirdLarge(76, 1) <= 0; angryBirdLarge(76, 2) <= 0; angryBirdLarge(76, 3) <= 0; angryBirdLarge(76, 4) <= 0; angryBirdLarge(76, 5) <= 0; angryBirdLarge(76, 6) <= 5; angryBirdLarge(76, 7) <= 5; angryBirdLarge(76, 8) <= 5; angryBirdLarge(76, 9) <= 5; angryBirdLarge(76, 10) <= 5; angryBirdLarge(76, 11) <= 5; angryBirdLarge(76, 12) <= 5; angryBirdLarge(76, 13) <= 5; angryBirdLarge(76, 14) <= 5; angryBirdLarge(76, 15) <= 5; angryBirdLarge(76, 16) <= 5; angryBirdLarge(76, 17) <= 5; angryBirdLarge(76, 18) <= 5; angryBirdLarge(76, 19) <= 5; angryBirdLarge(76, 20) <= 5; angryBirdLarge(76, 21) <= 5; angryBirdLarge(76, 22) <= 5; angryBirdLarge(76, 23) <= 5; angryBirdLarge(76, 24) <= 5; angryBirdLarge(76, 25) <= 5; angryBirdLarge(76, 26) <= 5; angryBirdLarge(76, 27) <= 5; angryBirdLarge(76, 28) <= 5; angryBirdLarge(76, 29) <= 5; angryBirdLarge(76, 30) <= 4; angryBirdLarge(76, 31) <= 4; angryBirdLarge(76, 32) <= 4; angryBirdLarge(76, 33) <= 4; angryBirdLarge(76, 34) <= 4; angryBirdLarge(76, 35) <= 4; angryBirdLarge(76, 36) <= 4; angryBirdLarge(76, 37) <= 4; angryBirdLarge(76, 38) <= 4; angryBirdLarge(76, 39) <= 4; angryBirdLarge(76, 40) <= 4; angryBirdLarge(76, 41) <= 4; angryBirdLarge(76, 42) <= 4; angryBirdLarge(76, 43) <= 4; angryBirdLarge(76, 44) <= 4; angryBirdLarge(76, 45) <= 4; angryBirdLarge(76, 46) <= 4; angryBirdLarge(76, 47) <= 4; angryBirdLarge(76, 48) <= 4; angryBirdLarge(76, 49) <= 4; angryBirdLarge(76, 50) <= 4; angryBirdLarge(76, 51) <= 4; angryBirdLarge(76, 52) <= 4; angryBirdLarge(76, 53) <= 4; angryBirdLarge(76, 54) <= 4; angryBirdLarge(76, 55) <= 4; angryBirdLarge(76, 56) <= 4; angryBirdLarge(76, 57) <= 4; angryBirdLarge(76, 58) <= 4; angryBirdLarge(76, 59) <= 4; angryBirdLarge(76, 60) <= 4; angryBirdLarge(76, 61) <= 4; angryBirdLarge(76, 62) <= 4; angryBirdLarge(76, 63) <= 4; angryBirdLarge(76, 64) <= 4; angryBirdLarge(76, 65) <= 4; angryBirdLarge(76, 66) <= 4; angryBirdLarge(76, 67) <= 4; angryBirdLarge(76, 68) <= 4; angryBirdLarge(76, 69) <= 4; angryBirdLarge(76, 70) <= 4; angryBirdLarge(76, 71) <= 4; angryBirdLarge(76, 72) <= 4; angryBirdLarge(76, 73) <= 4; angryBirdLarge(76, 74) <= 4; angryBirdLarge(76, 75) <= 4; angryBirdLarge(76, 76) <= 4; angryBirdLarge(76, 77) <= 4; angryBirdLarge(76, 78) <= 5; angryBirdLarge(76, 79) <= 5; angryBirdLarge(76, 80) <= 5; angryBirdLarge(76, 81) <= 5; angryBirdLarge(76, 82) <= 5; angryBirdLarge(76, 83) <= 5; angryBirdLarge(76, 84) <= 2; angryBirdLarge(76, 85) <= 2; angryBirdLarge(76, 86) <= 2; angryBirdLarge(76, 87) <= 2; angryBirdLarge(76, 88) <= 2; angryBirdLarge(76, 89) <= 2; angryBirdLarge(76, 90) <= 2; angryBirdLarge(76, 91) <= 2; angryBirdLarge(76, 92) <= 2; angryBirdLarge(76, 93) <= 2; angryBirdLarge(76, 94) <= 2; angryBirdLarge(76, 95) <= 2; angryBirdLarge(76, 96) <= 5; angryBirdLarge(76, 97) <= 5; angryBirdLarge(76, 98) <= 5; angryBirdLarge(76, 99) <= 5; angryBirdLarge(76, 100) <= 5; angryBirdLarge(76, 101) <= 5; angryBirdLarge(76, 102) <= 5; angryBirdLarge(76, 103) <= 5; angryBirdLarge(76, 104) <= 5; angryBirdLarge(76, 105) <= 5; angryBirdLarge(76, 106) <= 5; angryBirdLarge(76, 107) <= 5; angryBirdLarge(76, 108) <= 5; angryBirdLarge(76, 109) <= 5; angryBirdLarge(76, 110) <= 5; angryBirdLarge(76, 111) <= 5; angryBirdLarge(76, 112) <= 5; angryBirdLarge(76, 113) <= 5; angryBirdLarge(76, 114) <= 5; angryBirdLarge(76, 115) <= 5; angryBirdLarge(76, 116) <= 5; angryBirdLarge(76, 117) <= 5; angryBirdLarge(76, 118) <= 5; angryBirdLarge(76, 119) <= 5; angryBirdLarge(76, 120) <= 5; angryBirdLarge(76, 121) <= 5; angryBirdLarge(76, 122) <= 5; angryBirdLarge(76, 123) <= 5; angryBirdLarge(76, 124) <= 5; angryBirdLarge(76, 125) <= 5; angryBirdLarge(76, 126) <= 5; angryBirdLarge(76, 127) <= 5; angryBirdLarge(76, 128) <= 5; angryBirdLarge(76, 129) <= 5; angryBirdLarge(76, 130) <= 5; angryBirdLarge(76, 131) <= 5; angryBirdLarge(76, 132) <= 5; angryBirdLarge(76, 133) <= 5; angryBirdLarge(76, 134) <= 5; angryBirdLarge(76, 135) <= 5; angryBirdLarge(76, 136) <= 5; angryBirdLarge(76, 137) <= 5; angryBirdLarge(76, 138) <= 4; angryBirdLarge(76, 139) <= 4; angryBirdLarge(76, 140) <= 4; angryBirdLarge(76, 141) <= 4; angryBirdLarge(76, 142) <= 4; angryBirdLarge(76, 143) <= 4; angryBirdLarge(76, 144) <= 5; angryBirdLarge(76, 145) <= 5; angryBirdLarge(76, 146) <= 5; angryBirdLarge(76, 147) <= 5; angryBirdLarge(76, 148) <= 5; angryBirdLarge(76, 149) <= 5; 
angryBirdLarge(77, 0) <= 0; angryBirdLarge(77, 1) <= 0; angryBirdLarge(77, 2) <= 0; angryBirdLarge(77, 3) <= 0; angryBirdLarge(77, 4) <= 0; angryBirdLarge(77, 5) <= 0; angryBirdLarge(77, 6) <= 5; angryBirdLarge(77, 7) <= 5; angryBirdLarge(77, 8) <= 5; angryBirdLarge(77, 9) <= 5; angryBirdLarge(77, 10) <= 5; angryBirdLarge(77, 11) <= 5; angryBirdLarge(77, 12) <= 5; angryBirdLarge(77, 13) <= 5; angryBirdLarge(77, 14) <= 5; angryBirdLarge(77, 15) <= 5; angryBirdLarge(77, 16) <= 5; angryBirdLarge(77, 17) <= 5; angryBirdLarge(77, 18) <= 5; angryBirdLarge(77, 19) <= 5; angryBirdLarge(77, 20) <= 5; angryBirdLarge(77, 21) <= 5; angryBirdLarge(77, 22) <= 5; angryBirdLarge(77, 23) <= 5; angryBirdLarge(77, 24) <= 5; angryBirdLarge(77, 25) <= 5; angryBirdLarge(77, 26) <= 5; angryBirdLarge(77, 27) <= 5; angryBirdLarge(77, 28) <= 5; angryBirdLarge(77, 29) <= 5; angryBirdLarge(77, 30) <= 4; angryBirdLarge(77, 31) <= 4; angryBirdLarge(77, 32) <= 4; angryBirdLarge(77, 33) <= 4; angryBirdLarge(77, 34) <= 4; angryBirdLarge(77, 35) <= 4; angryBirdLarge(77, 36) <= 4; angryBirdLarge(77, 37) <= 4; angryBirdLarge(77, 38) <= 4; angryBirdLarge(77, 39) <= 4; angryBirdLarge(77, 40) <= 4; angryBirdLarge(77, 41) <= 4; angryBirdLarge(77, 42) <= 4; angryBirdLarge(77, 43) <= 4; angryBirdLarge(77, 44) <= 4; angryBirdLarge(77, 45) <= 4; angryBirdLarge(77, 46) <= 4; angryBirdLarge(77, 47) <= 4; angryBirdLarge(77, 48) <= 4; angryBirdLarge(77, 49) <= 4; angryBirdLarge(77, 50) <= 4; angryBirdLarge(77, 51) <= 4; angryBirdLarge(77, 52) <= 4; angryBirdLarge(77, 53) <= 4; angryBirdLarge(77, 54) <= 4; angryBirdLarge(77, 55) <= 4; angryBirdLarge(77, 56) <= 4; angryBirdLarge(77, 57) <= 4; angryBirdLarge(77, 58) <= 4; angryBirdLarge(77, 59) <= 4; angryBirdLarge(77, 60) <= 4; angryBirdLarge(77, 61) <= 4; angryBirdLarge(77, 62) <= 4; angryBirdLarge(77, 63) <= 4; angryBirdLarge(77, 64) <= 4; angryBirdLarge(77, 65) <= 4; angryBirdLarge(77, 66) <= 4; angryBirdLarge(77, 67) <= 4; angryBirdLarge(77, 68) <= 4; angryBirdLarge(77, 69) <= 4; angryBirdLarge(77, 70) <= 4; angryBirdLarge(77, 71) <= 4; angryBirdLarge(77, 72) <= 4; angryBirdLarge(77, 73) <= 4; angryBirdLarge(77, 74) <= 4; angryBirdLarge(77, 75) <= 4; angryBirdLarge(77, 76) <= 4; angryBirdLarge(77, 77) <= 4; angryBirdLarge(77, 78) <= 5; angryBirdLarge(77, 79) <= 5; angryBirdLarge(77, 80) <= 5; angryBirdLarge(77, 81) <= 5; angryBirdLarge(77, 82) <= 5; angryBirdLarge(77, 83) <= 5; angryBirdLarge(77, 84) <= 2; angryBirdLarge(77, 85) <= 2; angryBirdLarge(77, 86) <= 2; angryBirdLarge(77, 87) <= 2; angryBirdLarge(77, 88) <= 2; angryBirdLarge(77, 89) <= 2; angryBirdLarge(77, 90) <= 2; angryBirdLarge(77, 91) <= 2; angryBirdLarge(77, 92) <= 2; angryBirdLarge(77, 93) <= 2; angryBirdLarge(77, 94) <= 2; angryBirdLarge(77, 95) <= 2; angryBirdLarge(77, 96) <= 5; angryBirdLarge(77, 97) <= 5; angryBirdLarge(77, 98) <= 5; angryBirdLarge(77, 99) <= 5; angryBirdLarge(77, 100) <= 5; angryBirdLarge(77, 101) <= 5; angryBirdLarge(77, 102) <= 5; angryBirdLarge(77, 103) <= 5; angryBirdLarge(77, 104) <= 5; angryBirdLarge(77, 105) <= 5; angryBirdLarge(77, 106) <= 5; angryBirdLarge(77, 107) <= 5; angryBirdLarge(77, 108) <= 5; angryBirdLarge(77, 109) <= 5; angryBirdLarge(77, 110) <= 5; angryBirdLarge(77, 111) <= 5; angryBirdLarge(77, 112) <= 5; angryBirdLarge(77, 113) <= 5; angryBirdLarge(77, 114) <= 5; angryBirdLarge(77, 115) <= 5; angryBirdLarge(77, 116) <= 5; angryBirdLarge(77, 117) <= 5; angryBirdLarge(77, 118) <= 5; angryBirdLarge(77, 119) <= 5; angryBirdLarge(77, 120) <= 5; angryBirdLarge(77, 121) <= 5; angryBirdLarge(77, 122) <= 5; angryBirdLarge(77, 123) <= 5; angryBirdLarge(77, 124) <= 5; angryBirdLarge(77, 125) <= 5; angryBirdLarge(77, 126) <= 5; angryBirdLarge(77, 127) <= 5; angryBirdLarge(77, 128) <= 5; angryBirdLarge(77, 129) <= 5; angryBirdLarge(77, 130) <= 5; angryBirdLarge(77, 131) <= 5; angryBirdLarge(77, 132) <= 5; angryBirdLarge(77, 133) <= 5; angryBirdLarge(77, 134) <= 5; angryBirdLarge(77, 135) <= 5; angryBirdLarge(77, 136) <= 5; angryBirdLarge(77, 137) <= 5; angryBirdLarge(77, 138) <= 4; angryBirdLarge(77, 139) <= 4; angryBirdLarge(77, 140) <= 4; angryBirdLarge(77, 141) <= 4; angryBirdLarge(77, 142) <= 4; angryBirdLarge(77, 143) <= 4; angryBirdLarge(77, 144) <= 5; angryBirdLarge(77, 145) <= 5; angryBirdLarge(77, 146) <= 5; angryBirdLarge(77, 147) <= 5; angryBirdLarge(77, 148) <= 5; angryBirdLarge(77, 149) <= 5; 
angryBirdLarge(78, 0) <= 0; angryBirdLarge(78, 1) <= 0; angryBirdLarge(78, 2) <= 0; angryBirdLarge(78, 3) <= 0; angryBirdLarge(78, 4) <= 0; angryBirdLarge(78, 5) <= 0; angryBirdLarge(78, 6) <= 5; angryBirdLarge(78, 7) <= 5; angryBirdLarge(78, 8) <= 5; angryBirdLarge(78, 9) <= 5; angryBirdLarge(78, 10) <= 5; angryBirdLarge(78, 11) <= 5; angryBirdLarge(78, 12) <= 5; angryBirdLarge(78, 13) <= 5; angryBirdLarge(78, 14) <= 5; angryBirdLarge(78, 15) <= 5; angryBirdLarge(78, 16) <= 5; angryBirdLarge(78, 17) <= 5; angryBirdLarge(78, 18) <= 5; angryBirdLarge(78, 19) <= 5; angryBirdLarge(78, 20) <= 5; angryBirdLarge(78, 21) <= 5; angryBirdLarge(78, 22) <= 5; angryBirdLarge(78, 23) <= 5; angryBirdLarge(78, 24) <= 5; angryBirdLarge(78, 25) <= 5; angryBirdLarge(78, 26) <= 5; angryBirdLarge(78, 27) <= 5; angryBirdLarge(78, 28) <= 5; angryBirdLarge(78, 29) <= 5; angryBirdLarge(78, 30) <= 4; angryBirdLarge(78, 31) <= 4; angryBirdLarge(78, 32) <= 4; angryBirdLarge(78, 33) <= 4; angryBirdLarge(78, 34) <= 4; angryBirdLarge(78, 35) <= 4; angryBirdLarge(78, 36) <= 4; angryBirdLarge(78, 37) <= 4; angryBirdLarge(78, 38) <= 4; angryBirdLarge(78, 39) <= 4; angryBirdLarge(78, 40) <= 4; angryBirdLarge(78, 41) <= 4; angryBirdLarge(78, 42) <= 4; angryBirdLarge(78, 43) <= 4; angryBirdLarge(78, 44) <= 4; angryBirdLarge(78, 45) <= 4; angryBirdLarge(78, 46) <= 4; angryBirdLarge(78, 47) <= 4; angryBirdLarge(78, 48) <= 4; angryBirdLarge(78, 49) <= 4; angryBirdLarge(78, 50) <= 4; angryBirdLarge(78, 51) <= 4; angryBirdLarge(78, 52) <= 4; angryBirdLarge(78, 53) <= 4; angryBirdLarge(78, 54) <= 4; angryBirdLarge(78, 55) <= 4; angryBirdLarge(78, 56) <= 4; angryBirdLarge(78, 57) <= 4; angryBirdLarge(78, 58) <= 4; angryBirdLarge(78, 59) <= 4; angryBirdLarge(78, 60) <= 4; angryBirdLarge(78, 61) <= 4; angryBirdLarge(78, 62) <= 4; angryBirdLarge(78, 63) <= 4; angryBirdLarge(78, 64) <= 4; angryBirdLarge(78, 65) <= 4; angryBirdLarge(78, 66) <= 4; angryBirdLarge(78, 67) <= 4; angryBirdLarge(78, 68) <= 4; angryBirdLarge(78, 69) <= 4; angryBirdLarge(78, 70) <= 4; angryBirdLarge(78, 71) <= 4; angryBirdLarge(78, 72) <= 4; angryBirdLarge(78, 73) <= 4; angryBirdLarge(78, 74) <= 4; angryBirdLarge(78, 75) <= 4; angryBirdLarge(78, 76) <= 4; angryBirdLarge(78, 77) <= 4; angryBirdLarge(78, 78) <= 5; angryBirdLarge(78, 79) <= 5; angryBirdLarge(78, 80) <= 5; angryBirdLarge(78, 81) <= 5; angryBirdLarge(78, 82) <= 5; angryBirdLarge(78, 83) <= 5; angryBirdLarge(78, 84) <= 2; angryBirdLarge(78, 85) <= 2; angryBirdLarge(78, 86) <= 2; angryBirdLarge(78, 87) <= 2; angryBirdLarge(78, 88) <= 2; angryBirdLarge(78, 89) <= 2; angryBirdLarge(78, 90) <= 2; angryBirdLarge(78, 91) <= 2; angryBirdLarge(78, 92) <= 2; angryBirdLarge(78, 93) <= 2; angryBirdLarge(78, 94) <= 2; angryBirdLarge(78, 95) <= 2; angryBirdLarge(78, 96) <= 2; angryBirdLarge(78, 97) <= 2; angryBirdLarge(78, 98) <= 2; angryBirdLarge(78, 99) <= 2; angryBirdLarge(78, 100) <= 2; angryBirdLarge(78, 101) <= 2; angryBirdLarge(78, 102) <= 5; angryBirdLarge(78, 103) <= 5; angryBirdLarge(78, 104) <= 5; angryBirdLarge(78, 105) <= 5; angryBirdLarge(78, 106) <= 5; angryBirdLarge(78, 107) <= 5; angryBirdLarge(78, 108) <= 2; angryBirdLarge(78, 109) <= 2; angryBirdLarge(78, 110) <= 2; angryBirdLarge(78, 111) <= 2; angryBirdLarge(78, 112) <= 2; angryBirdLarge(78, 113) <= 2; angryBirdLarge(78, 114) <= 2; angryBirdLarge(78, 115) <= 2; angryBirdLarge(78, 116) <= 2; angryBirdLarge(78, 117) <= 2; angryBirdLarge(78, 118) <= 2; angryBirdLarge(78, 119) <= 2; angryBirdLarge(78, 120) <= 5; angryBirdLarge(78, 121) <= 5; angryBirdLarge(78, 122) <= 5; angryBirdLarge(78, 123) <= 5; angryBirdLarge(78, 124) <= 5; angryBirdLarge(78, 125) <= 5; angryBirdLarge(78, 126) <= 2; angryBirdLarge(78, 127) <= 2; angryBirdLarge(78, 128) <= 2; angryBirdLarge(78, 129) <= 2; angryBirdLarge(78, 130) <= 2; angryBirdLarge(78, 131) <= 2; angryBirdLarge(78, 132) <= 5; angryBirdLarge(78, 133) <= 5; angryBirdLarge(78, 134) <= 5; angryBirdLarge(78, 135) <= 5; angryBirdLarge(78, 136) <= 5; angryBirdLarge(78, 137) <= 5; angryBirdLarge(78, 138) <= 4; angryBirdLarge(78, 139) <= 4; angryBirdLarge(78, 140) <= 4; angryBirdLarge(78, 141) <= 4; angryBirdLarge(78, 142) <= 4; angryBirdLarge(78, 143) <= 4; angryBirdLarge(78, 144) <= 5; angryBirdLarge(78, 145) <= 5; angryBirdLarge(78, 146) <= 5; angryBirdLarge(78, 147) <= 5; angryBirdLarge(78, 148) <= 5; angryBirdLarge(78, 149) <= 5; 
angryBirdLarge(79, 0) <= 0; angryBirdLarge(79, 1) <= 0; angryBirdLarge(79, 2) <= 0; angryBirdLarge(79, 3) <= 0; angryBirdLarge(79, 4) <= 0; angryBirdLarge(79, 5) <= 0; angryBirdLarge(79, 6) <= 5; angryBirdLarge(79, 7) <= 5; angryBirdLarge(79, 8) <= 5; angryBirdLarge(79, 9) <= 5; angryBirdLarge(79, 10) <= 5; angryBirdLarge(79, 11) <= 5; angryBirdLarge(79, 12) <= 5; angryBirdLarge(79, 13) <= 5; angryBirdLarge(79, 14) <= 5; angryBirdLarge(79, 15) <= 5; angryBirdLarge(79, 16) <= 5; angryBirdLarge(79, 17) <= 5; angryBirdLarge(79, 18) <= 5; angryBirdLarge(79, 19) <= 5; angryBirdLarge(79, 20) <= 5; angryBirdLarge(79, 21) <= 5; angryBirdLarge(79, 22) <= 5; angryBirdLarge(79, 23) <= 5; angryBirdLarge(79, 24) <= 5; angryBirdLarge(79, 25) <= 5; angryBirdLarge(79, 26) <= 5; angryBirdLarge(79, 27) <= 5; angryBirdLarge(79, 28) <= 5; angryBirdLarge(79, 29) <= 5; angryBirdLarge(79, 30) <= 4; angryBirdLarge(79, 31) <= 4; angryBirdLarge(79, 32) <= 4; angryBirdLarge(79, 33) <= 4; angryBirdLarge(79, 34) <= 4; angryBirdLarge(79, 35) <= 4; angryBirdLarge(79, 36) <= 4; angryBirdLarge(79, 37) <= 4; angryBirdLarge(79, 38) <= 4; angryBirdLarge(79, 39) <= 4; angryBirdLarge(79, 40) <= 4; angryBirdLarge(79, 41) <= 4; angryBirdLarge(79, 42) <= 4; angryBirdLarge(79, 43) <= 4; angryBirdLarge(79, 44) <= 4; angryBirdLarge(79, 45) <= 4; angryBirdLarge(79, 46) <= 4; angryBirdLarge(79, 47) <= 4; angryBirdLarge(79, 48) <= 4; angryBirdLarge(79, 49) <= 4; angryBirdLarge(79, 50) <= 4; angryBirdLarge(79, 51) <= 4; angryBirdLarge(79, 52) <= 4; angryBirdLarge(79, 53) <= 4; angryBirdLarge(79, 54) <= 4; angryBirdLarge(79, 55) <= 4; angryBirdLarge(79, 56) <= 4; angryBirdLarge(79, 57) <= 4; angryBirdLarge(79, 58) <= 4; angryBirdLarge(79, 59) <= 4; angryBirdLarge(79, 60) <= 4; angryBirdLarge(79, 61) <= 4; angryBirdLarge(79, 62) <= 4; angryBirdLarge(79, 63) <= 4; angryBirdLarge(79, 64) <= 4; angryBirdLarge(79, 65) <= 4; angryBirdLarge(79, 66) <= 4; angryBirdLarge(79, 67) <= 4; angryBirdLarge(79, 68) <= 4; angryBirdLarge(79, 69) <= 4; angryBirdLarge(79, 70) <= 4; angryBirdLarge(79, 71) <= 4; angryBirdLarge(79, 72) <= 4; angryBirdLarge(79, 73) <= 4; angryBirdLarge(79, 74) <= 4; angryBirdLarge(79, 75) <= 4; angryBirdLarge(79, 76) <= 4; angryBirdLarge(79, 77) <= 4; angryBirdLarge(79, 78) <= 5; angryBirdLarge(79, 79) <= 5; angryBirdLarge(79, 80) <= 5; angryBirdLarge(79, 81) <= 5; angryBirdLarge(79, 82) <= 5; angryBirdLarge(79, 83) <= 5; angryBirdLarge(79, 84) <= 2; angryBirdLarge(79, 85) <= 2; angryBirdLarge(79, 86) <= 2; angryBirdLarge(79, 87) <= 2; angryBirdLarge(79, 88) <= 2; angryBirdLarge(79, 89) <= 2; angryBirdLarge(79, 90) <= 2; angryBirdLarge(79, 91) <= 2; angryBirdLarge(79, 92) <= 2; angryBirdLarge(79, 93) <= 2; angryBirdLarge(79, 94) <= 2; angryBirdLarge(79, 95) <= 2; angryBirdLarge(79, 96) <= 2; angryBirdLarge(79, 97) <= 2; angryBirdLarge(79, 98) <= 2; angryBirdLarge(79, 99) <= 2; angryBirdLarge(79, 100) <= 2; angryBirdLarge(79, 101) <= 2; angryBirdLarge(79, 102) <= 5; angryBirdLarge(79, 103) <= 5; angryBirdLarge(79, 104) <= 5; angryBirdLarge(79, 105) <= 5; angryBirdLarge(79, 106) <= 5; angryBirdLarge(79, 107) <= 5; angryBirdLarge(79, 108) <= 2; angryBirdLarge(79, 109) <= 2; angryBirdLarge(79, 110) <= 2; angryBirdLarge(79, 111) <= 2; angryBirdLarge(79, 112) <= 2; angryBirdLarge(79, 113) <= 2; angryBirdLarge(79, 114) <= 2; angryBirdLarge(79, 115) <= 2; angryBirdLarge(79, 116) <= 2; angryBirdLarge(79, 117) <= 2; angryBirdLarge(79, 118) <= 2; angryBirdLarge(79, 119) <= 2; angryBirdLarge(79, 120) <= 5; angryBirdLarge(79, 121) <= 5; angryBirdLarge(79, 122) <= 5; angryBirdLarge(79, 123) <= 5; angryBirdLarge(79, 124) <= 5; angryBirdLarge(79, 125) <= 5; angryBirdLarge(79, 126) <= 2; angryBirdLarge(79, 127) <= 2; angryBirdLarge(79, 128) <= 2; angryBirdLarge(79, 129) <= 2; angryBirdLarge(79, 130) <= 2; angryBirdLarge(79, 131) <= 2; angryBirdLarge(79, 132) <= 5; angryBirdLarge(79, 133) <= 5; angryBirdLarge(79, 134) <= 5; angryBirdLarge(79, 135) <= 5; angryBirdLarge(79, 136) <= 5; angryBirdLarge(79, 137) <= 5; angryBirdLarge(79, 138) <= 4; angryBirdLarge(79, 139) <= 4; angryBirdLarge(79, 140) <= 4; angryBirdLarge(79, 141) <= 4; angryBirdLarge(79, 142) <= 4; angryBirdLarge(79, 143) <= 4; angryBirdLarge(79, 144) <= 5; angryBirdLarge(79, 145) <= 5; angryBirdLarge(79, 146) <= 5; angryBirdLarge(79, 147) <= 5; angryBirdLarge(79, 148) <= 5; angryBirdLarge(79, 149) <= 5; 
angryBirdLarge(80, 0) <= 0; angryBirdLarge(80, 1) <= 0; angryBirdLarge(80, 2) <= 0; angryBirdLarge(80, 3) <= 0; angryBirdLarge(80, 4) <= 0; angryBirdLarge(80, 5) <= 0; angryBirdLarge(80, 6) <= 5; angryBirdLarge(80, 7) <= 5; angryBirdLarge(80, 8) <= 5; angryBirdLarge(80, 9) <= 5; angryBirdLarge(80, 10) <= 5; angryBirdLarge(80, 11) <= 5; angryBirdLarge(80, 12) <= 5; angryBirdLarge(80, 13) <= 5; angryBirdLarge(80, 14) <= 5; angryBirdLarge(80, 15) <= 5; angryBirdLarge(80, 16) <= 5; angryBirdLarge(80, 17) <= 5; angryBirdLarge(80, 18) <= 5; angryBirdLarge(80, 19) <= 5; angryBirdLarge(80, 20) <= 5; angryBirdLarge(80, 21) <= 5; angryBirdLarge(80, 22) <= 5; angryBirdLarge(80, 23) <= 5; angryBirdLarge(80, 24) <= 5; angryBirdLarge(80, 25) <= 5; angryBirdLarge(80, 26) <= 5; angryBirdLarge(80, 27) <= 5; angryBirdLarge(80, 28) <= 5; angryBirdLarge(80, 29) <= 5; angryBirdLarge(80, 30) <= 4; angryBirdLarge(80, 31) <= 4; angryBirdLarge(80, 32) <= 4; angryBirdLarge(80, 33) <= 4; angryBirdLarge(80, 34) <= 4; angryBirdLarge(80, 35) <= 4; angryBirdLarge(80, 36) <= 4; angryBirdLarge(80, 37) <= 4; angryBirdLarge(80, 38) <= 4; angryBirdLarge(80, 39) <= 4; angryBirdLarge(80, 40) <= 4; angryBirdLarge(80, 41) <= 4; angryBirdLarge(80, 42) <= 4; angryBirdLarge(80, 43) <= 4; angryBirdLarge(80, 44) <= 4; angryBirdLarge(80, 45) <= 4; angryBirdLarge(80, 46) <= 4; angryBirdLarge(80, 47) <= 4; angryBirdLarge(80, 48) <= 4; angryBirdLarge(80, 49) <= 4; angryBirdLarge(80, 50) <= 4; angryBirdLarge(80, 51) <= 4; angryBirdLarge(80, 52) <= 4; angryBirdLarge(80, 53) <= 4; angryBirdLarge(80, 54) <= 4; angryBirdLarge(80, 55) <= 4; angryBirdLarge(80, 56) <= 4; angryBirdLarge(80, 57) <= 4; angryBirdLarge(80, 58) <= 4; angryBirdLarge(80, 59) <= 4; angryBirdLarge(80, 60) <= 4; angryBirdLarge(80, 61) <= 4; angryBirdLarge(80, 62) <= 4; angryBirdLarge(80, 63) <= 4; angryBirdLarge(80, 64) <= 4; angryBirdLarge(80, 65) <= 4; angryBirdLarge(80, 66) <= 4; angryBirdLarge(80, 67) <= 4; angryBirdLarge(80, 68) <= 4; angryBirdLarge(80, 69) <= 4; angryBirdLarge(80, 70) <= 4; angryBirdLarge(80, 71) <= 4; angryBirdLarge(80, 72) <= 4; angryBirdLarge(80, 73) <= 4; angryBirdLarge(80, 74) <= 4; angryBirdLarge(80, 75) <= 4; angryBirdLarge(80, 76) <= 4; angryBirdLarge(80, 77) <= 4; angryBirdLarge(80, 78) <= 5; angryBirdLarge(80, 79) <= 5; angryBirdLarge(80, 80) <= 5; angryBirdLarge(80, 81) <= 5; angryBirdLarge(80, 82) <= 5; angryBirdLarge(80, 83) <= 5; angryBirdLarge(80, 84) <= 2; angryBirdLarge(80, 85) <= 2; angryBirdLarge(80, 86) <= 2; angryBirdLarge(80, 87) <= 2; angryBirdLarge(80, 88) <= 2; angryBirdLarge(80, 89) <= 2; angryBirdLarge(80, 90) <= 2; angryBirdLarge(80, 91) <= 2; angryBirdLarge(80, 92) <= 2; angryBirdLarge(80, 93) <= 2; angryBirdLarge(80, 94) <= 2; angryBirdLarge(80, 95) <= 2; angryBirdLarge(80, 96) <= 2; angryBirdLarge(80, 97) <= 2; angryBirdLarge(80, 98) <= 2; angryBirdLarge(80, 99) <= 2; angryBirdLarge(80, 100) <= 2; angryBirdLarge(80, 101) <= 2; angryBirdLarge(80, 102) <= 5; angryBirdLarge(80, 103) <= 5; angryBirdLarge(80, 104) <= 5; angryBirdLarge(80, 105) <= 5; angryBirdLarge(80, 106) <= 5; angryBirdLarge(80, 107) <= 5; angryBirdLarge(80, 108) <= 2; angryBirdLarge(80, 109) <= 2; angryBirdLarge(80, 110) <= 2; angryBirdLarge(80, 111) <= 2; angryBirdLarge(80, 112) <= 2; angryBirdLarge(80, 113) <= 2; angryBirdLarge(80, 114) <= 2; angryBirdLarge(80, 115) <= 2; angryBirdLarge(80, 116) <= 2; angryBirdLarge(80, 117) <= 2; angryBirdLarge(80, 118) <= 2; angryBirdLarge(80, 119) <= 2; angryBirdLarge(80, 120) <= 5; angryBirdLarge(80, 121) <= 5; angryBirdLarge(80, 122) <= 5; angryBirdLarge(80, 123) <= 5; angryBirdLarge(80, 124) <= 5; angryBirdLarge(80, 125) <= 5; angryBirdLarge(80, 126) <= 2; angryBirdLarge(80, 127) <= 2; angryBirdLarge(80, 128) <= 2; angryBirdLarge(80, 129) <= 2; angryBirdLarge(80, 130) <= 2; angryBirdLarge(80, 131) <= 2; angryBirdLarge(80, 132) <= 5; angryBirdLarge(80, 133) <= 5; angryBirdLarge(80, 134) <= 5; angryBirdLarge(80, 135) <= 5; angryBirdLarge(80, 136) <= 5; angryBirdLarge(80, 137) <= 5; angryBirdLarge(80, 138) <= 4; angryBirdLarge(80, 139) <= 4; angryBirdLarge(80, 140) <= 4; angryBirdLarge(80, 141) <= 4; angryBirdLarge(80, 142) <= 4; angryBirdLarge(80, 143) <= 4; angryBirdLarge(80, 144) <= 5; angryBirdLarge(80, 145) <= 5; angryBirdLarge(80, 146) <= 5; angryBirdLarge(80, 147) <= 5; angryBirdLarge(80, 148) <= 5; angryBirdLarge(80, 149) <= 5; 
angryBirdLarge(81, 0) <= 0; angryBirdLarge(81, 1) <= 0; angryBirdLarge(81, 2) <= 0; angryBirdLarge(81, 3) <= 0; angryBirdLarge(81, 4) <= 0; angryBirdLarge(81, 5) <= 0; angryBirdLarge(81, 6) <= 5; angryBirdLarge(81, 7) <= 5; angryBirdLarge(81, 8) <= 5; angryBirdLarge(81, 9) <= 5; angryBirdLarge(81, 10) <= 5; angryBirdLarge(81, 11) <= 5; angryBirdLarge(81, 12) <= 5; angryBirdLarge(81, 13) <= 5; angryBirdLarge(81, 14) <= 5; angryBirdLarge(81, 15) <= 5; angryBirdLarge(81, 16) <= 5; angryBirdLarge(81, 17) <= 5; angryBirdLarge(81, 18) <= 5; angryBirdLarge(81, 19) <= 5; angryBirdLarge(81, 20) <= 5; angryBirdLarge(81, 21) <= 5; angryBirdLarge(81, 22) <= 5; angryBirdLarge(81, 23) <= 5; angryBirdLarge(81, 24) <= 5; angryBirdLarge(81, 25) <= 5; angryBirdLarge(81, 26) <= 5; angryBirdLarge(81, 27) <= 5; angryBirdLarge(81, 28) <= 5; angryBirdLarge(81, 29) <= 5; angryBirdLarge(81, 30) <= 4; angryBirdLarge(81, 31) <= 4; angryBirdLarge(81, 32) <= 4; angryBirdLarge(81, 33) <= 4; angryBirdLarge(81, 34) <= 4; angryBirdLarge(81, 35) <= 4; angryBirdLarge(81, 36) <= 4; angryBirdLarge(81, 37) <= 4; angryBirdLarge(81, 38) <= 4; angryBirdLarge(81, 39) <= 4; angryBirdLarge(81, 40) <= 4; angryBirdLarge(81, 41) <= 4; angryBirdLarge(81, 42) <= 4; angryBirdLarge(81, 43) <= 4; angryBirdLarge(81, 44) <= 4; angryBirdLarge(81, 45) <= 4; angryBirdLarge(81, 46) <= 4; angryBirdLarge(81, 47) <= 4; angryBirdLarge(81, 48) <= 4; angryBirdLarge(81, 49) <= 4; angryBirdLarge(81, 50) <= 4; angryBirdLarge(81, 51) <= 4; angryBirdLarge(81, 52) <= 4; angryBirdLarge(81, 53) <= 4; angryBirdLarge(81, 54) <= 4; angryBirdLarge(81, 55) <= 4; angryBirdLarge(81, 56) <= 4; angryBirdLarge(81, 57) <= 4; angryBirdLarge(81, 58) <= 4; angryBirdLarge(81, 59) <= 4; angryBirdLarge(81, 60) <= 4; angryBirdLarge(81, 61) <= 4; angryBirdLarge(81, 62) <= 4; angryBirdLarge(81, 63) <= 4; angryBirdLarge(81, 64) <= 4; angryBirdLarge(81, 65) <= 4; angryBirdLarge(81, 66) <= 4; angryBirdLarge(81, 67) <= 4; angryBirdLarge(81, 68) <= 4; angryBirdLarge(81, 69) <= 4; angryBirdLarge(81, 70) <= 4; angryBirdLarge(81, 71) <= 4; angryBirdLarge(81, 72) <= 4; angryBirdLarge(81, 73) <= 4; angryBirdLarge(81, 74) <= 4; angryBirdLarge(81, 75) <= 4; angryBirdLarge(81, 76) <= 4; angryBirdLarge(81, 77) <= 4; angryBirdLarge(81, 78) <= 5; angryBirdLarge(81, 79) <= 5; angryBirdLarge(81, 80) <= 5; angryBirdLarge(81, 81) <= 5; angryBirdLarge(81, 82) <= 5; angryBirdLarge(81, 83) <= 5; angryBirdLarge(81, 84) <= 2; angryBirdLarge(81, 85) <= 2; angryBirdLarge(81, 86) <= 2; angryBirdLarge(81, 87) <= 2; angryBirdLarge(81, 88) <= 2; angryBirdLarge(81, 89) <= 2; angryBirdLarge(81, 90) <= 2; angryBirdLarge(81, 91) <= 2; angryBirdLarge(81, 92) <= 2; angryBirdLarge(81, 93) <= 2; angryBirdLarge(81, 94) <= 2; angryBirdLarge(81, 95) <= 2; angryBirdLarge(81, 96) <= 2; angryBirdLarge(81, 97) <= 2; angryBirdLarge(81, 98) <= 2; angryBirdLarge(81, 99) <= 2; angryBirdLarge(81, 100) <= 2; angryBirdLarge(81, 101) <= 2; angryBirdLarge(81, 102) <= 5; angryBirdLarge(81, 103) <= 5; angryBirdLarge(81, 104) <= 5; angryBirdLarge(81, 105) <= 5; angryBirdLarge(81, 106) <= 5; angryBirdLarge(81, 107) <= 5; angryBirdLarge(81, 108) <= 2; angryBirdLarge(81, 109) <= 2; angryBirdLarge(81, 110) <= 2; angryBirdLarge(81, 111) <= 2; angryBirdLarge(81, 112) <= 2; angryBirdLarge(81, 113) <= 2; angryBirdLarge(81, 114) <= 2; angryBirdLarge(81, 115) <= 2; angryBirdLarge(81, 116) <= 2; angryBirdLarge(81, 117) <= 2; angryBirdLarge(81, 118) <= 2; angryBirdLarge(81, 119) <= 2; angryBirdLarge(81, 120) <= 5; angryBirdLarge(81, 121) <= 5; angryBirdLarge(81, 122) <= 5; angryBirdLarge(81, 123) <= 5; angryBirdLarge(81, 124) <= 5; angryBirdLarge(81, 125) <= 5; angryBirdLarge(81, 126) <= 2; angryBirdLarge(81, 127) <= 2; angryBirdLarge(81, 128) <= 2; angryBirdLarge(81, 129) <= 2; angryBirdLarge(81, 130) <= 2; angryBirdLarge(81, 131) <= 2; angryBirdLarge(81, 132) <= 5; angryBirdLarge(81, 133) <= 5; angryBirdLarge(81, 134) <= 5; angryBirdLarge(81, 135) <= 5; angryBirdLarge(81, 136) <= 5; angryBirdLarge(81, 137) <= 5; angryBirdLarge(81, 138) <= 4; angryBirdLarge(81, 139) <= 4; angryBirdLarge(81, 140) <= 4; angryBirdLarge(81, 141) <= 4; angryBirdLarge(81, 142) <= 4; angryBirdLarge(81, 143) <= 4; angryBirdLarge(81, 144) <= 5; angryBirdLarge(81, 145) <= 5; angryBirdLarge(81, 146) <= 5; angryBirdLarge(81, 147) <= 5; angryBirdLarge(81, 148) <= 5; angryBirdLarge(81, 149) <= 5; 
angryBirdLarge(82, 0) <= 0; angryBirdLarge(82, 1) <= 0; angryBirdLarge(82, 2) <= 0; angryBirdLarge(82, 3) <= 0; angryBirdLarge(82, 4) <= 0; angryBirdLarge(82, 5) <= 0; angryBirdLarge(82, 6) <= 5; angryBirdLarge(82, 7) <= 5; angryBirdLarge(82, 8) <= 5; angryBirdLarge(82, 9) <= 5; angryBirdLarge(82, 10) <= 5; angryBirdLarge(82, 11) <= 5; angryBirdLarge(82, 12) <= 5; angryBirdLarge(82, 13) <= 5; angryBirdLarge(82, 14) <= 5; angryBirdLarge(82, 15) <= 5; angryBirdLarge(82, 16) <= 5; angryBirdLarge(82, 17) <= 5; angryBirdLarge(82, 18) <= 5; angryBirdLarge(82, 19) <= 5; angryBirdLarge(82, 20) <= 5; angryBirdLarge(82, 21) <= 5; angryBirdLarge(82, 22) <= 5; angryBirdLarge(82, 23) <= 5; angryBirdLarge(82, 24) <= 5; angryBirdLarge(82, 25) <= 5; angryBirdLarge(82, 26) <= 5; angryBirdLarge(82, 27) <= 5; angryBirdLarge(82, 28) <= 5; angryBirdLarge(82, 29) <= 5; angryBirdLarge(82, 30) <= 4; angryBirdLarge(82, 31) <= 4; angryBirdLarge(82, 32) <= 4; angryBirdLarge(82, 33) <= 4; angryBirdLarge(82, 34) <= 4; angryBirdLarge(82, 35) <= 4; angryBirdLarge(82, 36) <= 4; angryBirdLarge(82, 37) <= 4; angryBirdLarge(82, 38) <= 4; angryBirdLarge(82, 39) <= 4; angryBirdLarge(82, 40) <= 4; angryBirdLarge(82, 41) <= 4; angryBirdLarge(82, 42) <= 4; angryBirdLarge(82, 43) <= 4; angryBirdLarge(82, 44) <= 4; angryBirdLarge(82, 45) <= 4; angryBirdLarge(82, 46) <= 4; angryBirdLarge(82, 47) <= 4; angryBirdLarge(82, 48) <= 4; angryBirdLarge(82, 49) <= 4; angryBirdLarge(82, 50) <= 4; angryBirdLarge(82, 51) <= 4; angryBirdLarge(82, 52) <= 4; angryBirdLarge(82, 53) <= 4; angryBirdLarge(82, 54) <= 4; angryBirdLarge(82, 55) <= 4; angryBirdLarge(82, 56) <= 4; angryBirdLarge(82, 57) <= 4; angryBirdLarge(82, 58) <= 4; angryBirdLarge(82, 59) <= 4; angryBirdLarge(82, 60) <= 4; angryBirdLarge(82, 61) <= 4; angryBirdLarge(82, 62) <= 4; angryBirdLarge(82, 63) <= 4; angryBirdLarge(82, 64) <= 4; angryBirdLarge(82, 65) <= 4; angryBirdLarge(82, 66) <= 4; angryBirdLarge(82, 67) <= 4; angryBirdLarge(82, 68) <= 4; angryBirdLarge(82, 69) <= 4; angryBirdLarge(82, 70) <= 4; angryBirdLarge(82, 71) <= 4; angryBirdLarge(82, 72) <= 4; angryBirdLarge(82, 73) <= 4; angryBirdLarge(82, 74) <= 4; angryBirdLarge(82, 75) <= 4; angryBirdLarge(82, 76) <= 4; angryBirdLarge(82, 77) <= 4; angryBirdLarge(82, 78) <= 5; angryBirdLarge(82, 79) <= 5; angryBirdLarge(82, 80) <= 5; angryBirdLarge(82, 81) <= 5; angryBirdLarge(82, 82) <= 5; angryBirdLarge(82, 83) <= 5; angryBirdLarge(82, 84) <= 2; angryBirdLarge(82, 85) <= 2; angryBirdLarge(82, 86) <= 2; angryBirdLarge(82, 87) <= 2; angryBirdLarge(82, 88) <= 2; angryBirdLarge(82, 89) <= 2; angryBirdLarge(82, 90) <= 2; angryBirdLarge(82, 91) <= 2; angryBirdLarge(82, 92) <= 2; angryBirdLarge(82, 93) <= 2; angryBirdLarge(82, 94) <= 2; angryBirdLarge(82, 95) <= 2; angryBirdLarge(82, 96) <= 2; angryBirdLarge(82, 97) <= 2; angryBirdLarge(82, 98) <= 2; angryBirdLarge(82, 99) <= 2; angryBirdLarge(82, 100) <= 2; angryBirdLarge(82, 101) <= 2; angryBirdLarge(82, 102) <= 5; angryBirdLarge(82, 103) <= 5; angryBirdLarge(82, 104) <= 5; angryBirdLarge(82, 105) <= 5; angryBirdLarge(82, 106) <= 5; angryBirdLarge(82, 107) <= 5; angryBirdLarge(82, 108) <= 2; angryBirdLarge(82, 109) <= 2; angryBirdLarge(82, 110) <= 2; angryBirdLarge(82, 111) <= 2; angryBirdLarge(82, 112) <= 2; angryBirdLarge(82, 113) <= 2; angryBirdLarge(82, 114) <= 2; angryBirdLarge(82, 115) <= 2; angryBirdLarge(82, 116) <= 2; angryBirdLarge(82, 117) <= 2; angryBirdLarge(82, 118) <= 2; angryBirdLarge(82, 119) <= 2; angryBirdLarge(82, 120) <= 5; angryBirdLarge(82, 121) <= 5; angryBirdLarge(82, 122) <= 5; angryBirdLarge(82, 123) <= 5; angryBirdLarge(82, 124) <= 5; angryBirdLarge(82, 125) <= 5; angryBirdLarge(82, 126) <= 2; angryBirdLarge(82, 127) <= 2; angryBirdLarge(82, 128) <= 2; angryBirdLarge(82, 129) <= 2; angryBirdLarge(82, 130) <= 2; angryBirdLarge(82, 131) <= 2; angryBirdLarge(82, 132) <= 5; angryBirdLarge(82, 133) <= 5; angryBirdLarge(82, 134) <= 5; angryBirdLarge(82, 135) <= 5; angryBirdLarge(82, 136) <= 5; angryBirdLarge(82, 137) <= 5; angryBirdLarge(82, 138) <= 4; angryBirdLarge(82, 139) <= 4; angryBirdLarge(82, 140) <= 4; angryBirdLarge(82, 141) <= 4; angryBirdLarge(82, 142) <= 4; angryBirdLarge(82, 143) <= 4; angryBirdLarge(82, 144) <= 5; angryBirdLarge(82, 145) <= 5; angryBirdLarge(82, 146) <= 5; angryBirdLarge(82, 147) <= 5; angryBirdLarge(82, 148) <= 5; angryBirdLarge(82, 149) <= 5; 
angryBirdLarge(83, 0) <= 0; angryBirdLarge(83, 1) <= 0; angryBirdLarge(83, 2) <= 0; angryBirdLarge(83, 3) <= 0; angryBirdLarge(83, 4) <= 0; angryBirdLarge(83, 5) <= 0; angryBirdLarge(83, 6) <= 5; angryBirdLarge(83, 7) <= 5; angryBirdLarge(83, 8) <= 5; angryBirdLarge(83, 9) <= 5; angryBirdLarge(83, 10) <= 5; angryBirdLarge(83, 11) <= 5; angryBirdLarge(83, 12) <= 5; angryBirdLarge(83, 13) <= 5; angryBirdLarge(83, 14) <= 5; angryBirdLarge(83, 15) <= 5; angryBirdLarge(83, 16) <= 5; angryBirdLarge(83, 17) <= 5; angryBirdLarge(83, 18) <= 5; angryBirdLarge(83, 19) <= 5; angryBirdLarge(83, 20) <= 5; angryBirdLarge(83, 21) <= 5; angryBirdLarge(83, 22) <= 5; angryBirdLarge(83, 23) <= 5; angryBirdLarge(83, 24) <= 5; angryBirdLarge(83, 25) <= 5; angryBirdLarge(83, 26) <= 5; angryBirdLarge(83, 27) <= 5; angryBirdLarge(83, 28) <= 5; angryBirdLarge(83, 29) <= 5; angryBirdLarge(83, 30) <= 4; angryBirdLarge(83, 31) <= 4; angryBirdLarge(83, 32) <= 4; angryBirdLarge(83, 33) <= 4; angryBirdLarge(83, 34) <= 4; angryBirdLarge(83, 35) <= 4; angryBirdLarge(83, 36) <= 4; angryBirdLarge(83, 37) <= 4; angryBirdLarge(83, 38) <= 4; angryBirdLarge(83, 39) <= 4; angryBirdLarge(83, 40) <= 4; angryBirdLarge(83, 41) <= 4; angryBirdLarge(83, 42) <= 4; angryBirdLarge(83, 43) <= 4; angryBirdLarge(83, 44) <= 4; angryBirdLarge(83, 45) <= 4; angryBirdLarge(83, 46) <= 4; angryBirdLarge(83, 47) <= 4; angryBirdLarge(83, 48) <= 4; angryBirdLarge(83, 49) <= 4; angryBirdLarge(83, 50) <= 4; angryBirdLarge(83, 51) <= 4; angryBirdLarge(83, 52) <= 4; angryBirdLarge(83, 53) <= 4; angryBirdLarge(83, 54) <= 4; angryBirdLarge(83, 55) <= 4; angryBirdLarge(83, 56) <= 4; angryBirdLarge(83, 57) <= 4; angryBirdLarge(83, 58) <= 4; angryBirdLarge(83, 59) <= 4; angryBirdLarge(83, 60) <= 4; angryBirdLarge(83, 61) <= 4; angryBirdLarge(83, 62) <= 4; angryBirdLarge(83, 63) <= 4; angryBirdLarge(83, 64) <= 4; angryBirdLarge(83, 65) <= 4; angryBirdLarge(83, 66) <= 4; angryBirdLarge(83, 67) <= 4; angryBirdLarge(83, 68) <= 4; angryBirdLarge(83, 69) <= 4; angryBirdLarge(83, 70) <= 4; angryBirdLarge(83, 71) <= 4; angryBirdLarge(83, 72) <= 4; angryBirdLarge(83, 73) <= 4; angryBirdLarge(83, 74) <= 4; angryBirdLarge(83, 75) <= 4; angryBirdLarge(83, 76) <= 4; angryBirdLarge(83, 77) <= 4; angryBirdLarge(83, 78) <= 5; angryBirdLarge(83, 79) <= 5; angryBirdLarge(83, 80) <= 5; angryBirdLarge(83, 81) <= 5; angryBirdLarge(83, 82) <= 5; angryBirdLarge(83, 83) <= 5; angryBirdLarge(83, 84) <= 2; angryBirdLarge(83, 85) <= 2; angryBirdLarge(83, 86) <= 2; angryBirdLarge(83, 87) <= 2; angryBirdLarge(83, 88) <= 2; angryBirdLarge(83, 89) <= 2; angryBirdLarge(83, 90) <= 2; angryBirdLarge(83, 91) <= 2; angryBirdLarge(83, 92) <= 2; angryBirdLarge(83, 93) <= 2; angryBirdLarge(83, 94) <= 2; angryBirdLarge(83, 95) <= 2; angryBirdLarge(83, 96) <= 2; angryBirdLarge(83, 97) <= 2; angryBirdLarge(83, 98) <= 2; angryBirdLarge(83, 99) <= 2; angryBirdLarge(83, 100) <= 2; angryBirdLarge(83, 101) <= 2; angryBirdLarge(83, 102) <= 5; angryBirdLarge(83, 103) <= 5; angryBirdLarge(83, 104) <= 5; angryBirdLarge(83, 105) <= 5; angryBirdLarge(83, 106) <= 5; angryBirdLarge(83, 107) <= 5; angryBirdLarge(83, 108) <= 2; angryBirdLarge(83, 109) <= 2; angryBirdLarge(83, 110) <= 2; angryBirdLarge(83, 111) <= 2; angryBirdLarge(83, 112) <= 2; angryBirdLarge(83, 113) <= 2; angryBirdLarge(83, 114) <= 2; angryBirdLarge(83, 115) <= 2; angryBirdLarge(83, 116) <= 2; angryBirdLarge(83, 117) <= 2; angryBirdLarge(83, 118) <= 2; angryBirdLarge(83, 119) <= 2; angryBirdLarge(83, 120) <= 5; angryBirdLarge(83, 121) <= 5; angryBirdLarge(83, 122) <= 5; angryBirdLarge(83, 123) <= 5; angryBirdLarge(83, 124) <= 5; angryBirdLarge(83, 125) <= 5; angryBirdLarge(83, 126) <= 2; angryBirdLarge(83, 127) <= 2; angryBirdLarge(83, 128) <= 2; angryBirdLarge(83, 129) <= 2; angryBirdLarge(83, 130) <= 2; angryBirdLarge(83, 131) <= 2; angryBirdLarge(83, 132) <= 5; angryBirdLarge(83, 133) <= 5; angryBirdLarge(83, 134) <= 5; angryBirdLarge(83, 135) <= 5; angryBirdLarge(83, 136) <= 5; angryBirdLarge(83, 137) <= 5; angryBirdLarge(83, 138) <= 4; angryBirdLarge(83, 139) <= 4; angryBirdLarge(83, 140) <= 4; angryBirdLarge(83, 141) <= 4; angryBirdLarge(83, 142) <= 4; angryBirdLarge(83, 143) <= 4; angryBirdLarge(83, 144) <= 5; angryBirdLarge(83, 145) <= 5; angryBirdLarge(83, 146) <= 5; angryBirdLarge(83, 147) <= 5; angryBirdLarge(83, 148) <= 5; angryBirdLarge(83, 149) <= 5; 
angryBirdLarge(84, 0) <= 0; angryBirdLarge(84, 1) <= 0; angryBirdLarge(84, 2) <= 0; angryBirdLarge(84, 3) <= 0; angryBirdLarge(84, 4) <= 0; angryBirdLarge(84, 5) <= 0; angryBirdLarge(84, 6) <= 5; angryBirdLarge(84, 7) <= 5; angryBirdLarge(84, 8) <= 5; angryBirdLarge(84, 9) <= 5; angryBirdLarge(84, 10) <= 5; angryBirdLarge(84, 11) <= 5; angryBirdLarge(84, 12) <= 5; angryBirdLarge(84, 13) <= 5; angryBirdLarge(84, 14) <= 5; angryBirdLarge(84, 15) <= 5; angryBirdLarge(84, 16) <= 5; angryBirdLarge(84, 17) <= 5; angryBirdLarge(84, 18) <= 5; angryBirdLarge(84, 19) <= 5; angryBirdLarge(84, 20) <= 5; angryBirdLarge(84, 21) <= 5; angryBirdLarge(84, 22) <= 5; angryBirdLarge(84, 23) <= 5; angryBirdLarge(84, 24) <= 5; angryBirdLarge(84, 25) <= 5; angryBirdLarge(84, 26) <= 5; angryBirdLarge(84, 27) <= 5; angryBirdLarge(84, 28) <= 5; angryBirdLarge(84, 29) <= 5; angryBirdLarge(84, 30) <= 4; angryBirdLarge(84, 31) <= 4; angryBirdLarge(84, 32) <= 4; angryBirdLarge(84, 33) <= 4; angryBirdLarge(84, 34) <= 4; angryBirdLarge(84, 35) <= 4; angryBirdLarge(84, 36) <= 4; angryBirdLarge(84, 37) <= 4; angryBirdLarge(84, 38) <= 4; angryBirdLarge(84, 39) <= 4; angryBirdLarge(84, 40) <= 4; angryBirdLarge(84, 41) <= 4; angryBirdLarge(84, 42) <= 4; angryBirdLarge(84, 43) <= 4; angryBirdLarge(84, 44) <= 4; angryBirdLarge(84, 45) <= 4; angryBirdLarge(84, 46) <= 4; angryBirdLarge(84, 47) <= 4; angryBirdLarge(84, 48) <= 4; angryBirdLarge(84, 49) <= 4; angryBirdLarge(84, 50) <= 4; angryBirdLarge(84, 51) <= 4; angryBirdLarge(84, 52) <= 4; angryBirdLarge(84, 53) <= 4; angryBirdLarge(84, 54) <= 4; angryBirdLarge(84, 55) <= 4; angryBirdLarge(84, 56) <= 4; angryBirdLarge(84, 57) <= 4; angryBirdLarge(84, 58) <= 4; angryBirdLarge(84, 59) <= 4; angryBirdLarge(84, 60) <= 4; angryBirdLarge(84, 61) <= 4; angryBirdLarge(84, 62) <= 4; angryBirdLarge(84, 63) <= 4; angryBirdLarge(84, 64) <= 4; angryBirdLarge(84, 65) <= 4; angryBirdLarge(84, 66) <= 4; angryBirdLarge(84, 67) <= 4; angryBirdLarge(84, 68) <= 4; angryBirdLarge(84, 69) <= 4; angryBirdLarge(84, 70) <= 4; angryBirdLarge(84, 71) <= 4; angryBirdLarge(84, 72) <= 4; angryBirdLarge(84, 73) <= 4; angryBirdLarge(84, 74) <= 4; angryBirdLarge(84, 75) <= 4; angryBirdLarge(84, 76) <= 4; angryBirdLarge(84, 77) <= 4; angryBirdLarge(84, 78) <= 4; angryBirdLarge(84, 79) <= 4; angryBirdLarge(84, 80) <= 4; angryBirdLarge(84, 81) <= 4; angryBirdLarge(84, 82) <= 4; angryBirdLarge(84, 83) <= 4; angryBirdLarge(84, 84) <= 5; angryBirdLarge(84, 85) <= 5; angryBirdLarge(84, 86) <= 5; angryBirdLarge(84, 87) <= 5; angryBirdLarge(84, 88) <= 5; angryBirdLarge(84, 89) <= 5; angryBirdLarge(84, 90) <= 2; angryBirdLarge(84, 91) <= 2; angryBirdLarge(84, 92) <= 2; angryBirdLarge(84, 93) <= 2; angryBirdLarge(84, 94) <= 2; angryBirdLarge(84, 95) <= 2; angryBirdLarge(84, 96) <= 2; angryBirdLarge(84, 97) <= 2; angryBirdLarge(84, 98) <= 2; angryBirdLarge(84, 99) <= 2; angryBirdLarge(84, 100) <= 2; angryBirdLarge(84, 101) <= 2; angryBirdLarge(84, 102) <= 2; angryBirdLarge(84, 103) <= 2; angryBirdLarge(84, 104) <= 2; angryBirdLarge(84, 105) <= 2; angryBirdLarge(84, 106) <= 2; angryBirdLarge(84, 107) <= 2; angryBirdLarge(84, 108) <= 5; angryBirdLarge(84, 109) <= 5; angryBirdLarge(84, 110) <= 5; angryBirdLarge(84, 111) <= 5; angryBirdLarge(84, 112) <= 5; angryBirdLarge(84, 113) <= 5; angryBirdLarge(84, 114) <= 5; angryBirdLarge(84, 115) <= 5; angryBirdLarge(84, 116) <= 5; angryBirdLarge(84, 117) <= 5; angryBirdLarge(84, 118) <= 5; angryBirdLarge(84, 119) <= 5; angryBirdLarge(84, 120) <= 2; angryBirdLarge(84, 121) <= 2; angryBirdLarge(84, 122) <= 2; angryBirdLarge(84, 123) <= 2; angryBirdLarge(84, 124) <= 2; angryBirdLarge(84, 125) <= 2; angryBirdLarge(84, 126) <= 2; angryBirdLarge(84, 127) <= 2; angryBirdLarge(84, 128) <= 2; angryBirdLarge(84, 129) <= 2; angryBirdLarge(84, 130) <= 2; angryBirdLarge(84, 131) <= 2; angryBirdLarge(84, 132) <= 5; angryBirdLarge(84, 133) <= 5; angryBirdLarge(84, 134) <= 5; angryBirdLarge(84, 135) <= 5; angryBirdLarge(84, 136) <= 5; angryBirdLarge(84, 137) <= 5; angryBirdLarge(84, 138) <= 4; angryBirdLarge(84, 139) <= 4; angryBirdLarge(84, 140) <= 4; angryBirdLarge(84, 141) <= 4; angryBirdLarge(84, 142) <= 4; angryBirdLarge(84, 143) <= 4; angryBirdLarge(84, 144) <= 5; angryBirdLarge(84, 145) <= 5; angryBirdLarge(84, 146) <= 5; angryBirdLarge(84, 147) <= 5; angryBirdLarge(84, 148) <= 5; angryBirdLarge(84, 149) <= 5; 
angryBirdLarge(85, 0) <= 0; angryBirdLarge(85, 1) <= 0; angryBirdLarge(85, 2) <= 0; angryBirdLarge(85, 3) <= 0; angryBirdLarge(85, 4) <= 0; angryBirdLarge(85, 5) <= 0; angryBirdLarge(85, 6) <= 5; angryBirdLarge(85, 7) <= 5; angryBirdLarge(85, 8) <= 5; angryBirdLarge(85, 9) <= 5; angryBirdLarge(85, 10) <= 5; angryBirdLarge(85, 11) <= 5; angryBirdLarge(85, 12) <= 5; angryBirdLarge(85, 13) <= 5; angryBirdLarge(85, 14) <= 5; angryBirdLarge(85, 15) <= 5; angryBirdLarge(85, 16) <= 5; angryBirdLarge(85, 17) <= 5; angryBirdLarge(85, 18) <= 5; angryBirdLarge(85, 19) <= 5; angryBirdLarge(85, 20) <= 5; angryBirdLarge(85, 21) <= 5; angryBirdLarge(85, 22) <= 5; angryBirdLarge(85, 23) <= 5; angryBirdLarge(85, 24) <= 5; angryBirdLarge(85, 25) <= 5; angryBirdLarge(85, 26) <= 5; angryBirdLarge(85, 27) <= 5; angryBirdLarge(85, 28) <= 5; angryBirdLarge(85, 29) <= 5; angryBirdLarge(85, 30) <= 4; angryBirdLarge(85, 31) <= 4; angryBirdLarge(85, 32) <= 4; angryBirdLarge(85, 33) <= 4; angryBirdLarge(85, 34) <= 4; angryBirdLarge(85, 35) <= 4; angryBirdLarge(85, 36) <= 4; angryBirdLarge(85, 37) <= 4; angryBirdLarge(85, 38) <= 4; angryBirdLarge(85, 39) <= 4; angryBirdLarge(85, 40) <= 4; angryBirdLarge(85, 41) <= 4; angryBirdLarge(85, 42) <= 4; angryBirdLarge(85, 43) <= 4; angryBirdLarge(85, 44) <= 4; angryBirdLarge(85, 45) <= 4; angryBirdLarge(85, 46) <= 4; angryBirdLarge(85, 47) <= 4; angryBirdLarge(85, 48) <= 4; angryBirdLarge(85, 49) <= 4; angryBirdLarge(85, 50) <= 4; angryBirdLarge(85, 51) <= 4; angryBirdLarge(85, 52) <= 4; angryBirdLarge(85, 53) <= 4; angryBirdLarge(85, 54) <= 4; angryBirdLarge(85, 55) <= 4; angryBirdLarge(85, 56) <= 4; angryBirdLarge(85, 57) <= 4; angryBirdLarge(85, 58) <= 4; angryBirdLarge(85, 59) <= 4; angryBirdLarge(85, 60) <= 4; angryBirdLarge(85, 61) <= 4; angryBirdLarge(85, 62) <= 4; angryBirdLarge(85, 63) <= 4; angryBirdLarge(85, 64) <= 4; angryBirdLarge(85, 65) <= 4; angryBirdLarge(85, 66) <= 4; angryBirdLarge(85, 67) <= 4; angryBirdLarge(85, 68) <= 4; angryBirdLarge(85, 69) <= 4; angryBirdLarge(85, 70) <= 4; angryBirdLarge(85, 71) <= 4; angryBirdLarge(85, 72) <= 4; angryBirdLarge(85, 73) <= 4; angryBirdLarge(85, 74) <= 4; angryBirdLarge(85, 75) <= 4; angryBirdLarge(85, 76) <= 4; angryBirdLarge(85, 77) <= 4; angryBirdLarge(85, 78) <= 4; angryBirdLarge(85, 79) <= 4; angryBirdLarge(85, 80) <= 4; angryBirdLarge(85, 81) <= 4; angryBirdLarge(85, 82) <= 4; angryBirdLarge(85, 83) <= 4; angryBirdLarge(85, 84) <= 5; angryBirdLarge(85, 85) <= 5; angryBirdLarge(85, 86) <= 5; angryBirdLarge(85, 87) <= 5; angryBirdLarge(85, 88) <= 5; angryBirdLarge(85, 89) <= 5; angryBirdLarge(85, 90) <= 2; angryBirdLarge(85, 91) <= 2; angryBirdLarge(85, 92) <= 2; angryBirdLarge(85, 93) <= 2; angryBirdLarge(85, 94) <= 2; angryBirdLarge(85, 95) <= 2; angryBirdLarge(85, 96) <= 2; angryBirdLarge(85, 97) <= 2; angryBirdLarge(85, 98) <= 2; angryBirdLarge(85, 99) <= 2; angryBirdLarge(85, 100) <= 2; angryBirdLarge(85, 101) <= 2; angryBirdLarge(85, 102) <= 2; angryBirdLarge(85, 103) <= 2; angryBirdLarge(85, 104) <= 2; angryBirdLarge(85, 105) <= 2; angryBirdLarge(85, 106) <= 2; angryBirdLarge(85, 107) <= 2; angryBirdLarge(85, 108) <= 5; angryBirdLarge(85, 109) <= 5; angryBirdLarge(85, 110) <= 5; angryBirdLarge(85, 111) <= 5; angryBirdLarge(85, 112) <= 5; angryBirdLarge(85, 113) <= 5; angryBirdLarge(85, 114) <= 5; angryBirdLarge(85, 115) <= 5; angryBirdLarge(85, 116) <= 5; angryBirdLarge(85, 117) <= 5; angryBirdLarge(85, 118) <= 5; angryBirdLarge(85, 119) <= 5; angryBirdLarge(85, 120) <= 2; angryBirdLarge(85, 121) <= 2; angryBirdLarge(85, 122) <= 2; angryBirdLarge(85, 123) <= 2; angryBirdLarge(85, 124) <= 2; angryBirdLarge(85, 125) <= 2; angryBirdLarge(85, 126) <= 2; angryBirdLarge(85, 127) <= 2; angryBirdLarge(85, 128) <= 2; angryBirdLarge(85, 129) <= 2; angryBirdLarge(85, 130) <= 2; angryBirdLarge(85, 131) <= 2; angryBirdLarge(85, 132) <= 5; angryBirdLarge(85, 133) <= 5; angryBirdLarge(85, 134) <= 5; angryBirdLarge(85, 135) <= 5; angryBirdLarge(85, 136) <= 5; angryBirdLarge(85, 137) <= 5; angryBirdLarge(85, 138) <= 4; angryBirdLarge(85, 139) <= 4; angryBirdLarge(85, 140) <= 4; angryBirdLarge(85, 141) <= 4; angryBirdLarge(85, 142) <= 4; angryBirdLarge(85, 143) <= 4; angryBirdLarge(85, 144) <= 5; angryBirdLarge(85, 145) <= 5; angryBirdLarge(85, 146) <= 5; angryBirdLarge(85, 147) <= 5; angryBirdLarge(85, 148) <= 5; angryBirdLarge(85, 149) <= 5; 
angryBirdLarge(86, 0) <= 0; angryBirdLarge(86, 1) <= 0; angryBirdLarge(86, 2) <= 0; angryBirdLarge(86, 3) <= 0; angryBirdLarge(86, 4) <= 0; angryBirdLarge(86, 5) <= 0; angryBirdLarge(86, 6) <= 5; angryBirdLarge(86, 7) <= 5; angryBirdLarge(86, 8) <= 5; angryBirdLarge(86, 9) <= 5; angryBirdLarge(86, 10) <= 5; angryBirdLarge(86, 11) <= 5; angryBirdLarge(86, 12) <= 5; angryBirdLarge(86, 13) <= 5; angryBirdLarge(86, 14) <= 5; angryBirdLarge(86, 15) <= 5; angryBirdLarge(86, 16) <= 5; angryBirdLarge(86, 17) <= 5; angryBirdLarge(86, 18) <= 5; angryBirdLarge(86, 19) <= 5; angryBirdLarge(86, 20) <= 5; angryBirdLarge(86, 21) <= 5; angryBirdLarge(86, 22) <= 5; angryBirdLarge(86, 23) <= 5; angryBirdLarge(86, 24) <= 5; angryBirdLarge(86, 25) <= 5; angryBirdLarge(86, 26) <= 5; angryBirdLarge(86, 27) <= 5; angryBirdLarge(86, 28) <= 5; angryBirdLarge(86, 29) <= 5; angryBirdLarge(86, 30) <= 4; angryBirdLarge(86, 31) <= 4; angryBirdLarge(86, 32) <= 4; angryBirdLarge(86, 33) <= 4; angryBirdLarge(86, 34) <= 4; angryBirdLarge(86, 35) <= 4; angryBirdLarge(86, 36) <= 4; angryBirdLarge(86, 37) <= 4; angryBirdLarge(86, 38) <= 4; angryBirdLarge(86, 39) <= 4; angryBirdLarge(86, 40) <= 4; angryBirdLarge(86, 41) <= 4; angryBirdLarge(86, 42) <= 4; angryBirdLarge(86, 43) <= 4; angryBirdLarge(86, 44) <= 4; angryBirdLarge(86, 45) <= 4; angryBirdLarge(86, 46) <= 4; angryBirdLarge(86, 47) <= 4; angryBirdLarge(86, 48) <= 4; angryBirdLarge(86, 49) <= 4; angryBirdLarge(86, 50) <= 4; angryBirdLarge(86, 51) <= 4; angryBirdLarge(86, 52) <= 4; angryBirdLarge(86, 53) <= 4; angryBirdLarge(86, 54) <= 4; angryBirdLarge(86, 55) <= 4; angryBirdLarge(86, 56) <= 4; angryBirdLarge(86, 57) <= 4; angryBirdLarge(86, 58) <= 4; angryBirdLarge(86, 59) <= 4; angryBirdLarge(86, 60) <= 4; angryBirdLarge(86, 61) <= 4; angryBirdLarge(86, 62) <= 4; angryBirdLarge(86, 63) <= 4; angryBirdLarge(86, 64) <= 4; angryBirdLarge(86, 65) <= 4; angryBirdLarge(86, 66) <= 4; angryBirdLarge(86, 67) <= 4; angryBirdLarge(86, 68) <= 4; angryBirdLarge(86, 69) <= 4; angryBirdLarge(86, 70) <= 4; angryBirdLarge(86, 71) <= 4; angryBirdLarge(86, 72) <= 4; angryBirdLarge(86, 73) <= 4; angryBirdLarge(86, 74) <= 4; angryBirdLarge(86, 75) <= 4; angryBirdLarge(86, 76) <= 4; angryBirdLarge(86, 77) <= 4; angryBirdLarge(86, 78) <= 4; angryBirdLarge(86, 79) <= 4; angryBirdLarge(86, 80) <= 4; angryBirdLarge(86, 81) <= 4; angryBirdLarge(86, 82) <= 4; angryBirdLarge(86, 83) <= 4; angryBirdLarge(86, 84) <= 5; angryBirdLarge(86, 85) <= 5; angryBirdLarge(86, 86) <= 5; angryBirdLarge(86, 87) <= 5; angryBirdLarge(86, 88) <= 5; angryBirdLarge(86, 89) <= 5; angryBirdLarge(86, 90) <= 2; angryBirdLarge(86, 91) <= 2; angryBirdLarge(86, 92) <= 2; angryBirdLarge(86, 93) <= 2; angryBirdLarge(86, 94) <= 2; angryBirdLarge(86, 95) <= 2; angryBirdLarge(86, 96) <= 2; angryBirdLarge(86, 97) <= 2; angryBirdLarge(86, 98) <= 2; angryBirdLarge(86, 99) <= 2; angryBirdLarge(86, 100) <= 2; angryBirdLarge(86, 101) <= 2; angryBirdLarge(86, 102) <= 2; angryBirdLarge(86, 103) <= 2; angryBirdLarge(86, 104) <= 2; angryBirdLarge(86, 105) <= 2; angryBirdLarge(86, 106) <= 2; angryBirdLarge(86, 107) <= 2; angryBirdLarge(86, 108) <= 5; angryBirdLarge(86, 109) <= 5; angryBirdLarge(86, 110) <= 5; angryBirdLarge(86, 111) <= 5; angryBirdLarge(86, 112) <= 5; angryBirdLarge(86, 113) <= 5; angryBirdLarge(86, 114) <= 5; angryBirdLarge(86, 115) <= 5; angryBirdLarge(86, 116) <= 5; angryBirdLarge(86, 117) <= 5; angryBirdLarge(86, 118) <= 5; angryBirdLarge(86, 119) <= 5; angryBirdLarge(86, 120) <= 2; angryBirdLarge(86, 121) <= 2; angryBirdLarge(86, 122) <= 2; angryBirdLarge(86, 123) <= 2; angryBirdLarge(86, 124) <= 2; angryBirdLarge(86, 125) <= 2; angryBirdLarge(86, 126) <= 2; angryBirdLarge(86, 127) <= 2; angryBirdLarge(86, 128) <= 2; angryBirdLarge(86, 129) <= 2; angryBirdLarge(86, 130) <= 2; angryBirdLarge(86, 131) <= 2; angryBirdLarge(86, 132) <= 5; angryBirdLarge(86, 133) <= 5; angryBirdLarge(86, 134) <= 5; angryBirdLarge(86, 135) <= 5; angryBirdLarge(86, 136) <= 5; angryBirdLarge(86, 137) <= 5; angryBirdLarge(86, 138) <= 4; angryBirdLarge(86, 139) <= 4; angryBirdLarge(86, 140) <= 4; angryBirdLarge(86, 141) <= 4; angryBirdLarge(86, 142) <= 4; angryBirdLarge(86, 143) <= 4; angryBirdLarge(86, 144) <= 5; angryBirdLarge(86, 145) <= 5; angryBirdLarge(86, 146) <= 5; angryBirdLarge(86, 147) <= 5; angryBirdLarge(86, 148) <= 5; angryBirdLarge(86, 149) <= 5; 
angryBirdLarge(87, 0) <= 0; angryBirdLarge(87, 1) <= 0; angryBirdLarge(87, 2) <= 0; angryBirdLarge(87, 3) <= 0; angryBirdLarge(87, 4) <= 0; angryBirdLarge(87, 5) <= 0; angryBirdLarge(87, 6) <= 5; angryBirdLarge(87, 7) <= 5; angryBirdLarge(87, 8) <= 5; angryBirdLarge(87, 9) <= 5; angryBirdLarge(87, 10) <= 5; angryBirdLarge(87, 11) <= 5; angryBirdLarge(87, 12) <= 5; angryBirdLarge(87, 13) <= 5; angryBirdLarge(87, 14) <= 5; angryBirdLarge(87, 15) <= 5; angryBirdLarge(87, 16) <= 5; angryBirdLarge(87, 17) <= 5; angryBirdLarge(87, 18) <= 5; angryBirdLarge(87, 19) <= 5; angryBirdLarge(87, 20) <= 5; angryBirdLarge(87, 21) <= 5; angryBirdLarge(87, 22) <= 5; angryBirdLarge(87, 23) <= 5; angryBirdLarge(87, 24) <= 5; angryBirdLarge(87, 25) <= 5; angryBirdLarge(87, 26) <= 5; angryBirdLarge(87, 27) <= 5; angryBirdLarge(87, 28) <= 5; angryBirdLarge(87, 29) <= 5; angryBirdLarge(87, 30) <= 4; angryBirdLarge(87, 31) <= 4; angryBirdLarge(87, 32) <= 4; angryBirdLarge(87, 33) <= 4; angryBirdLarge(87, 34) <= 4; angryBirdLarge(87, 35) <= 4; angryBirdLarge(87, 36) <= 4; angryBirdLarge(87, 37) <= 4; angryBirdLarge(87, 38) <= 4; angryBirdLarge(87, 39) <= 4; angryBirdLarge(87, 40) <= 4; angryBirdLarge(87, 41) <= 4; angryBirdLarge(87, 42) <= 4; angryBirdLarge(87, 43) <= 4; angryBirdLarge(87, 44) <= 4; angryBirdLarge(87, 45) <= 4; angryBirdLarge(87, 46) <= 4; angryBirdLarge(87, 47) <= 4; angryBirdLarge(87, 48) <= 4; angryBirdLarge(87, 49) <= 4; angryBirdLarge(87, 50) <= 4; angryBirdLarge(87, 51) <= 4; angryBirdLarge(87, 52) <= 4; angryBirdLarge(87, 53) <= 4; angryBirdLarge(87, 54) <= 4; angryBirdLarge(87, 55) <= 4; angryBirdLarge(87, 56) <= 4; angryBirdLarge(87, 57) <= 4; angryBirdLarge(87, 58) <= 4; angryBirdLarge(87, 59) <= 4; angryBirdLarge(87, 60) <= 4; angryBirdLarge(87, 61) <= 4; angryBirdLarge(87, 62) <= 4; angryBirdLarge(87, 63) <= 4; angryBirdLarge(87, 64) <= 4; angryBirdLarge(87, 65) <= 4; angryBirdLarge(87, 66) <= 4; angryBirdLarge(87, 67) <= 4; angryBirdLarge(87, 68) <= 4; angryBirdLarge(87, 69) <= 4; angryBirdLarge(87, 70) <= 4; angryBirdLarge(87, 71) <= 4; angryBirdLarge(87, 72) <= 4; angryBirdLarge(87, 73) <= 4; angryBirdLarge(87, 74) <= 4; angryBirdLarge(87, 75) <= 4; angryBirdLarge(87, 76) <= 4; angryBirdLarge(87, 77) <= 4; angryBirdLarge(87, 78) <= 4; angryBirdLarge(87, 79) <= 4; angryBirdLarge(87, 80) <= 4; angryBirdLarge(87, 81) <= 4; angryBirdLarge(87, 82) <= 4; angryBirdLarge(87, 83) <= 4; angryBirdLarge(87, 84) <= 5; angryBirdLarge(87, 85) <= 5; angryBirdLarge(87, 86) <= 5; angryBirdLarge(87, 87) <= 5; angryBirdLarge(87, 88) <= 5; angryBirdLarge(87, 89) <= 5; angryBirdLarge(87, 90) <= 2; angryBirdLarge(87, 91) <= 2; angryBirdLarge(87, 92) <= 2; angryBirdLarge(87, 93) <= 2; angryBirdLarge(87, 94) <= 2; angryBirdLarge(87, 95) <= 2; angryBirdLarge(87, 96) <= 2; angryBirdLarge(87, 97) <= 2; angryBirdLarge(87, 98) <= 2; angryBirdLarge(87, 99) <= 2; angryBirdLarge(87, 100) <= 2; angryBirdLarge(87, 101) <= 2; angryBirdLarge(87, 102) <= 2; angryBirdLarge(87, 103) <= 2; angryBirdLarge(87, 104) <= 2; angryBirdLarge(87, 105) <= 2; angryBirdLarge(87, 106) <= 2; angryBirdLarge(87, 107) <= 2; angryBirdLarge(87, 108) <= 5; angryBirdLarge(87, 109) <= 5; angryBirdLarge(87, 110) <= 5; angryBirdLarge(87, 111) <= 5; angryBirdLarge(87, 112) <= 5; angryBirdLarge(87, 113) <= 5; angryBirdLarge(87, 114) <= 5; angryBirdLarge(87, 115) <= 5; angryBirdLarge(87, 116) <= 5; angryBirdLarge(87, 117) <= 5; angryBirdLarge(87, 118) <= 5; angryBirdLarge(87, 119) <= 5; angryBirdLarge(87, 120) <= 2; angryBirdLarge(87, 121) <= 2; angryBirdLarge(87, 122) <= 2; angryBirdLarge(87, 123) <= 2; angryBirdLarge(87, 124) <= 2; angryBirdLarge(87, 125) <= 2; angryBirdLarge(87, 126) <= 2; angryBirdLarge(87, 127) <= 2; angryBirdLarge(87, 128) <= 2; angryBirdLarge(87, 129) <= 2; angryBirdLarge(87, 130) <= 2; angryBirdLarge(87, 131) <= 2; angryBirdLarge(87, 132) <= 5; angryBirdLarge(87, 133) <= 5; angryBirdLarge(87, 134) <= 5; angryBirdLarge(87, 135) <= 5; angryBirdLarge(87, 136) <= 5; angryBirdLarge(87, 137) <= 5; angryBirdLarge(87, 138) <= 4; angryBirdLarge(87, 139) <= 4; angryBirdLarge(87, 140) <= 4; angryBirdLarge(87, 141) <= 4; angryBirdLarge(87, 142) <= 4; angryBirdLarge(87, 143) <= 4; angryBirdLarge(87, 144) <= 5; angryBirdLarge(87, 145) <= 5; angryBirdLarge(87, 146) <= 5; angryBirdLarge(87, 147) <= 5; angryBirdLarge(87, 148) <= 5; angryBirdLarge(87, 149) <= 5; 
angryBirdLarge(88, 0) <= 0; angryBirdLarge(88, 1) <= 0; angryBirdLarge(88, 2) <= 0; angryBirdLarge(88, 3) <= 0; angryBirdLarge(88, 4) <= 0; angryBirdLarge(88, 5) <= 0; angryBirdLarge(88, 6) <= 5; angryBirdLarge(88, 7) <= 5; angryBirdLarge(88, 8) <= 5; angryBirdLarge(88, 9) <= 5; angryBirdLarge(88, 10) <= 5; angryBirdLarge(88, 11) <= 5; angryBirdLarge(88, 12) <= 5; angryBirdLarge(88, 13) <= 5; angryBirdLarge(88, 14) <= 5; angryBirdLarge(88, 15) <= 5; angryBirdLarge(88, 16) <= 5; angryBirdLarge(88, 17) <= 5; angryBirdLarge(88, 18) <= 5; angryBirdLarge(88, 19) <= 5; angryBirdLarge(88, 20) <= 5; angryBirdLarge(88, 21) <= 5; angryBirdLarge(88, 22) <= 5; angryBirdLarge(88, 23) <= 5; angryBirdLarge(88, 24) <= 5; angryBirdLarge(88, 25) <= 5; angryBirdLarge(88, 26) <= 5; angryBirdLarge(88, 27) <= 5; angryBirdLarge(88, 28) <= 5; angryBirdLarge(88, 29) <= 5; angryBirdLarge(88, 30) <= 4; angryBirdLarge(88, 31) <= 4; angryBirdLarge(88, 32) <= 4; angryBirdLarge(88, 33) <= 4; angryBirdLarge(88, 34) <= 4; angryBirdLarge(88, 35) <= 4; angryBirdLarge(88, 36) <= 4; angryBirdLarge(88, 37) <= 4; angryBirdLarge(88, 38) <= 4; angryBirdLarge(88, 39) <= 4; angryBirdLarge(88, 40) <= 4; angryBirdLarge(88, 41) <= 4; angryBirdLarge(88, 42) <= 4; angryBirdLarge(88, 43) <= 4; angryBirdLarge(88, 44) <= 4; angryBirdLarge(88, 45) <= 4; angryBirdLarge(88, 46) <= 4; angryBirdLarge(88, 47) <= 4; angryBirdLarge(88, 48) <= 4; angryBirdLarge(88, 49) <= 4; angryBirdLarge(88, 50) <= 4; angryBirdLarge(88, 51) <= 4; angryBirdLarge(88, 52) <= 4; angryBirdLarge(88, 53) <= 4; angryBirdLarge(88, 54) <= 4; angryBirdLarge(88, 55) <= 4; angryBirdLarge(88, 56) <= 4; angryBirdLarge(88, 57) <= 4; angryBirdLarge(88, 58) <= 4; angryBirdLarge(88, 59) <= 4; angryBirdLarge(88, 60) <= 4; angryBirdLarge(88, 61) <= 4; angryBirdLarge(88, 62) <= 4; angryBirdLarge(88, 63) <= 4; angryBirdLarge(88, 64) <= 4; angryBirdLarge(88, 65) <= 4; angryBirdLarge(88, 66) <= 4; angryBirdLarge(88, 67) <= 4; angryBirdLarge(88, 68) <= 4; angryBirdLarge(88, 69) <= 4; angryBirdLarge(88, 70) <= 4; angryBirdLarge(88, 71) <= 4; angryBirdLarge(88, 72) <= 4; angryBirdLarge(88, 73) <= 4; angryBirdLarge(88, 74) <= 4; angryBirdLarge(88, 75) <= 4; angryBirdLarge(88, 76) <= 4; angryBirdLarge(88, 77) <= 4; angryBirdLarge(88, 78) <= 4; angryBirdLarge(88, 79) <= 4; angryBirdLarge(88, 80) <= 4; angryBirdLarge(88, 81) <= 4; angryBirdLarge(88, 82) <= 4; angryBirdLarge(88, 83) <= 4; angryBirdLarge(88, 84) <= 5; angryBirdLarge(88, 85) <= 5; angryBirdLarge(88, 86) <= 5; angryBirdLarge(88, 87) <= 5; angryBirdLarge(88, 88) <= 5; angryBirdLarge(88, 89) <= 5; angryBirdLarge(88, 90) <= 2; angryBirdLarge(88, 91) <= 2; angryBirdLarge(88, 92) <= 2; angryBirdLarge(88, 93) <= 2; angryBirdLarge(88, 94) <= 2; angryBirdLarge(88, 95) <= 2; angryBirdLarge(88, 96) <= 2; angryBirdLarge(88, 97) <= 2; angryBirdLarge(88, 98) <= 2; angryBirdLarge(88, 99) <= 2; angryBirdLarge(88, 100) <= 2; angryBirdLarge(88, 101) <= 2; angryBirdLarge(88, 102) <= 2; angryBirdLarge(88, 103) <= 2; angryBirdLarge(88, 104) <= 2; angryBirdLarge(88, 105) <= 2; angryBirdLarge(88, 106) <= 2; angryBirdLarge(88, 107) <= 2; angryBirdLarge(88, 108) <= 5; angryBirdLarge(88, 109) <= 5; angryBirdLarge(88, 110) <= 5; angryBirdLarge(88, 111) <= 5; angryBirdLarge(88, 112) <= 5; angryBirdLarge(88, 113) <= 5; angryBirdLarge(88, 114) <= 5; angryBirdLarge(88, 115) <= 5; angryBirdLarge(88, 116) <= 5; angryBirdLarge(88, 117) <= 5; angryBirdLarge(88, 118) <= 5; angryBirdLarge(88, 119) <= 5; angryBirdLarge(88, 120) <= 2; angryBirdLarge(88, 121) <= 2; angryBirdLarge(88, 122) <= 2; angryBirdLarge(88, 123) <= 2; angryBirdLarge(88, 124) <= 2; angryBirdLarge(88, 125) <= 2; angryBirdLarge(88, 126) <= 2; angryBirdLarge(88, 127) <= 2; angryBirdLarge(88, 128) <= 2; angryBirdLarge(88, 129) <= 2; angryBirdLarge(88, 130) <= 2; angryBirdLarge(88, 131) <= 2; angryBirdLarge(88, 132) <= 5; angryBirdLarge(88, 133) <= 5; angryBirdLarge(88, 134) <= 5; angryBirdLarge(88, 135) <= 5; angryBirdLarge(88, 136) <= 5; angryBirdLarge(88, 137) <= 5; angryBirdLarge(88, 138) <= 4; angryBirdLarge(88, 139) <= 4; angryBirdLarge(88, 140) <= 4; angryBirdLarge(88, 141) <= 4; angryBirdLarge(88, 142) <= 4; angryBirdLarge(88, 143) <= 4; angryBirdLarge(88, 144) <= 5; angryBirdLarge(88, 145) <= 5; angryBirdLarge(88, 146) <= 5; angryBirdLarge(88, 147) <= 5; angryBirdLarge(88, 148) <= 5; angryBirdLarge(88, 149) <= 5; 
angryBirdLarge(89, 0) <= 0; angryBirdLarge(89, 1) <= 0; angryBirdLarge(89, 2) <= 0; angryBirdLarge(89, 3) <= 0; angryBirdLarge(89, 4) <= 0; angryBirdLarge(89, 5) <= 0; angryBirdLarge(89, 6) <= 5; angryBirdLarge(89, 7) <= 5; angryBirdLarge(89, 8) <= 5; angryBirdLarge(89, 9) <= 5; angryBirdLarge(89, 10) <= 5; angryBirdLarge(89, 11) <= 5; angryBirdLarge(89, 12) <= 5; angryBirdLarge(89, 13) <= 5; angryBirdLarge(89, 14) <= 5; angryBirdLarge(89, 15) <= 5; angryBirdLarge(89, 16) <= 5; angryBirdLarge(89, 17) <= 5; angryBirdLarge(89, 18) <= 5; angryBirdLarge(89, 19) <= 5; angryBirdLarge(89, 20) <= 5; angryBirdLarge(89, 21) <= 5; angryBirdLarge(89, 22) <= 5; angryBirdLarge(89, 23) <= 5; angryBirdLarge(89, 24) <= 5; angryBirdLarge(89, 25) <= 5; angryBirdLarge(89, 26) <= 5; angryBirdLarge(89, 27) <= 5; angryBirdLarge(89, 28) <= 5; angryBirdLarge(89, 29) <= 5; angryBirdLarge(89, 30) <= 4; angryBirdLarge(89, 31) <= 4; angryBirdLarge(89, 32) <= 4; angryBirdLarge(89, 33) <= 4; angryBirdLarge(89, 34) <= 4; angryBirdLarge(89, 35) <= 4; angryBirdLarge(89, 36) <= 4; angryBirdLarge(89, 37) <= 4; angryBirdLarge(89, 38) <= 4; angryBirdLarge(89, 39) <= 4; angryBirdLarge(89, 40) <= 4; angryBirdLarge(89, 41) <= 4; angryBirdLarge(89, 42) <= 4; angryBirdLarge(89, 43) <= 4; angryBirdLarge(89, 44) <= 4; angryBirdLarge(89, 45) <= 4; angryBirdLarge(89, 46) <= 4; angryBirdLarge(89, 47) <= 4; angryBirdLarge(89, 48) <= 4; angryBirdLarge(89, 49) <= 4; angryBirdLarge(89, 50) <= 4; angryBirdLarge(89, 51) <= 4; angryBirdLarge(89, 52) <= 4; angryBirdLarge(89, 53) <= 4; angryBirdLarge(89, 54) <= 4; angryBirdLarge(89, 55) <= 4; angryBirdLarge(89, 56) <= 4; angryBirdLarge(89, 57) <= 4; angryBirdLarge(89, 58) <= 4; angryBirdLarge(89, 59) <= 4; angryBirdLarge(89, 60) <= 4; angryBirdLarge(89, 61) <= 4; angryBirdLarge(89, 62) <= 4; angryBirdLarge(89, 63) <= 4; angryBirdLarge(89, 64) <= 4; angryBirdLarge(89, 65) <= 4; angryBirdLarge(89, 66) <= 4; angryBirdLarge(89, 67) <= 4; angryBirdLarge(89, 68) <= 4; angryBirdLarge(89, 69) <= 4; angryBirdLarge(89, 70) <= 4; angryBirdLarge(89, 71) <= 4; angryBirdLarge(89, 72) <= 4; angryBirdLarge(89, 73) <= 4; angryBirdLarge(89, 74) <= 4; angryBirdLarge(89, 75) <= 4; angryBirdLarge(89, 76) <= 4; angryBirdLarge(89, 77) <= 4; angryBirdLarge(89, 78) <= 4; angryBirdLarge(89, 79) <= 4; angryBirdLarge(89, 80) <= 4; angryBirdLarge(89, 81) <= 4; angryBirdLarge(89, 82) <= 4; angryBirdLarge(89, 83) <= 4; angryBirdLarge(89, 84) <= 5; angryBirdLarge(89, 85) <= 5; angryBirdLarge(89, 86) <= 5; angryBirdLarge(89, 87) <= 5; angryBirdLarge(89, 88) <= 5; angryBirdLarge(89, 89) <= 5; angryBirdLarge(89, 90) <= 2; angryBirdLarge(89, 91) <= 2; angryBirdLarge(89, 92) <= 2; angryBirdLarge(89, 93) <= 2; angryBirdLarge(89, 94) <= 2; angryBirdLarge(89, 95) <= 2; angryBirdLarge(89, 96) <= 2; angryBirdLarge(89, 97) <= 2; angryBirdLarge(89, 98) <= 2; angryBirdLarge(89, 99) <= 2; angryBirdLarge(89, 100) <= 2; angryBirdLarge(89, 101) <= 2; angryBirdLarge(89, 102) <= 2; angryBirdLarge(89, 103) <= 2; angryBirdLarge(89, 104) <= 2; angryBirdLarge(89, 105) <= 2; angryBirdLarge(89, 106) <= 2; angryBirdLarge(89, 107) <= 2; angryBirdLarge(89, 108) <= 5; angryBirdLarge(89, 109) <= 5; angryBirdLarge(89, 110) <= 5; angryBirdLarge(89, 111) <= 5; angryBirdLarge(89, 112) <= 5; angryBirdLarge(89, 113) <= 5; angryBirdLarge(89, 114) <= 5; angryBirdLarge(89, 115) <= 5; angryBirdLarge(89, 116) <= 5; angryBirdLarge(89, 117) <= 5; angryBirdLarge(89, 118) <= 5; angryBirdLarge(89, 119) <= 5; angryBirdLarge(89, 120) <= 2; angryBirdLarge(89, 121) <= 2; angryBirdLarge(89, 122) <= 2; angryBirdLarge(89, 123) <= 2; angryBirdLarge(89, 124) <= 2; angryBirdLarge(89, 125) <= 2; angryBirdLarge(89, 126) <= 2; angryBirdLarge(89, 127) <= 2; angryBirdLarge(89, 128) <= 2; angryBirdLarge(89, 129) <= 2; angryBirdLarge(89, 130) <= 2; angryBirdLarge(89, 131) <= 2; angryBirdLarge(89, 132) <= 5; angryBirdLarge(89, 133) <= 5; angryBirdLarge(89, 134) <= 5; angryBirdLarge(89, 135) <= 5; angryBirdLarge(89, 136) <= 5; angryBirdLarge(89, 137) <= 5; angryBirdLarge(89, 138) <= 4; angryBirdLarge(89, 139) <= 4; angryBirdLarge(89, 140) <= 4; angryBirdLarge(89, 141) <= 4; angryBirdLarge(89, 142) <= 4; angryBirdLarge(89, 143) <= 4; angryBirdLarge(89, 144) <= 5; angryBirdLarge(89, 145) <= 5; angryBirdLarge(89, 146) <= 5; angryBirdLarge(89, 147) <= 5; angryBirdLarge(89, 148) <= 5; angryBirdLarge(89, 149) <= 5; 
angryBirdLarge(90, 0) <= 0; angryBirdLarge(90, 1) <= 0; angryBirdLarge(90, 2) <= 0; angryBirdLarge(90, 3) <= 0; angryBirdLarge(90, 4) <= 0; angryBirdLarge(90, 5) <= 0; angryBirdLarge(90, 6) <= 0; angryBirdLarge(90, 7) <= 0; angryBirdLarge(90, 8) <= 0; angryBirdLarge(90, 9) <= 0; angryBirdLarge(90, 10) <= 0; angryBirdLarge(90, 11) <= 0; angryBirdLarge(90, 12) <= 0; angryBirdLarge(90, 13) <= 0; angryBirdLarge(90, 14) <= 0; angryBirdLarge(90, 15) <= 0; angryBirdLarge(90, 16) <= 0; angryBirdLarge(90, 17) <= 0; angryBirdLarge(90, 18) <= 5; angryBirdLarge(90, 19) <= 5; angryBirdLarge(90, 20) <= 5; angryBirdLarge(90, 21) <= 5; angryBirdLarge(90, 22) <= 5; angryBirdLarge(90, 23) <= 5; angryBirdLarge(90, 24) <= 5; angryBirdLarge(90, 25) <= 5; angryBirdLarge(90, 26) <= 5; angryBirdLarge(90, 27) <= 5; angryBirdLarge(90, 28) <= 5; angryBirdLarge(90, 29) <= 5; angryBirdLarge(90, 30) <= 4; angryBirdLarge(90, 31) <= 4; angryBirdLarge(90, 32) <= 4; angryBirdLarge(90, 33) <= 4; angryBirdLarge(90, 34) <= 4; angryBirdLarge(90, 35) <= 4; angryBirdLarge(90, 36) <= 4; angryBirdLarge(90, 37) <= 4; angryBirdLarge(90, 38) <= 4; angryBirdLarge(90, 39) <= 4; angryBirdLarge(90, 40) <= 4; angryBirdLarge(90, 41) <= 4; angryBirdLarge(90, 42) <= 4; angryBirdLarge(90, 43) <= 4; angryBirdLarge(90, 44) <= 4; angryBirdLarge(90, 45) <= 4; angryBirdLarge(90, 46) <= 4; angryBirdLarge(90, 47) <= 4; angryBirdLarge(90, 48) <= 4; angryBirdLarge(90, 49) <= 4; angryBirdLarge(90, 50) <= 4; angryBirdLarge(90, 51) <= 4; angryBirdLarge(90, 52) <= 4; angryBirdLarge(90, 53) <= 4; angryBirdLarge(90, 54) <= 4; angryBirdLarge(90, 55) <= 4; angryBirdLarge(90, 56) <= 4; angryBirdLarge(90, 57) <= 4; angryBirdLarge(90, 58) <= 4; angryBirdLarge(90, 59) <= 4; angryBirdLarge(90, 60) <= 4; angryBirdLarge(90, 61) <= 4; angryBirdLarge(90, 62) <= 4; angryBirdLarge(90, 63) <= 4; angryBirdLarge(90, 64) <= 4; angryBirdLarge(90, 65) <= 4; angryBirdLarge(90, 66) <= 4; angryBirdLarge(90, 67) <= 4; angryBirdLarge(90, 68) <= 4; angryBirdLarge(90, 69) <= 4; angryBirdLarge(90, 70) <= 4; angryBirdLarge(90, 71) <= 4; angryBirdLarge(90, 72) <= 4; angryBirdLarge(90, 73) <= 4; angryBirdLarge(90, 74) <= 4; angryBirdLarge(90, 75) <= 4; angryBirdLarge(90, 76) <= 4; angryBirdLarge(90, 77) <= 4; angryBirdLarge(90, 78) <= 4; angryBirdLarge(90, 79) <= 4; angryBirdLarge(90, 80) <= 4; angryBirdLarge(90, 81) <= 4; angryBirdLarge(90, 82) <= 4; angryBirdLarge(90, 83) <= 4; angryBirdLarge(90, 84) <= 4; angryBirdLarge(90, 85) <= 4; angryBirdLarge(90, 86) <= 4; angryBirdLarge(90, 87) <= 4; angryBirdLarge(90, 88) <= 4; angryBirdLarge(90, 89) <= 4; angryBirdLarge(90, 90) <= 5; angryBirdLarge(90, 91) <= 5; angryBirdLarge(90, 92) <= 5; angryBirdLarge(90, 93) <= 5; angryBirdLarge(90, 94) <= 5; angryBirdLarge(90, 95) <= 5; angryBirdLarge(90, 96) <= 5; angryBirdLarge(90, 97) <= 5; angryBirdLarge(90, 98) <= 5; angryBirdLarge(90, 99) <= 5; angryBirdLarge(90, 100) <= 5; angryBirdLarge(90, 101) <= 5; angryBirdLarge(90, 102) <= 3; angryBirdLarge(90, 103) <= 3; angryBirdLarge(90, 104) <= 3; angryBirdLarge(90, 105) <= 3; angryBirdLarge(90, 106) <= 3; angryBirdLarge(90, 107) <= 3; angryBirdLarge(90, 108) <= 3; angryBirdLarge(90, 109) <= 3; angryBirdLarge(90, 110) <= 3; angryBirdLarge(90, 111) <= 3; angryBirdLarge(90, 112) <= 3; angryBirdLarge(90, 113) <= 3; angryBirdLarge(90, 114) <= 3; angryBirdLarge(90, 115) <= 3; angryBirdLarge(90, 116) <= 3; angryBirdLarge(90, 117) <= 3; angryBirdLarge(90, 118) <= 3; angryBirdLarge(90, 119) <= 3; angryBirdLarge(90, 120) <= 5; angryBirdLarge(90, 121) <= 5; angryBirdLarge(90, 122) <= 5; angryBirdLarge(90, 123) <= 5; angryBirdLarge(90, 124) <= 5; angryBirdLarge(90, 125) <= 5; angryBirdLarge(90, 126) <= 5; angryBirdLarge(90, 127) <= 5; angryBirdLarge(90, 128) <= 5; angryBirdLarge(90, 129) <= 5; angryBirdLarge(90, 130) <= 5; angryBirdLarge(90, 131) <= 5; angryBirdLarge(90, 132) <= 4; angryBirdLarge(90, 133) <= 4; angryBirdLarge(90, 134) <= 4; angryBirdLarge(90, 135) <= 4; angryBirdLarge(90, 136) <= 4; angryBirdLarge(90, 137) <= 4; angryBirdLarge(90, 138) <= 4; angryBirdLarge(90, 139) <= 4; angryBirdLarge(90, 140) <= 4; angryBirdLarge(90, 141) <= 4; angryBirdLarge(90, 142) <= 4; angryBirdLarge(90, 143) <= 4; angryBirdLarge(90, 144) <= 5; angryBirdLarge(90, 145) <= 5; angryBirdLarge(90, 146) <= 5; angryBirdLarge(90, 147) <= 5; angryBirdLarge(90, 148) <= 5; angryBirdLarge(90, 149) <= 5; 
angryBirdLarge(91, 0) <= 0; angryBirdLarge(91, 1) <= 0; angryBirdLarge(91, 2) <= 0; angryBirdLarge(91, 3) <= 0; angryBirdLarge(91, 4) <= 0; angryBirdLarge(91, 5) <= 0; angryBirdLarge(91, 6) <= 0; angryBirdLarge(91, 7) <= 0; angryBirdLarge(91, 8) <= 0; angryBirdLarge(91, 9) <= 0; angryBirdLarge(91, 10) <= 0; angryBirdLarge(91, 11) <= 0; angryBirdLarge(91, 12) <= 0; angryBirdLarge(91, 13) <= 0; angryBirdLarge(91, 14) <= 0; angryBirdLarge(91, 15) <= 0; angryBirdLarge(91, 16) <= 0; angryBirdLarge(91, 17) <= 0; angryBirdLarge(91, 18) <= 5; angryBirdLarge(91, 19) <= 5; angryBirdLarge(91, 20) <= 5; angryBirdLarge(91, 21) <= 5; angryBirdLarge(91, 22) <= 5; angryBirdLarge(91, 23) <= 5; angryBirdLarge(91, 24) <= 5; angryBirdLarge(91, 25) <= 5; angryBirdLarge(91, 26) <= 5; angryBirdLarge(91, 27) <= 5; angryBirdLarge(91, 28) <= 5; angryBirdLarge(91, 29) <= 5; angryBirdLarge(91, 30) <= 4; angryBirdLarge(91, 31) <= 4; angryBirdLarge(91, 32) <= 4; angryBirdLarge(91, 33) <= 4; angryBirdLarge(91, 34) <= 4; angryBirdLarge(91, 35) <= 4; angryBirdLarge(91, 36) <= 4; angryBirdLarge(91, 37) <= 4; angryBirdLarge(91, 38) <= 4; angryBirdLarge(91, 39) <= 4; angryBirdLarge(91, 40) <= 4; angryBirdLarge(91, 41) <= 4; angryBirdLarge(91, 42) <= 4; angryBirdLarge(91, 43) <= 4; angryBirdLarge(91, 44) <= 4; angryBirdLarge(91, 45) <= 4; angryBirdLarge(91, 46) <= 4; angryBirdLarge(91, 47) <= 4; angryBirdLarge(91, 48) <= 4; angryBirdLarge(91, 49) <= 4; angryBirdLarge(91, 50) <= 4; angryBirdLarge(91, 51) <= 4; angryBirdLarge(91, 52) <= 4; angryBirdLarge(91, 53) <= 4; angryBirdLarge(91, 54) <= 4; angryBirdLarge(91, 55) <= 4; angryBirdLarge(91, 56) <= 4; angryBirdLarge(91, 57) <= 4; angryBirdLarge(91, 58) <= 4; angryBirdLarge(91, 59) <= 4; angryBirdLarge(91, 60) <= 4; angryBirdLarge(91, 61) <= 4; angryBirdLarge(91, 62) <= 4; angryBirdLarge(91, 63) <= 4; angryBirdLarge(91, 64) <= 4; angryBirdLarge(91, 65) <= 4; angryBirdLarge(91, 66) <= 4; angryBirdLarge(91, 67) <= 4; angryBirdLarge(91, 68) <= 4; angryBirdLarge(91, 69) <= 4; angryBirdLarge(91, 70) <= 4; angryBirdLarge(91, 71) <= 4; angryBirdLarge(91, 72) <= 4; angryBirdLarge(91, 73) <= 4; angryBirdLarge(91, 74) <= 4; angryBirdLarge(91, 75) <= 4; angryBirdLarge(91, 76) <= 4; angryBirdLarge(91, 77) <= 4; angryBirdLarge(91, 78) <= 4; angryBirdLarge(91, 79) <= 4; angryBirdLarge(91, 80) <= 4; angryBirdLarge(91, 81) <= 4; angryBirdLarge(91, 82) <= 4; angryBirdLarge(91, 83) <= 4; angryBirdLarge(91, 84) <= 4; angryBirdLarge(91, 85) <= 4; angryBirdLarge(91, 86) <= 4; angryBirdLarge(91, 87) <= 4; angryBirdLarge(91, 88) <= 4; angryBirdLarge(91, 89) <= 4; angryBirdLarge(91, 90) <= 5; angryBirdLarge(91, 91) <= 5; angryBirdLarge(91, 92) <= 5; angryBirdLarge(91, 93) <= 5; angryBirdLarge(91, 94) <= 5; angryBirdLarge(91, 95) <= 5; angryBirdLarge(91, 96) <= 5; angryBirdLarge(91, 97) <= 5; angryBirdLarge(91, 98) <= 5; angryBirdLarge(91, 99) <= 5; angryBirdLarge(91, 100) <= 5; angryBirdLarge(91, 101) <= 5; angryBirdLarge(91, 102) <= 3; angryBirdLarge(91, 103) <= 3; angryBirdLarge(91, 104) <= 3; angryBirdLarge(91, 105) <= 3; angryBirdLarge(91, 106) <= 3; angryBirdLarge(91, 107) <= 3; angryBirdLarge(91, 108) <= 3; angryBirdLarge(91, 109) <= 3; angryBirdLarge(91, 110) <= 3; angryBirdLarge(91, 111) <= 3; angryBirdLarge(91, 112) <= 3; angryBirdLarge(91, 113) <= 3; angryBirdLarge(91, 114) <= 3; angryBirdLarge(91, 115) <= 3; angryBirdLarge(91, 116) <= 3; angryBirdLarge(91, 117) <= 3; angryBirdLarge(91, 118) <= 3; angryBirdLarge(91, 119) <= 3; angryBirdLarge(91, 120) <= 5; angryBirdLarge(91, 121) <= 5; angryBirdLarge(91, 122) <= 5; angryBirdLarge(91, 123) <= 5; angryBirdLarge(91, 124) <= 5; angryBirdLarge(91, 125) <= 5; angryBirdLarge(91, 126) <= 5; angryBirdLarge(91, 127) <= 5; angryBirdLarge(91, 128) <= 5; angryBirdLarge(91, 129) <= 5; angryBirdLarge(91, 130) <= 5; angryBirdLarge(91, 131) <= 5; angryBirdLarge(91, 132) <= 4; angryBirdLarge(91, 133) <= 4; angryBirdLarge(91, 134) <= 4; angryBirdLarge(91, 135) <= 4; angryBirdLarge(91, 136) <= 4; angryBirdLarge(91, 137) <= 4; angryBirdLarge(91, 138) <= 4; angryBirdLarge(91, 139) <= 4; angryBirdLarge(91, 140) <= 4; angryBirdLarge(91, 141) <= 4; angryBirdLarge(91, 142) <= 4; angryBirdLarge(91, 143) <= 4; angryBirdLarge(91, 144) <= 5; angryBirdLarge(91, 145) <= 5; angryBirdLarge(91, 146) <= 5; angryBirdLarge(91, 147) <= 5; angryBirdLarge(91, 148) <= 5; angryBirdLarge(91, 149) <= 5; 
angryBirdLarge(92, 0) <= 0; angryBirdLarge(92, 1) <= 0; angryBirdLarge(92, 2) <= 0; angryBirdLarge(92, 3) <= 0; angryBirdLarge(92, 4) <= 0; angryBirdLarge(92, 5) <= 0; angryBirdLarge(92, 6) <= 0; angryBirdLarge(92, 7) <= 0; angryBirdLarge(92, 8) <= 0; angryBirdLarge(92, 9) <= 0; angryBirdLarge(92, 10) <= 0; angryBirdLarge(92, 11) <= 0; angryBirdLarge(92, 12) <= 0; angryBirdLarge(92, 13) <= 0; angryBirdLarge(92, 14) <= 0; angryBirdLarge(92, 15) <= 0; angryBirdLarge(92, 16) <= 0; angryBirdLarge(92, 17) <= 0; angryBirdLarge(92, 18) <= 5; angryBirdLarge(92, 19) <= 5; angryBirdLarge(92, 20) <= 5; angryBirdLarge(92, 21) <= 5; angryBirdLarge(92, 22) <= 5; angryBirdLarge(92, 23) <= 5; angryBirdLarge(92, 24) <= 5; angryBirdLarge(92, 25) <= 5; angryBirdLarge(92, 26) <= 5; angryBirdLarge(92, 27) <= 5; angryBirdLarge(92, 28) <= 5; angryBirdLarge(92, 29) <= 5; angryBirdLarge(92, 30) <= 4; angryBirdLarge(92, 31) <= 4; angryBirdLarge(92, 32) <= 4; angryBirdLarge(92, 33) <= 4; angryBirdLarge(92, 34) <= 4; angryBirdLarge(92, 35) <= 4; angryBirdLarge(92, 36) <= 4; angryBirdLarge(92, 37) <= 4; angryBirdLarge(92, 38) <= 4; angryBirdLarge(92, 39) <= 4; angryBirdLarge(92, 40) <= 4; angryBirdLarge(92, 41) <= 4; angryBirdLarge(92, 42) <= 4; angryBirdLarge(92, 43) <= 4; angryBirdLarge(92, 44) <= 4; angryBirdLarge(92, 45) <= 4; angryBirdLarge(92, 46) <= 4; angryBirdLarge(92, 47) <= 4; angryBirdLarge(92, 48) <= 4; angryBirdLarge(92, 49) <= 4; angryBirdLarge(92, 50) <= 4; angryBirdLarge(92, 51) <= 4; angryBirdLarge(92, 52) <= 4; angryBirdLarge(92, 53) <= 4; angryBirdLarge(92, 54) <= 4; angryBirdLarge(92, 55) <= 4; angryBirdLarge(92, 56) <= 4; angryBirdLarge(92, 57) <= 4; angryBirdLarge(92, 58) <= 4; angryBirdLarge(92, 59) <= 4; angryBirdLarge(92, 60) <= 4; angryBirdLarge(92, 61) <= 4; angryBirdLarge(92, 62) <= 4; angryBirdLarge(92, 63) <= 4; angryBirdLarge(92, 64) <= 4; angryBirdLarge(92, 65) <= 4; angryBirdLarge(92, 66) <= 4; angryBirdLarge(92, 67) <= 4; angryBirdLarge(92, 68) <= 4; angryBirdLarge(92, 69) <= 4; angryBirdLarge(92, 70) <= 4; angryBirdLarge(92, 71) <= 4; angryBirdLarge(92, 72) <= 4; angryBirdLarge(92, 73) <= 4; angryBirdLarge(92, 74) <= 4; angryBirdLarge(92, 75) <= 4; angryBirdLarge(92, 76) <= 4; angryBirdLarge(92, 77) <= 4; angryBirdLarge(92, 78) <= 4; angryBirdLarge(92, 79) <= 4; angryBirdLarge(92, 80) <= 4; angryBirdLarge(92, 81) <= 4; angryBirdLarge(92, 82) <= 4; angryBirdLarge(92, 83) <= 4; angryBirdLarge(92, 84) <= 4; angryBirdLarge(92, 85) <= 4; angryBirdLarge(92, 86) <= 4; angryBirdLarge(92, 87) <= 4; angryBirdLarge(92, 88) <= 4; angryBirdLarge(92, 89) <= 4; angryBirdLarge(92, 90) <= 5; angryBirdLarge(92, 91) <= 5; angryBirdLarge(92, 92) <= 5; angryBirdLarge(92, 93) <= 5; angryBirdLarge(92, 94) <= 5; angryBirdLarge(92, 95) <= 5; angryBirdLarge(92, 96) <= 5; angryBirdLarge(92, 97) <= 5; angryBirdLarge(92, 98) <= 5; angryBirdLarge(92, 99) <= 5; angryBirdLarge(92, 100) <= 5; angryBirdLarge(92, 101) <= 5; angryBirdLarge(92, 102) <= 3; angryBirdLarge(92, 103) <= 3; angryBirdLarge(92, 104) <= 3; angryBirdLarge(92, 105) <= 3; angryBirdLarge(92, 106) <= 3; angryBirdLarge(92, 107) <= 3; angryBirdLarge(92, 108) <= 3; angryBirdLarge(92, 109) <= 3; angryBirdLarge(92, 110) <= 3; angryBirdLarge(92, 111) <= 3; angryBirdLarge(92, 112) <= 3; angryBirdLarge(92, 113) <= 3; angryBirdLarge(92, 114) <= 3; angryBirdLarge(92, 115) <= 3; angryBirdLarge(92, 116) <= 3; angryBirdLarge(92, 117) <= 3; angryBirdLarge(92, 118) <= 3; angryBirdLarge(92, 119) <= 3; angryBirdLarge(92, 120) <= 5; angryBirdLarge(92, 121) <= 5; angryBirdLarge(92, 122) <= 5; angryBirdLarge(92, 123) <= 5; angryBirdLarge(92, 124) <= 5; angryBirdLarge(92, 125) <= 5; angryBirdLarge(92, 126) <= 5; angryBirdLarge(92, 127) <= 5; angryBirdLarge(92, 128) <= 5; angryBirdLarge(92, 129) <= 5; angryBirdLarge(92, 130) <= 5; angryBirdLarge(92, 131) <= 5; angryBirdLarge(92, 132) <= 4; angryBirdLarge(92, 133) <= 4; angryBirdLarge(92, 134) <= 4; angryBirdLarge(92, 135) <= 4; angryBirdLarge(92, 136) <= 4; angryBirdLarge(92, 137) <= 4; angryBirdLarge(92, 138) <= 4; angryBirdLarge(92, 139) <= 4; angryBirdLarge(92, 140) <= 4; angryBirdLarge(92, 141) <= 4; angryBirdLarge(92, 142) <= 4; angryBirdLarge(92, 143) <= 4; angryBirdLarge(92, 144) <= 5; angryBirdLarge(92, 145) <= 5; angryBirdLarge(92, 146) <= 5; angryBirdLarge(92, 147) <= 5; angryBirdLarge(92, 148) <= 5; angryBirdLarge(92, 149) <= 5; 
angryBirdLarge(93, 0) <= 0; angryBirdLarge(93, 1) <= 0; angryBirdLarge(93, 2) <= 0; angryBirdLarge(93, 3) <= 0; angryBirdLarge(93, 4) <= 0; angryBirdLarge(93, 5) <= 0; angryBirdLarge(93, 6) <= 0; angryBirdLarge(93, 7) <= 0; angryBirdLarge(93, 8) <= 0; angryBirdLarge(93, 9) <= 0; angryBirdLarge(93, 10) <= 0; angryBirdLarge(93, 11) <= 0; angryBirdLarge(93, 12) <= 0; angryBirdLarge(93, 13) <= 0; angryBirdLarge(93, 14) <= 0; angryBirdLarge(93, 15) <= 0; angryBirdLarge(93, 16) <= 0; angryBirdLarge(93, 17) <= 0; angryBirdLarge(93, 18) <= 5; angryBirdLarge(93, 19) <= 5; angryBirdLarge(93, 20) <= 5; angryBirdLarge(93, 21) <= 5; angryBirdLarge(93, 22) <= 5; angryBirdLarge(93, 23) <= 5; angryBirdLarge(93, 24) <= 5; angryBirdLarge(93, 25) <= 5; angryBirdLarge(93, 26) <= 5; angryBirdLarge(93, 27) <= 5; angryBirdLarge(93, 28) <= 5; angryBirdLarge(93, 29) <= 5; angryBirdLarge(93, 30) <= 4; angryBirdLarge(93, 31) <= 4; angryBirdLarge(93, 32) <= 4; angryBirdLarge(93, 33) <= 4; angryBirdLarge(93, 34) <= 4; angryBirdLarge(93, 35) <= 4; angryBirdLarge(93, 36) <= 4; angryBirdLarge(93, 37) <= 4; angryBirdLarge(93, 38) <= 4; angryBirdLarge(93, 39) <= 4; angryBirdLarge(93, 40) <= 4; angryBirdLarge(93, 41) <= 4; angryBirdLarge(93, 42) <= 4; angryBirdLarge(93, 43) <= 4; angryBirdLarge(93, 44) <= 4; angryBirdLarge(93, 45) <= 4; angryBirdLarge(93, 46) <= 4; angryBirdLarge(93, 47) <= 4; angryBirdLarge(93, 48) <= 4; angryBirdLarge(93, 49) <= 4; angryBirdLarge(93, 50) <= 4; angryBirdLarge(93, 51) <= 4; angryBirdLarge(93, 52) <= 4; angryBirdLarge(93, 53) <= 4; angryBirdLarge(93, 54) <= 4; angryBirdLarge(93, 55) <= 4; angryBirdLarge(93, 56) <= 4; angryBirdLarge(93, 57) <= 4; angryBirdLarge(93, 58) <= 4; angryBirdLarge(93, 59) <= 4; angryBirdLarge(93, 60) <= 4; angryBirdLarge(93, 61) <= 4; angryBirdLarge(93, 62) <= 4; angryBirdLarge(93, 63) <= 4; angryBirdLarge(93, 64) <= 4; angryBirdLarge(93, 65) <= 4; angryBirdLarge(93, 66) <= 4; angryBirdLarge(93, 67) <= 4; angryBirdLarge(93, 68) <= 4; angryBirdLarge(93, 69) <= 4; angryBirdLarge(93, 70) <= 4; angryBirdLarge(93, 71) <= 4; angryBirdLarge(93, 72) <= 4; angryBirdLarge(93, 73) <= 4; angryBirdLarge(93, 74) <= 4; angryBirdLarge(93, 75) <= 4; angryBirdLarge(93, 76) <= 4; angryBirdLarge(93, 77) <= 4; angryBirdLarge(93, 78) <= 4; angryBirdLarge(93, 79) <= 4; angryBirdLarge(93, 80) <= 4; angryBirdLarge(93, 81) <= 4; angryBirdLarge(93, 82) <= 4; angryBirdLarge(93, 83) <= 4; angryBirdLarge(93, 84) <= 4; angryBirdLarge(93, 85) <= 4; angryBirdLarge(93, 86) <= 4; angryBirdLarge(93, 87) <= 4; angryBirdLarge(93, 88) <= 4; angryBirdLarge(93, 89) <= 4; angryBirdLarge(93, 90) <= 5; angryBirdLarge(93, 91) <= 5; angryBirdLarge(93, 92) <= 5; angryBirdLarge(93, 93) <= 5; angryBirdLarge(93, 94) <= 5; angryBirdLarge(93, 95) <= 5; angryBirdLarge(93, 96) <= 5; angryBirdLarge(93, 97) <= 5; angryBirdLarge(93, 98) <= 5; angryBirdLarge(93, 99) <= 5; angryBirdLarge(93, 100) <= 5; angryBirdLarge(93, 101) <= 5; angryBirdLarge(93, 102) <= 3; angryBirdLarge(93, 103) <= 3; angryBirdLarge(93, 104) <= 3; angryBirdLarge(93, 105) <= 3; angryBirdLarge(93, 106) <= 3; angryBirdLarge(93, 107) <= 3; angryBirdLarge(93, 108) <= 3; angryBirdLarge(93, 109) <= 3; angryBirdLarge(93, 110) <= 3; angryBirdLarge(93, 111) <= 3; angryBirdLarge(93, 112) <= 3; angryBirdLarge(93, 113) <= 3; angryBirdLarge(93, 114) <= 3; angryBirdLarge(93, 115) <= 3; angryBirdLarge(93, 116) <= 3; angryBirdLarge(93, 117) <= 3; angryBirdLarge(93, 118) <= 3; angryBirdLarge(93, 119) <= 3; angryBirdLarge(93, 120) <= 5; angryBirdLarge(93, 121) <= 5; angryBirdLarge(93, 122) <= 5; angryBirdLarge(93, 123) <= 5; angryBirdLarge(93, 124) <= 5; angryBirdLarge(93, 125) <= 5; angryBirdLarge(93, 126) <= 5; angryBirdLarge(93, 127) <= 5; angryBirdLarge(93, 128) <= 5; angryBirdLarge(93, 129) <= 5; angryBirdLarge(93, 130) <= 5; angryBirdLarge(93, 131) <= 5; angryBirdLarge(93, 132) <= 4; angryBirdLarge(93, 133) <= 4; angryBirdLarge(93, 134) <= 4; angryBirdLarge(93, 135) <= 4; angryBirdLarge(93, 136) <= 4; angryBirdLarge(93, 137) <= 4; angryBirdLarge(93, 138) <= 4; angryBirdLarge(93, 139) <= 4; angryBirdLarge(93, 140) <= 4; angryBirdLarge(93, 141) <= 4; angryBirdLarge(93, 142) <= 4; angryBirdLarge(93, 143) <= 4; angryBirdLarge(93, 144) <= 5; angryBirdLarge(93, 145) <= 5; angryBirdLarge(93, 146) <= 5; angryBirdLarge(93, 147) <= 5; angryBirdLarge(93, 148) <= 5; angryBirdLarge(93, 149) <= 5; 
angryBirdLarge(94, 0) <= 0; angryBirdLarge(94, 1) <= 0; angryBirdLarge(94, 2) <= 0; angryBirdLarge(94, 3) <= 0; angryBirdLarge(94, 4) <= 0; angryBirdLarge(94, 5) <= 0; angryBirdLarge(94, 6) <= 0; angryBirdLarge(94, 7) <= 0; angryBirdLarge(94, 8) <= 0; angryBirdLarge(94, 9) <= 0; angryBirdLarge(94, 10) <= 0; angryBirdLarge(94, 11) <= 0; angryBirdLarge(94, 12) <= 0; angryBirdLarge(94, 13) <= 0; angryBirdLarge(94, 14) <= 0; angryBirdLarge(94, 15) <= 0; angryBirdLarge(94, 16) <= 0; angryBirdLarge(94, 17) <= 0; angryBirdLarge(94, 18) <= 5; angryBirdLarge(94, 19) <= 5; angryBirdLarge(94, 20) <= 5; angryBirdLarge(94, 21) <= 5; angryBirdLarge(94, 22) <= 5; angryBirdLarge(94, 23) <= 5; angryBirdLarge(94, 24) <= 5; angryBirdLarge(94, 25) <= 5; angryBirdLarge(94, 26) <= 5; angryBirdLarge(94, 27) <= 5; angryBirdLarge(94, 28) <= 5; angryBirdLarge(94, 29) <= 5; angryBirdLarge(94, 30) <= 4; angryBirdLarge(94, 31) <= 4; angryBirdLarge(94, 32) <= 4; angryBirdLarge(94, 33) <= 4; angryBirdLarge(94, 34) <= 4; angryBirdLarge(94, 35) <= 4; angryBirdLarge(94, 36) <= 4; angryBirdLarge(94, 37) <= 4; angryBirdLarge(94, 38) <= 4; angryBirdLarge(94, 39) <= 4; angryBirdLarge(94, 40) <= 4; angryBirdLarge(94, 41) <= 4; angryBirdLarge(94, 42) <= 4; angryBirdLarge(94, 43) <= 4; angryBirdLarge(94, 44) <= 4; angryBirdLarge(94, 45) <= 4; angryBirdLarge(94, 46) <= 4; angryBirdLarge(94, 47) <= 4; angryBirdLarge(94, 48) <= 4; angryBirdLarge(94, 49) <= 4; angryBirdLarge(94, 50) <= 4; angryBirdLarge(94, 51) <= 4; angryBirdLarge(94, 52) <= 4; angryBirdLarge(94, 53) <= 4; angryBirdLarge(94, 54) <= 4; angryBirdLarge(94, 55) <= 4; angryBirdLarge(94, 56) <= 4; angryBirdLarge(94, 57) <= 4; angryBirdLarge(94, 58) <= 4; angryBirdLarge(94, 59) <= 4; angryBirdLarge(94, 60) <= 4; angryBirdLarge(94, 61) <= 4; angryBirdLarge(94, 62) <= 4; angryBirdLarge(94, 63) <= 4; angryBirdLarge(94, 64) <= 4; angryBirdLarge(94, 65) <= 4; angryBirdLarge(94, 66) <= 4; angryBirdLarge(94, 67) <= 4; angryBirdLarge(94, 68) <= 4; angryBirdLarge(94, 69) <= 4; angryBirdLarge(94, 70) <= 4; angryBirdLarge(94, 71) <= 4; angryBirdLarge(94, 72) <= 4; angryBirdLarge(94, 73) <= 4; angryBirdLarge(94, 74) <= 4; angryBirdLarge(94, 75) <= 4; angryBirdLarge(94, 76) <= 4; angryBirdLarge(94, 77) <= 4; angryBirdLarge(94, 78) <= 4; angryBirdLarge(94, 79) <= 4; angryBirdLarge(94, 80) <= 4; angryBirdLarge(94, 81) <= 4; angryBirdLarge(94, 82) <= 4; angryBirdLarge(94, 83) <= 4; angryBirdLarge(94, 84) <= 4; angryBirdLarge(94, 85) <= 4; angryBirdLarge(94, 86) <= 4; angryBirdLarge(94, 87) <= 4; angryBirdLarge(94, 88) <= 4; angryBirdLarge(94, 89) <= 4; angryBirdLarge(94, 90) <= 5; angryBirdLarge(94, 91) <= 5; angryBirdLarge(94, 92) <= 5; angryBirdLarge(94, 93) <= 5; angryBirdLarge(94, 94) <= 5; angryBirdLarge(94, 95) <= 5; angryBirdLarge(94, 96) <= 5; angryBirdLarge(94, 97) <= 5; angryBirdLarge(94, 98) <= 5; angryBirdLarge(94, 99) <= 5; angryBirdLarge(94, 100) <= 5; angryBirdLarge(94, 101) <= 5; angryBirdLarge(94, 102) <= 3; angryBirdLarge(94, 103) <= 3; angryBirdLarge(94, 104) <= 3; angryBirdLarge(94, 105) <= 3; angryBirdLarge(94, 106) <= 3; angryBirdLarge(94, 107) <= 3; angryBirdLarge(94, 108) <= 3; angryBirdLarge(94, 109) <= 3; angryBirdLarge(94, 110) <= 3; angryBirdLarge(94, 111) <= 3; angryBirdLarge(94, 112) <= 3; angryBirdLarge(94, 113) <= 3; angryBirdLarge(94, 114) <= 3; angryBirdLarge(94, 115) <= 3; angryBirdLarge(94, 116) <= 3; angryBirdLarge(94, 117) <= 3; angryBirdLarge(94, 118) <= 3; angryBirdLarge(94, 119) <= 3; angryBirdLarge(94, 120) <= 5; angryBirdLarge(94, 121) <= 5; angryBirdLarge(94, 122) <= 5; angryBirdLarge(94, 123) <= 5; angryBirdLarge(94, 124) <= 5; angryBirdLarge(94, 125) <= 5; angryBirdLarge(94, 126) <= 5; angryBirdLarge(94, 127) <= 5; angryBirdLarge(94, 128) <= 5; angryBirdLarge(94, 129) <= 5; angryBirdLarge(94, 130) <= 5; angryBirdLarge(94, 131) <= 5; angryBirdLarge(94, 132) <= 4; angryBirdLarge(94, 133) <= 4; angryBirdLarge(94, 134) <= 4; angryBirdLarge(94, 135) <= 4; angryBirdLarge(94, 136) <= 4; angryBirdLarge(94, 137) <= 4; angryBirdLarge(94, 138) <= 4; angryBirdLarge(94, 139) <= 4; angryBirdLarge(94, 140) <= 4; angryBirdLarge(94, 141) <= 4; angryBirdLarge(94, 142) <= 4; angryBirdLarge(94, 143) <= 4; angryBirdLarge(94, 144) <= 5; angryBirdLarge(94, 145) <= 5; angryBirdLarge(94, 146) <= 5; angryBirdLarge(94, 147) <= 5; angryBirdLarge(94, 148) <= 5; angryBirdLarge(94, 149) <= 5; 
angryBirdLarge(95, 0) <= 0; angryBirdLarge(95, 1) <= 0; angryBirdLarge(95, 2) <= 0; angryBirdLarge(95, 3) <= 0; angryBirdLarge(95, 4) <= 0; angryBirdLarge(95, 5) <= 0; angryBirdLarge(95, 6) <= 0; angryBirdLarge(95, 7) <= 0; angryBirdLarge(95, 8) <= 0; angryBirdLarge(95, 9) <= 0; angryBirdLarge(95, 10) <= 0; angryBirdLarge(95, 11) <= 0; angryBirdLarge(95, 12) <= 0; angryBirdLarge(95, 13) <= 0; angryBirdLarge(95, 14) <= 0; angryBirdLarge(95, 15) <= 0; angryBirdLarge(95, 16) <= 0; angryBirdLarge(95, 17) <= 0; angryBirdLarge(95, 18) <= 5; angryBirdLarge(95, 19) <= 5; angryBirdLarge(95, 20) <= 5; angryBirdLarge(95, 21) <= 5; angryBirdLarge(95, 22) <= 5; angryBirdLarge(95, 23) <= 5; angryBirdLarge(95, 24) <= 5; angryBirdLarge(95, 25) <= 5; angryBirdLarge(95, 26) <= 5; angryBirdLarge(95, 27) <= 5; angryBirdLarge(95, 28) <= 5; angryBirdLarge(95, 29) <= 5; angryBirdLarge(95, 30) <= 4; angryBirdLarge(95, 31) <= 4; angryBirdLarge(95, 32) <= 4; angryBirdLarge(95, 33) <= 4; angryBirdLarge(95, 34) <= 4; angryBirdLarge(95, 35) <= 4; angryBirdLarge(95, 36) <= 4; angryBirdLarge(95, 37) <= 4; angryBirdLarge(95, 38) <= 4; angryBirdLarge(95, 39) <= 4; angryBirdLarge(95, 40) <= 4; angryBirdLarge(95, 41) <= 4; angryBirdLarge(95, 42) <= 4; angryBirdLarge(95, 43) <= 4; angryBirdLarge(95, 44) <= 4; angryBirdLarge(95, 45) <= 4; angryBirdLarge(95, 46) <= 4; angryBirdLarge(95, 47) <= 4; angryBirdLarge(95, 48) <= 4; angryBirdLarge(95, 49) <= 4; angryBirdLarge(95, 50) <= 4; angryBirdLarge(95, 51) <= 4; angryBirdLarge(95, 52) <= 4; angryBirdLarge(95, 53) <= 4; angryBirdLarge(95, 54) <= 4; angryBirdLarge(95, 55) <= 4; angryBirdLarge(95, 56) <= 4; angryBirdLarge(95, 57) <= 4; angryBirdLarge(95, 58) <= 4; angryBirdLarge(95, 59) <= 4; angryBirdLarge(95, 60) <= 4; angryBirdLarge(95, 61) <= 4; angryBirdLarge(95, 62) <= 4; angryBirdLarge(95, 63) <= 4; angryBirdLarge(95, 64) <= 4; angryBirdLarge(95, 65) <= 4; angryBirdLarge(95, 66) <= 4; angryBirdLarge(95, 67) <= 4; angryBirdLarge(95, 68) <= 4; angryBirdLarge(95, 69) <= 4; angryBirdLarge(95, 70) <= 4; angryBirdLarge(95, 71) <= 4; angryBirdLarge(95, 72) <= 4; angryBirdLarge(95, 73) <= 4; angryBirdLarge(95, 74) <= 4; angryBirdLarge(95, 75) <= 4; angryBirdLarge(95, 76) <= 4; angryBirdLarge(95, 77) <= 4; angryBirdLarge(95, 78) <= 4; angryBirdLarge(95, 79) <= 4; angryBirdLarge(95, 80) <= 4; angryBirdLarge(95, 81) <= 4; angryBirdLarge(95, 82) <= 4; angryBirdLarge(95, 83) <= 4; angryBirdLarge(95, 84) <= 4; angryBirdLarge(95, 85) <= 4; angryBirdLarge(95, 86) <= 4; angryBirdLarge(95, 87) <= 4; angryBirdLarge(95, 88) <= 4; angryBirdLarge(95, 89) <= 4; angryBirdLarge(95, 90) <= 5; angryBirdLarge(95, 91) <= 5; angryBirdLarge(95, 92) <= 5; angryBirdLarge(95, 93) <= 5; angryBirdLarge(95, 94) <= 5; angryBirdLarge(95, 95) <= 5; angryBirdLarge(95, 96) <= 5; angryBirdLarge(95, 97) <= 5; angryBirdLarge(95, 98) <= 5; angryBirdLarge(95, 99) <= 5; angryBirdLarge(95, 100) <= 5; angryBirdLarge(95, 101) <= 5; angryBirdLarge(95, 102) <= 3; angryBirdLarge(95, 103) <= 3; angryBirdLarge(95, 104) <= 3; angryBirdLarge(95, 105) <= 3; angryBirdLarge(95, 106) <= 3; angryBirdLarge(95, 107) <= 3; angryBirdLarge(95, 108) <= 3; angryBirdLarge(95, 109) <= 3; angryBirdLarge(95, 110) <= 3; angryBirdLarge(95, 111) <= 3; angryBirdLarge(95, 112) <= 3; angryBirdLarge(95, 113) <= 3; angryBirdLarge(95, 114) <= 3; angryBirdLarge(95, 115) <= 3; angryBirdLarge(95, 116) <= 3; angryBirdLarge(95, 117) <= 3; angryBirdLarge(95, 118) <= 3; angryBirdLarge(95, 119) <= 3; angryBirdLarge(95, 120) <= 5; angryBirdLarge(95, 121) <= 5; angryBirdLarge(95, 122) <= 5; angryBirdLarge(95, 123) <= 5; angryBirdLarge(95, 124) <= 5; angryBirdLarge(95, 125) <= 5; angryBirdLarge(95, 126) <= 5; angryBirdLarge(95, 127) <= 5; angryBirdLarge(95, 128) <= 5; angryBirdLarge(95, 129) <= 5; angryBirdLarge(95, 130) <= 5; angryBirdLarge(95, 131) <= 5; angryBirdLarge(95, 132) <= 4; angryBirdLarge(95, 133) <= 4; angryBirdLarge(95, 134) <= 4; angryBirdLarge(95, 135) <= 4; angryBirdLarge(95, 136) <= 4; angryBirdLarge(95, 137) <= 4; angryBirdLarge(95, 138) <= 4; angryBirdLarge(95, 139) <= 4; angryBirdLarge(95, 140) <= 4; angryBirdLarge(95, 141) <= 4; angryBirdLarge(95, 142) <= 4; angryBirdLarge(95, 143) <= 4; angryBirdLarge(95, 144) <= 5; angryBirdLarge(95, 145) <= 5; angryBirdLarge(95, 146) <= 5; angryBirdLarge(95, 147) <= 5; angryBirdLarge(95, 148) <= 5; angryBirdLarge(95, 149) <= 5; 
angryBirdLarge(96, 0) <= 0; angryBirdLarge(96, 1) <= 0; angryBirdLarge(96, 2) <= 0; angryBirdLarge(96, 3) <= 0; angryBirdLarge(96, 4) <= 0; angryBirdLarge(96, 5) <= 0; angryBirdLarge(96, 6) <= 5; angryBirdLarge(96, 7) <= 5; angryBirdLarge(96, 8) <= 5; angryBirdLarge(96, 9) <= 5; angryBirdLarge(96, 10) <= 5; angryBirdLarge(96, 11) <= 5; angryBirdLarge(96, 12) <= 5; angryBirdLarge(96, 13) <= 5; angryBirdLarge(96, 14) <= 5; angryBirdLarge(96, 15) <= 5; angryBirdLarge(96, 16) <= 5; angryBirdLarge(96, 17) <= 5; angryBirdLarge(96, 18) <= 0; angryBirdLarge(96, 19) <= 0; angryBirdLarge(96, 20) <= 0; angryBirdLarge(96, 21) <= 0; angryBirdLarge(96, 22) <= 0; angryBirdLarge(96, 23) <= 0; angryBirdLarge(96, 24) <= 4; angryBirdLarge(96, 25) <= 4; angryBirdLarge(96, 26) <= 4; angryBirdLarge(96, 27) <= 4; angryBirdLarge(96, 28) <= 4; angryBirdLarge(96, 29) <= 4; angryBirdLarge(96, 30) <= 4; angryBirdLarge(96, 31) <= 4; angryBirdLarge(96, 32) <= 4; angryBirdLarge(96, 33) <= 4; angryBirdLarge(96, 34) <= 4; angryBirdLarge(96, 35) <= 4; angryBirdLarge(96, 36) <= 4; angryBirdLarge(96, 37) <= 4; angryBirdLarge(96, 38) <= 4; angryBirdLarge(96, 39) <= 4; angryBirdLarge(96, 40) <= 4; angryBirdLarge(96, 41) <= 4; angryBirdLarge(96, 42) <= 4; angryBirdLarge(96, 43) <= 4; angryBirdLarge(96, 44) <= 4; angryBirdLarge(96, 45) <= 4; angryBirdLarge(96, 46) <= 4; angryBirdLarge(96, 47) <= 4; angryBirdLarge(96, 48) <= 4; angryBirdLarge(96, 49) <= 4; angryBirdLarge(96, 50) <= 4; angryBirdLarge(96, 51) <= 4; angryBirdLarge(96, 52) <= 4; angryBirdLarge(96, 53) <= 4; angryBirdLarge(96, 54) <= 4; angryBirdLarge(96, 55) <= 4; angryBirdLarge(96, 56) <= 4; angryBirdLarge(96, 57) <= 4; angryBirdLarge(96, 58) <= 4; angryBirdLarge(96, 59) <= 4; angryBirdLarge(96, 60) <= 4; angryBirdLarge(96, 61) <= 4; angryBirdLarge(96, 62) <= 4; angryBirdLarge(96, 63) <= 4; angryBirdLarge(96, 64) <= 4; angryBirdLarge(96, 65) <= 4; angryBirdLarge(96, 66) <= 4; angryBirdLarge(96, 67) <= 4; angryBirdLarge(96, 68) <= 4; angryBirdLarge(96, 69) <= 4; angryBirdLarge(96, 70) <= 4; angryBirdLarge(96, 71) <= 4; angryBirdLarge(96, 72) <= 4; angryBirdLarge(96, 73) <= 4; angryBirdLarge(96, 74) <= 4; angryBirdLarge(96, 75) <= 4; angryBirdLarge(96, 76) <= 4; angryBirdLarge(96, 77) <= 4; angryBirdLarge(96, 78) <= 4; angryBirdLarge(96, 79) <= 4; angryBirdLarge(96, 80) <= 4; angryBirdLarge(96, 81) <= 4; angryBirdLarge(96, 82) <= 4; angryBirdLarge(96, 83) <= 4; angryBirdLarge(96, 84) <= 4; angryBirdLarge(96, 85) <= 4; angryBirdLarge(96, 86) <= 4; angryBirdLarge(96, 87) <= 4; angryBirdLarge(96, 88) <= 4; angryBirdLarge(96, 89) <= 4; angryBirdLarge(96, 90) <= 5; angryBirdLarge(96, 91) <= 5; angryBirdLarge(96, 92) <= 5; angryBirdLarge(96, 93) <= 5; angryBirdLarge(96, 94) <= 5; angryBirdLarge(96, 95) <= 5; angryBirdLarge(96, 96) <= 3; angryBirdLarge(96, 97) <= 3; angryBirdLarge(96, 98) <= 3; angryBirdLarge(96, 99) <= 3; angryBirdLarge(96, 100) <= 3; angryBirdLarge(96, 101) <= 3; angryBirdLarge(96, 102) <= 3; angryBirdLarge(96, 103) <= 3; angryBirdLarge(96, 104) <= 3; angryBirdLarge(96, 105) <= 3; angryBirdLarge(96, 106) <= 3; angryBirdLarge(96, 107) <= 3; angryBirdLarge(96, 108) <= 3; angryBirdLarge(96, 109) <= 3; angryBirdLarge(96, 110) <= 3; angryBirdLarge(96, 111) <= 3; angryBirdLarge(96, 112) <= 3; angryBirdLarge(96, 113) <= 3; angryBirdLarge(96, 114) <= 3; angryBirdLarge(96, 115) <= 3; angryBirdLarge(96, 116) <= 3; angryBirdLarge(96, 117) <= 3; angryBirdLarge(96, 118) <= 3; angryBirdLarge(96, 119) <= 3; angryBirdLarge(96, 120) <= 3; angryBirdLarge(96, 121) <= 3; angryBirdLarge(96, 122) <= 3; angryBirdLarge(96, 123) <= 3; angryBirdLarge(96, 124) <= 3; angryBirdLarge(96, 125) <= 3; angryBirdLarge(96, 126) <= 3; angryBirdLarge(96, 127) <= 3; angryBirdLarge(96, 128) <= 3; angryBirdLarge(96, 129) <= 3; angryBirdLarge(96, 130) <= 3; angryBirdLarge(96, 131) <= 3; angryBirdLarge(96, 132) <= 5; angryBirdLarge(96, 133) <= 5; angryBirdLarge(96, 134) <= 5; angryBirdLarge(96, 135) <= 5; angryBirdLarge(96, 136) <= 5; angryBirdLarge(96, 137) <= 5; angryBirdLarge(96, 138) <= 4; angryBirdLarge(96, 139) <= 4; angryBirdLarge(96, 140) <= 4; angryBirdLarge(96, 141) <= 4; angryBirdLarge(96, 142) <= 4; angryBirdLarge(96, 143) <= 4; angryBirdLarge(96, 144) <= 5; angryBirdLarge(96, 145) <= 5; angryBirdLarge(96, 146) <= 5; angryBirdLarge(96, 147) <= 5; angryBirdLarge(96, 148) <= 5; angryBirdLarge(96, 149) <= 5; 
angryBirdLarge(97, 0) <= 0; angryBirdLarge(97, 1) <= 0; angryBirdLarge(97, 2) <= 0; angryBirdLarge(97, 3) <= 0; angryBirdLarge(97, 4) <= 0; angryBirdLarge(97, 5) <= 0; angryBirdLarge(97, 6) <= 5; angryBirdLarge(97, 7) <= 5; angryBirdLarge(97, 8) <= 5; angryBirdLarge(97, 9) <= 5; angryBirdLarge(97, 10) <= 5; angryBirdLarge(97, 11) <= 5; angryBirdLarge(97, 12) <= 5; angryBirdLarge(97, 13) <= 5; angryBirdLarge(97, 14) <= 5; angryBirdLarge(97, 15) <= 5; angryBirdLarge(97, 16) <= 5; angryBirdLarge(97, 17) <= 5; angryBirdLarge(97, 18) <= 0; angryBirdLarge(97, 19) <= 0; angryBirdLarge(97, 20) <= 0; angryBirdLarge(97, 21) <= 0; angryBirdLarge(97, 22) <= 0; angryBirdLarge(97, 23) <= 0; angryBirdLarge(97, 24) <= 4; angryBirdLarge(97, 25) <= 4; angryBirdLarge(97, 26) <= 4; angryBirdLarge(97, 27) <= 4; angryBirdLarge(97, 28) <= 4; angryBirdLarge(97, 29) <= 4; angryBirdLarge(97, 30) <= 4; angryBirdLarge(97, 31) <= 4; angryBirdLarge(97, 32) <= 4; angryBirdLarge(97, 33) <= 4; angryBirdLarge(97, 34) <= 4; angryBirdLarge(97, 35) <= 4; angryBirdLarge(97, 36) <= 4; angryBirdLarge(97, 37) <= 4; angryBirdLarge(97, 38) <= 4; angryBirdLarge(97, 39) <= 4; angryBirdLarge(97, 40) <= 4; angryBirdLarge(97, 41) <= 4; angryBirdLarge(97, 42) <= 4; angryBirdLarge(97, 43) <= 4; angryBirdLarge(97, 44) <= 4; angryBirdLarge(97, 45) <= 4; angryBirdLarge(97, 46) <= 4; angryBirdLarge(97, 47) <= 4; angryBirdLarge(97, 48) <= 4; angryBirdLarge(97, 49) <= 4; angryBirdLarge(97, 50) <= 4; angryBirdLarge(97, 51) <= 4; angryBirdLarge(97, 52) <= 4; angryBirdLarge(97, 53) <= 4; angryBirdLarge(97, 54) <= 4; angryBirdLarge(97, 55) <= 4; angryBirdLarge(97, 56) <= 4; angryBirdLarge(97, 57) <= 4; angryBirdLarge(97, 58) <= 4; angryBirdLarge(97, 59) <= 4; angryBirdLarge(97, 60) <= 4; angryBirdLarge(97, 61) <= 4; angryBirdLarge(97, 62) <= 4; angryBirdLarge(97, 63) <= 4; angryBirdLarge(97, 64) <= 4; angryBirdLarge(97, 65) <= 4; angryBirdLarge(97, 66) <= 4; angryBirdLarge(97, 67) <= 4; angryBirdLarge(97, 68) <= 4; angryBirdLarge(97, 69) <= 4; angryBirdLarge(97, 70) <= 4; angryBirdLarge(97, 71) <= 4; angryBirdLarge(97, 72) <= 4; angryBirdLarge(97, 73) <= 4; angryBirdLarge(97, 74) <= 4; angryBirdLarge(97, 75) <= 4; angryBirdLarge(97, 76) <= 4; angryBirdLarge(97, 77) <= 4; angryBirdLarge(97, 78) <= 4; angryBirdLarge(97, 79) <= 4; angryBirdLarge(97, 80) <= 4; angryBirdLarge(97, 81) <= 4; angryBirdLarge(97, 82) <= 4; angryBirdLarge(97, 83) <= 4; angryBirdLarge(97, 84) <= 4; angryBirdLarge(97, 85) <= 4; angryBirdLarge(97, 86) <= 4; angryBirdLarge(97, 87) <= 4; angryBirdLarge(97, 88) <= 4; angryBirdLarge(97, 89) <= 4; angryBirdLarge(97, 90) <= 5; angryBirdLarge(97, 91) <= 5; angryBirdLarge(97, 92) <= 5; angryBirdLarge(97, 93) <= 5; angryBirdLarge(97, 94) <= 5; angryBirdLarge(97, 95) <= 5; angryBirdLarge(97, 96) <= 3; angryBirdLarge(97, 97) <= 3; angryBirdLarge(97, 98) <= 3; angryBirdLarge(97, 99) <= 3; angryBirdLarge(97, 100) <= 3; angryBirdLarge(97, 101) <= 3; angryBirdLarge(97, 102) <= 3; angryBirdLarge(97, 103) <= 3; angryBirdLarge(97, 104) <= 3; angryBirdLarge(97, 105) <= 3; angryBirdLarge(97, 106) <= 3; angryBirdLarge(97, 107) <= 3; angryBirdLarge(97, 108) <= 3; angryBirdLarge(97, 109) <= 3; angryBirdLarge(97, 110) <= 3; angryBirdLarge(97, 111) <= 3; angryBirdLarge(97, 112) <= 3; angryBirdLarge(97, 113) <= 3; angryBirdLarge(97, 114) <= 3; angryBirdLarge(97, 115) <= 3; angryBirdLarge(97, 116) <= 3; angryBirdLarge(97, 117) <= 3; angryBirdLarge(97, 118) <= 3; angryBirdLarge(97, 119) <= 3; angryBirdLarge(97, 120) <= 3; angryBirdLarge(97, 121) <= 3; angryBirdLarge(97, 122) <= 3; angryBirdLarge(97, 123) <= 3; angryBirdLarge(97, 124) <= 3; angryBirdLarge(97, 125) <= 3; angryBirdLarge(97, 126) <= 3; angryBirdLarge(97, 127) <= 3; angryBirdLarge(97, 128) <= 3; angryBirdLarge(97, 129) <= 3; angryBirdLarge(97, 130) <= 3; angryBirdLarge(97, 131) <= 3; angryBirdLarge(97, 132) <= 5; angryBirdLarge(97, 133) <= 5; angryBirdLarge(97, 134) <= 5; angryBirdLarge(97, 135) <= 5; angryBirdLarge(97, 136) <= 5; angryBirdLarge(97, 137) <= 5; angryBirdLarge(97, 138) <= 4; angryBirdLarge(97, 139) <= 4; angryBirdLarge(97, 140) <= 4; angryBirdLarge(97, 141) <= 4; angryBirdLarge(97, 142) <= 4; angryBirdLarge(97, 143) <= 4; angryBirdLarge(97, 144) <= 5; angryBirdLarge(97, 145) <= 5; angryBirdLarge(97, 146) <= 5; angryBirdLarge(97, 147) <= 5; angryBirdLarge(97, 148) <= 5; angryBirdLarge(97, 149) <= 5; 
angryBirdLarge(98, 0) <= 0; angryBirdLarge(98, 1) <= 0; angryBirdLarge(98, 2) <= 0; angryBirdLarge(98, 3) <= 0; angryBirdLarge(98, 4) <= 0; angryBirdLarge(98, 5) <= 0; angryBirdLarge(98, 6) <= 5; angryBirdLarge(98, 7) <= 5; angryBirdLarge(98, 8) <= 5; angryBirdLarge(98, 9) <= 5; angryBirdLarge(98, 10) <= 5; angryBirdLarge(98, 11) <= 5; angryBirdLarge(98, 12) <= 5; angryBirdLarge(98, 13) <= 5; angryBirdLarge(98, 14) <= 5; angryBirdLarge(98, 15) <= 5; angryBirdLarge(98, 16) <= 5; angryBirdLarge(98, 17) <= 5; angryBirdLarge(98, 18) <= 0; angryBirdLarge(98, 19) <= 0; angryBirdLarge(98, 20) <= 0; angryBirdLarge(98, 21) <= 0; angryBirdLarge(98, 22) <= 0; angryBirdLarge(98, 23) <= 0; angryBirdLarge(98, 24) <= 4; angryBirdLarge(98, 25) <= 4; angryBirdLarge(98, 26) <= 4; angryBirdLarge(98, 27) <= 4; angryBirdLarge(98, 28) <= 4; angryBirdLarge(98, 29) <= 4; angryBirdLarge(98, 30) <= 4; angryBirdLarge(98, 31) <= 4; angryBirdLarge(98, 32) <= 4; angryBirdLarge(98, 33) <= 4; angryBirdLarge(98, 34) <= 4; angryBirdLarge(98, 35) <= 4; angryBirdLarge(98, 36) <= 4; angryBirdLarge(98, 37) <= 4; angryBirdLarge(98, 38) <= 4; angryBirdLarge(98, 39) <= 4; angryBirdLarge(98, 40) <= 4; angryBirdLarge(98, 41) <= 4; angryBirdLarge(98, 42) <= 4; angryBirdLarge(98, 43) <= 4; angryBirdLarge(98, 44) <= 4; angryBirdLarge(98, 45) <= 4; angryBirdLarge(98, 46) <= 4; angryBirdLarge(98, 47) <= 4; angryBirdLarge(98, 48) <= 4; angryBirdLarge(98, 49) <= 4; angryBirdLarge(98, 50) <= 4; angryBirdLarge(98, 51) <= 4; angryBirdLarge(98, 52) <= 4; angryBirdLarge(98, 53) <= 4; angryBirdLarge(98, 54) <= 4; angryBirdLarge(98, 55) <= 4; angryBirdLarge(98, 56) <= 4; angryBirdLarge(98, 57) <= 4; angryBirdLarge(98, 58) <= 4; angryBirdLarge(98, 59) <= 4; angryBirdLarge(98, 60) <= 4; angryBirdLarge(98, 61) <= 4; angryBirdLarge(98, 62) <= 4; angryBirdLarge(98, 63) <= 4; angryBirdLarge(98, 64) <= 4; angryBirdLarge(98, 65) <= 4; angryBirdLarge(98, 66) <= 4; angryBirdLarge(98, 67) <= 4; angryBirdLarge(98, 68) <= 4; angryBirdLarge(98, 69) <= 4; angryBirdLarge(98, 70) <= 4; angryBirdLarge(98, 71) <= 4; angryBirdLarge(98, 72) <= 4; angryBirdLarge(98, 73) <= 4; angryBirdLarge(98, 74) <= 4; angryBirdLarge(98, 75) <= 4; angryBirdLarge(98, 76) <= 4; angryBirdLarge(98, 77) <= 4; angryBirdLarge(98, 78) <= 4; angryBirdLarge(98, 79) <= 4; angryBirdLarge(98, 80) <= 4; angryBirdLarge(98, 81) <= 4; angryBirdLarge(98, 82) <= 4; angryBirdLarge(98, 83) <= 4; angryBirdLarge(98, 84) <= 4; angryBirdLarge(98, 85) <= 4; angryBirdLarge(98, 86) <= 4; angryBirdLarge(98, 87) <= 4; angryBirdLarge(98, 88) <= 4; angryBirdLarge(98, 89) <= 4; angryBirdLarge(98, 90) <= 5; angryBirdLarge(98, 91) <= 5; angryBirdLarge(98, 92) <= 5; angryBirdLarge(98, 93) <= 5; angryBirdLarge(98, 94) <= 5; angryBirdLarge(98, 95) <= 5; angryBirdLarge(98, 96) <= 3; angryBirdLarge(98, 97) <= 3; angryBirdLarge(98, 98) <= 3; angryBirdLarge(98, 99) <= 3; angryBirdLarge(98, 100) <= 3; angryBirdLarge(98, 101) <= 3; angryBirdLarge(98, 102) <= 3; angryBirdLarge(98, 103) <= 3; angryBirdLarge(98, 104) <= 3; angryBirdLarge(98, 105) <= 3; angryBirdLarge(98, 106) <= 3; angryBirdLarge(98, 107) <= 3; angryBirdLarge(98, 108) <= 3; angryBirdLarge(98, 109) <= 3; angryBirdLarge(98, 110) <= 3; angryBirdLarge(98, 111) <= 3; angryBirdLarge(98, 112) <= 3; angryBirdLarge(98, 113) <= 3; angryBirdLarge(98, 114) <= 3; angryBirdLarge(98, 115) <= 3; angryBirdLarge(98, 116) <= 3; angryBirdLarge(98, 117) <= 3; angryBirdLarge(98, 118) <= 3; angryBirdLarge(98, 119) <= 3; angryBirdLarge(98, 120) <= 3; angryBirdLarge(98, 121) <= 3; angryBirdLarge(98, 122) <= 3; angryBirdLarge(98, 123) <= 3; angryBirdLarge(98, 124) <= 3; angryBirdLarge(98, 125) <= 3; angryBirdLarge(98, 126) <= 3; angryBirdLarge(98, 127) <= 3; angryBirdLarge(98, 128) <= 3; angryBirdLarge(98, 129) <= 3; angryBirdLarge(98, 130) <= 3; angryBirdLarge(98, 131) <= 3; angryBirdLarge(98, 132) <= 5; angryBirdLarge(98, 133) <= 5; angryBirdLarge(98, 134) <= 5; angryBirdLarge(98, 135) <= 5; angryBirdLarge(98, 136) <= 5; angryBirdLarge(98, 137) <= 5; angryBirdLarge(98, 138) <= 4; angryBirdLarge(98, 139) <= 4; angryBirdLarge(98, 140) <= 4; angryBirdLarge(98, 141) <= 4; angryBirdLarge(98, 142) <= 4; angryBirdLarge(98, 143) <= 4; angryBirdLarge(98, 144) <= 5; angryBirdLarge(98, 145) <= 5; angryBirdLarge(98, 146) <= 5; angryBirdLarge(98, 147) <= 5; angryBirdLarge(98, 148) <= 5; angryBirdLarge(98, 149) <= 5; 
angryBirdLarge(99, 0) <= 0; angryBirdLarge(99, 1) <= 0; angryBirdLarge(99, 2) <= 0; angryBirdLarge(99, 3) <= 0; angryBirdLarge(99, 4) <= 0; angryBirdLarge(99, 5) <= 0; angryBirdLarge(99, 6) <= 5; angryBirdLarge(99, 7) <= 5; angryBirdLarge(99, 8) <= 5; angryBirdLarge(99, 9) <= 5; angryBirdLarge(99, 10) <= 5; angryBirdLarge(99, 11) <= 5; angryBirdLarge(99, 12) <= 5; angryBirdLarge(99, 13) <= 5; angryBirdLarge(99, 14) <= 5; angryBirdLarge(99, 15) <= 5; angryBirdLarge(99, 16) <= 5; angryBirdLarge(99, 17) <= 5; angryBirdLarge(99, 18) <= 0; angryBirdLarge(99, 19) <= 0; angryBirdLarge(99, 20) <= 0; angryBirdLarge(99, 21) <= 0; angryBirdLarge(99, 22) <= 0; angryBirdLarge(99, 23) <= 0; angryBirdLarge(99, 24) <= 4; angryBirdLarge(99, 25) <= 4; angryBirdLarge(99, 26) <= 4; angryBirdLarge(99, 27) <= 4; angryBirdLarge(99, 28) <= 4; angryBirdLarge(99, 29) <= 4; angryBirdLarge(99, 30) <= 4; angryBirdLarge(99, 31) <= 4; angryBirdLarge(99, 32) <= 4; angryBirdLarge(99, 33) <= 4; angryBirdLarge(99, 34) <= 4; angryBirdLarge(99, 35) <= 4; angryBirdLarge(99, 36) <= 4; angryBirdLarge(99, 37) <= 4; angryBirdLarge(99, 38) <= 4; angryBirdLarge(99, 39) <= 4; angryBirdLarge(99, 40) <= 4; angryBirdLarge(99, 41) <= 4; angryBirdLarge(99, 42) <= 4; angryBirdLarge(99, 43) <= 4; angryBirdLarge(99, 44) <= 4; angryBirdLarge(99, 45) <= 4; angryBirdLarge(99, 46) <= 4; angryBirdLarge(99, 47) <= 4; angryBirdLarge(99, 48) <= 4; angryBirdLarge(99, 49) <= 4; angryBirdLarge(99, 50) <= 4; angryBirdLarge(99, 51) <= 4; angryBirdLarge(99, 52) <= 4; angryBirdLarge(99, 53) <= 4; angryBirdLarge(99, 54) <= 4; angryBirdLarge(99, 55) <= 4; angryBirdLarge(99, 56) <= 4; angryBirdLarge(99, 57) <= 4; angryBirdLarge(99, 58) <= 4; angryBirdLarge(99, 59) <= 4; angryBirdLarge(99, 60) <= 4; angryBirdLarge(99, 61) <= 4; angryBirdLarge(99, 62) <= 4; angryBirdLarge(99, 63) <= 4; angryBirdLarge(99, 64) <= 4; angryBirdLarge(99, 65) <= 4; angryBirdLarge(99, 66) <= 4; angryBirdLarge(99, 67) <= 4; angryBirdLarge(99, 68) <= 4; angryBirdLarge(99, 69) <= 4; angryBirdLarge(99, 70) <= 4; angryBirdLarge(99, 71) <= 4; angryBirdLarge(99, 72) <= 4; angryBirdLarge(99, 73) <= 4; angryBirdLarge(99, 74) <= 4; angryBirdLarge(99, 75) <= 4; angryBirdLarge(99, 76) <= 4; angryBirdLarge(99, 77) <= 4; angryBirdLarge(99, 78) <= 4; angryBirdLarge(99, 79) <= 4; angryBirdLarge(99, 80) <= 4; angryBirdLarge(99, 81) <= 4; angryBirdLarge(99, 82) <= 4; angryBirdLarge(99, 83) <= 4; angryBirdLarge(99, 84) <= 4; angryBirdLarge(99, 85) <= 4; angryBirdLarge(99, 86) <= 4; angryBirdLarge(99, 87) <= 4; angryBirdLarge(99, 88) <= 4; angryBirdLarge(99, 89) <= 4; angryBirdLarge(99, 90) <= 5; angryBirdLarge(99, 91) <= 5; angryBirdLarge(99, 92) <= 5; angryBirdLarge(99, 93) <= 5; angryBirdLarge(99, 94) <= 5; angryBirdLarge(99, 95) <= 5; angryBirdLarge(99, 96) <= 3; angryBirdLarge(99, 97) <= 3; angryBirdLarge(99, 98) <= 3; angryBirdLarge(99, 99) <= 3; angryBirdLarge(99, 100) <= 3; angryBirdLarge(99, 101) <= 3; angryBirdLarge(99, 102) <= 3; angryBirdLarge(99, 103) <= 3; angryBirdLarge(99, 104) <= 3; angryBirdLarge(99, 105) <= 3; angryBirdLarge(99, 106) <= 3; angryBirdLarge(99, 107) <= 3; angryBirdLarge(99, 108) <= 3; angryBirdLarge(99, 109) <= 3; angryBirdLarge(99, 110) <= 3; angryBirdLarge(99, 111) <= 3; angryBirdLarge(99, 112) <= 3; angryBirdLarge(99, 113) <= 3; angryBirdLarge(99, 114) <= 3; angryBirdLarge(99, 115) <= 3; angryBirdLarge(99, 116) <= 3; angryBirdLarge(99, 117) <= 3; angryBirdLarge(99, 118) <= 3; angryBirdLarge(99, 119) <= 3; angryBirdLarge(99, 120) <= 3; angryBirdLarge(99, 121) <= 3; angryBirdLarge(99, 122) <= 3; angryBirdLarge(99, 123) <= 3; angryBirdLarge(99, 124) <= 3; angryBirdLarge(99, 125) <= 3; angryBirdLarge(99, 126) <= 3; angryBirdLarge(99, 127) <= 3; angryBirdLarge(99, 128) <= 3; angryBirdLarge(99, 129) <= 3; angryBirdLarge(99, 130) <= 3; angryBirdLarge(99, 131) <= 3; angryBirdLarge(99, 132) <= 5; angryBirdLarge(99, 133) <= 5; angryBirdLarge(99, 134) <= 5; angryBirdLarge(99, 135) <= 5; angryBirdLarge(99, 136) <= 5; angryBirdLarge(99, 137) <= 5; angryBirdLarge(99, 138) <= 4; angryBirdLarge(99, 139) <= 4; angryBirdLarge(99, 140) <= 4; angryBirdLarge(99, 141) <= 4; angryBirdLarge(99, 142) <= 4; angryBirdLarge(99, 143) <= 4; angryBirdLarge(99, 144) <= 5; angryBirdLarge(99, 145) <= 5; angryBirdLarge(99, 146) <= 5; angryBirdLarge(99, 147) <= 5; angryBirdLarge(99, 148) <= 5; angryBirdLarge(99, 149) <= 5; 
angryBirdLarge(100, 0) <= 0; angryBirdLarge(100, 1) <= 0; angryBirdLarge(100, 2) <= 0; angryBirdLarge(100, 3) <= 0; angryBirdLarge(100, 4) <= 0; angryBirdLarge(100, 5) <= 0; angryBirdLarge(100, 6) <= 5; angryBirdLarge(100, 7) <= 5; angryBirdLarge(100, 8) <= 5; angryBirdLarge(100, 9) <= 5; angryBirdLarge(100, 10) <= 5; angryBirdLarge(100, 11) <= 5; angryBirdLarge(100, 12) <= 5; angryBirdLarge(100, 13) <= 5; angryBirdLarge(100, 14) <= 5; angryBirdLarge(100, 15) <= 5; angryBirdLarge(100, 16) <= 5; angryBirdLarge(100, 17) <= 5; angryBirdLarge(100, 18) <= 0; angryBirdLarge(100, 19) <= 0; angryBirdLarge(100, 20) <= 0; angryBirdLarge(100, 21) <= 0; angryBirdLarge(100, 22) <= 0; angryBirdLarge(100, 23) <= 0; angryBirdLarge(100, 24) <= 4; angryBirdLarge(100, 25) <= 4; angryBirdLarge(100, 26) <= 4; angryBirdLarge(100, 27) <= 4; angryBirdLarge(100, 28) <= 4; angryBirdLarge(100, 29) <= 4; angryBirdLarge(100, 30) <= 4; angryBirdLarge(100, 31) <= 4; angryBirdLarge(100, 32) <= 4; angryBirdLarge(100, 33) <= 4; angryBirdLarge(100, 34) <= 4; angryBirdLarge(100, 35) <= 4; angryBirdLarge(100, 36) <= 4; angryBirdLarge(100, 37) <= 4; angryBirdLarge(100, 38) <= 4; angryBirdLarge(100, 39) <= 4; angryBirdLarge(100, 40) <= 4; angryBirdLarge(100, 41) <= 4; angryBirdLarge(100, 42) <= 4; angryBirdLarge(100, 43) <= 4; angryBirdLarge(100, 44) <= 4; angryBirdLarge(100, 45) <= 4; angryBirdLarge(100, 46) <= 4; angryBirdLarge(100, 47) <= 4; angryBirdLarge(100, 48) <= 4; angryBirdLarge(100, 49) <= 4; angryBirdLarge(100, 50) <= 4; angryBirdLarge(100, 51) <= 4; angryBirdLarge(100, 52) <= 4; angryBirdLarge(100, 53) <= 4; angryBirdLarge(100, 54) <= 4; angryBirdLarge(100, 55) <= 4; angryBirdLarge(100, 56) <= 4; angryBirdLarge(100, 57) <= 4; angryBirdLarge(100, 58) <= 4; angryBirdLarge(100, 59) <= 4; angryBirdLarge(100, 60) <= 4; angryBirdLarge(100, 61) <= 4; angryBirdLarge(100, 62) <= 4; angryBirdLarge(100, 63) <= 4; angryBirdLarge(100, 64) <= 4; angryBirdLarge(100, 65) <= 4; angryBirdLarge(100, 66) <= 4; angryBirdLarge(100, 67) <= 4; angryBirdLarge(100, 68) <= 4; angryBirdLarge(100, 69) <= 4; angryBirdLarge(100, 70) <= 4; angryBirdLarge(100, 71) <= 4; angryBirdLarge(100, 72) <= 4; angryBirdLarge(100, 73) <= 4; angryBirdLarge(100, 74) <= 4; angryBirdLarge(100, 75) <= 4; angryBirdLarge(100, 76) <= 4; angryBirdLarge(100, 77) <= 4; angryBirdLarge(100, 78) <= 4; angryBirdLarge(100, 79) <= 4; angryBirdLarge(100, 80) <= 4; angryBirdLarge(100, 81) <= 4; angryBirdLarge(100, 82) <= 4; angryBirdLarge(100, 83) <= 4; angryBirdLarge(100, 84) <= 4; angryBirdLarge(100, 85) <= 4; angryBirdLarge(100, 86) <= 4; angryBirdLarge(100, 87) <= 4; angryBirdLarge(100, 88) <= 4; angryBirdLarge(100, 89) <= 4; angryBirdLarge(100, 90) <= 5; angryBirdLarge(100, 91) <= 5; angryBirdLarge(100, 92) <= 5; angryBirdLarge(100, 93) <= 5; angryBirdLarge(100, 94) <= 5; angryBirdLarge(100, 95) <= 5; angryBirdLarge(100, 96) <= 3; angryBirdLarge(100, 97) <= 3; angryBirdLarge(100, 98) <= 3; angryBirdLarge(100, 99) <= 3; angryBirdLarge(100, 100) <= 3; angryBirdLarge(100, 101) <= 3; angryBirdLarge(100, 102) <= 3; angryBirdLarge(100, 103) <= 3; angryBirdLarge(100, 104) <= 3; angryBirdLarge(100, 105) <= 3; angryBirdLarge(100, 106) <= 3; angryBirdLarge(100, 107) <= 3; angryBirdLarge(100, 108) <= 3; angryBirdLarge(100, 109) <= 3; angryBirdLarge(100, 110) <= 3; angryBirdLarge(100, 111) <= 3; angryBirdLarge(100, 112) <= 3; angryBirdLarge(100, 113) <= 3; angryBirdLarge(100, 114) <= 3; angryBirdLarge(100, 115) <= 3; angryBirdLarge(100, 116) <= 3; angryBirdLarge(100, 117) <= 3; angryBirdLarge(100, 118) <= 3; angryBirdLarge(100, 119) <= 3; angryBirdLarge(100, 120) <= 3; angryBirdLarge(100, 121) <= 3; angryBirdLarge(100, 122) <= 3; angryBirdLarge(100, 123) <= 3; angryBirdLarge(100, 124) <= 3; angryBirdLarge(100, 125) <= 3; angryBirdLarge(100, 126) <= 3; angryBirdLarge(100, 127) <= 3; angryBirdLarge(100, 128) <= 3; angryBirdLarge(100, 129) <= 3; angryBirdLarge(100, 130) <= 3; angryBirdLarge(100, 131) <= 3; angryBirdLarge(100, 132) <= 5; angryBirdLarge(100, 133) <= 5; angryBirdLarge(100, 134) <= 5; angryBirdLarge(100, 135) <= 5; angryBirdLarge(100, 136) <= 5; angryBirdLarge(100, 137) <= 5; angryBirdLarge(100, 138) <= 4; angryBirdLarge(100, 139) <= 4; angryBirdLarge(100, 140) <= 4; angryBirdLarge(100, 141) <= 4; angryBirdLarge(100, 142) <= 4; angryBirdLarge(100, 143) <= 4; angryBirdLarge(100, 144) <= 5; angryBirdLarge(100, 145) <= 5; angryBirdLarge(100, 146) <= 5; angryBirdLarge(100, 147) <= 5; angryBirdLarge(100, 148) <= 5; angryBirdLarge(100, 149) <= 5; 
angryBirdLarge(101, 0) <= 0; angryBirdLarge(101, 1) <= 0; angryBirdLarge(101, 2) <= 0; angryBirdLarge(101, 3) <= 0; angryBirdLarge(101, 4) <= 0; angryBirdLarge(101, 5) <= 0; angryBirdLarge(101, 6) <= 5; angryBirdLarge(101, 7) <= 5; angryBirdLarge(101, 8) <= 5; angryBirdLarge(101, 9) <= 5; angryBirdLarge(101, 10) <= 5; angryBirdLarge(101, 11) <= 5; angryBirdLarge(101, 12) <= 5; angryBirdLarge(101, 13) <= 5; angryBirdLarge(101, 14) <= 5; angryBirdLarge(101, 15) <= 5; angryBirdLarge(101, 16) <= 5; angryBirdLarge(101, 17) <= 5; angryBirdLarge(101, 18) <= 0; angryBirdLarge(101, 19) <= 0; angryBirdLarge(101, 20) <= 0; angryBirdLarge(101, 21) <= 0; angryBirdLarge(101, 22) <= 0; angryBirdLarge(101, 23) <= 0; angryBirdLarge(101, 24) <= 4; angryBirdLarge(101, 25) <= 4; angryBirdLarge(101, 26) <= 4; angryBirdLarge(101, 27) <= 4; angryBirdLarge(101, 28) <= 4; angryBirdLarge(101, 29) <= 4; angryBirdLarge(101, 30) <= 4; angryBirdLarge(101, 31) <= 4; angryBirdLarge(101, 32) <= 4; angryBirdLarge(101, 33) <= 4; angryBirdLarge(101, 34) <= 4; angryBirdLarge(101, 35) <= 4; angryBirdLarge(101, 36) <= 4; angryBirdLarge(101, 37) <= 4; angryBirdLarge(101, 38) <= 4; angryBirdLarge(101, 39) <= 4; angryBirdLarge(101, 40) <= 4; angryBirdLarge(101, 41) <= 4; angryBirdLarge(101, 42) <= 4; angryBirdLarge(101, 43) <= 4; angryBirdLarge(101, 44) <= 4; angryBirdLarge(101, 45) <= 4; angryBirdLarge(101, 46) <= 4; angryBirdLarge(101, 47) <= 4; angryBirdLarge(101, 48) <= 4; angryBirdLarge(101, 49) <= 4; angryBirdLarge(101, 50) <= 4; angryBirdLarge(101, 51) <= 4; angryBirdLarge(101, 52) <= 4; angryBirdLarge(101, 53) <= 4; angryBirdLarge(101, 54) <= 4; angryBirdLarge(101, 55) <= 4; angryBirdLarge(101, 56) <= 4; angryBirdLarge(101, 57) <= 4; angryBirdLarge(101, 58) <= 4; angryBirdLarge(101, 59) <= 4; angryBirdLarge(101, 60) <= 4; angryBirdLarge(101, 61) <= 4; angryBirdLarge(101, 62) <= 4; angryBirdLarge(101, 63) <= 4; angryBirdLarge(101, 64) <= 4; angryBirdLarge(101, 65) <= 4; angryBirdLarge(101, 66) <= 4; angryBirdLarge(101, 67) <= 4; angryBirdLarge(101, 68) <= 4; angryBirdLarge(101, 69) <= 4; angryBirdLarge(101, 70) <= 4; angryBirdLarge(101, 71) <= 4; angryBirdLarge(101, 72) <= 4; angryBirdLarge(101, 73) <= 4; angryBirdLarge(101, 74) <= 4; angryBirdLarge(101, 75) <= 4; angryBirdLarge(101, 76) <= 4; angryBirdLarge(101, 77) <= 4; angryBirdLarge(101, 78) <= 4; angryBirdLarge(101, 79) <= 4; angryBirdLarge(101, 80) <= 4; angryBirdLarge(101, 81) <= 4; angryBirdLarge(101, 82) <= 4; angryBirdLarge(101, 83) <= 4; angryBirdLarge(101, 84) <= 4; angryBirdLarge(101, 85) <= 4; angryBirdLarge(101, 86) <= 4; angryBirdLarge(101, 87) <= 4; angryBirdLarge(101, 88) <= 4; angryBirdLarge(101, 89) <= 4; angryBirdLarge(101, 90) <= 5; angryBirdLarge(101, 91) <= 5; angryBirdLarge(101, 92) <= 5; angryBirdLarge(101, 93) <= 5; angryBirdLarge(101, 94) <= 5; angryBirdLarge(101, 95) <= 5; angryBirdLarge(101, 96) <= 3; angryBirdLarge(101, 97) <= 3; angryBirdLarge(101, 98) <= 3; angryBirdLarge(101, 99) <= 3; angryBirdLarge(101, 100) <= 3; angryBirdLarge(101, 101) <= 3; angryBirdLarge(101, 102) <= 3; angryBirdLarge(101, 103) <= 3; angryBirdLarge(101, 104) <= 3; angryBirdLarge(101, 105) <= 3; angryBirdLarge(101, 106) <= 3; angryBirdLarge(101, 107) <= 3; angryBirdLarge(101, 108) <= 3; angryBirdLarge(101, 109) <= 3; angryBirdLarge(101, 110) <= 3; angryBirdLarge(101, 111) <= 3; angryBirdLarge(101, 112) <= 3; angryBirdLarge(101, 113) <= 3; angryBirdLarge(101, 114) <= 3; angryBirdLarge(101, 115) <= 3; angryBirdLarge(101, 116) <= 3; angryBirdLarge(101, 117) <= 3; angryBirdLarge(101, 118) <= 3; angryBirdLarge(101, 119) <= 3; angryBirdLarge(101, 120) <= 3; angryBirdLarge(101, 121) <= 3; angryBirdLarge(101, 122) <= 3; angryBirdLarge(101, 123) <= 3; angryBirdLarge(101, 124) <= 3; angryBirdLarge(101, 125) <= 3; angryBirdLarge(101, 126) <= 3; angryBirdLarge(101, 127) <= 3; angryBirdLarge(101, 128) <= 3; angryBirdLarge(101, 129) <= 3; angryBirdLarge(101, 130) <= 3; angryBirdLarge(101, 131) <= 3; angryBirdLarge(101, 132) <= 5; angryBirdLarge(101, 133) <= 5; angryBirdLarge(101, 134) <= 5; angryBirdLarge(101, 135) <= 5; angryBirdLarge(101, 136) <= 5; angryBirdLarge(101, 137) <= 5; angryBirdLarge(101, 138) <= 4; angryBirdLarge(101, 139) <= 4; angryBirdLarge(101, 140) <= 4; angryBirdLarge(101, 141) <= 4; angryBirdLarge(101, 142) <= 4; angryBirdLarge(101, 143) <= 4; angryBirdLarge(101, 144) <= 5; angryBirdLarge(101, 145) <= 5; angryBirdLarge(101, 146) <= 5; angryBirdLarge(101, 147) <= 5; angryBirdLarge(101, 148) <= 5; angryBirdLarge(101, 149) <= 5; 
angryBirdLarge(102, 0) <= 0; angryBirdLarge(102, 1) <= 0; angryBirdLarge(102, 2) <= 0; angryBirdLarge(102, 3) <= 0; angryBirdLarge(102, 4) <= 0; angryBirdLarge(102, 5) <= 0; angryBirdLarge(102, 6) <= 0; angryBirdLarge(102, 7) <= 0; angryBirdLarge(102, 8) <= 0; angryBirdLarge(102, 9) <= 0; angryBirdLarge(102, 10) <= 0; angryBirdLarge(102, 11) <= 0; angryBirdLarge(102, 12) <= 0; angryBirdLarge(102, 13) <= 0; angryBirdLarge(102, 14) <= 0; angryBirdLarge(102, 15) <= 0; angryBirdLarge(102, 16) <= 0; angryBirdLarge(102, 17) <= 0; angryBirdLarge(102, 18) <= 0; angryBirdLarge(102, 19) <= 0; angryBirdLarge(102, 20) <= 0; angryBirdLarge(102, 21) <= 0; angryBirdLarge(102, 22) <= 0; angryBirdLarge(102, 23) <= 0; angryBirdLarge(102, 24) <= 5; angryBirdLarge(102, 25) <= 5; angryBirdLarge(102, 26) <= 5; angryBirdLarge(102, 27) <= 5; angryBirdLarge(102, 28) <= 5; angryBirdLarge(102, 29) <= 5; angryBirdLarge(102, 30) <= 4; angryBirdLarge(102, 31) <= 4; angryBirdLarge(102, 32) <= 4; angryBirdLarge(102, 33) <= 4; angryBirdLarge(102, 34) <= 4; angryBirdLarge(102, 35) <= 4; angryBirdLarge(102, 36) <= 4; angryBirdLarge(102, 37) <= 4; angryBirdLarge(102, 38) <= 4; angryBirdLarge(102, 39) <= 4; angryBirdLarge(102, 40) <= 4; angryBirdLarge(102, 41) <= 4; angryBirdLarge(102, 42) <= 4; angryBirdLarge(102, 43) <= 4; angryBirdLarge(102, 44) <= 4; angryBirdLarge(102, 45) <= 4; angryBirdLarge(102, 46) <= 4; angryBirdLarge(102, 47) <= 4; angryBirdLarge(102, 48) <= 4; angryBirdLarge(102, 49) <= 4; angryBirdLarge(102, 50) <= 4; angryBirdLarge(102, 51) <= 4; angryBirdLarge(102, 52) <= 4; angryBirdLarge(102, 53) <= 4; angryBirdLarge(102, 54) <= 4; angryBirdLarge(102, 55) <= 4; angryBirdLarge(102, 56) <= 4; angryBirdLarge(102, 57) <= 4; angryBirdLarge(102, 58) <= 4; angryBirdLarge(102, 59) <= 4; angryBirdLarge(102, 60) <= 4; angryBirdLarge(102, 61) <= 4; angryBirdLarge(102, 62) <= 4; angryBirdLarge(102, 63) <= 4; angryBirdLarge(102, 64) <= 4; angryBirdLarge(102, 65) <= 4; angryBirdLarge(102, 66) <= 2; angryBirdLarge(102, 67) <= 2; angryBirdLarge(102, 68) <= 2; angryBirdLarge(102, 69) <= 2; angryBirdLarge(102, 70) <= 2; angryBirdLarge(102, 71) <= 2; angryBirdLarge(102, 72) <= 2; angryBirdLarge(102, 73) <= 2; angryBirdLarge(102, 74) <= 2; angryBirdLarge(102, 75) <= 2; angryBirdLarge(102, 76) <= 2; angryBirdLarge(102, 77) <= 2; angryBirdLarge(102, 78) <= 2; angryBirdLarge(102, 79) <= 2; angryBirdLarge(102, 80) <= 2; angryBirdLarge(102, 81) <= 2; angryBirdLarge(102, 82) <= 2; angryBirdLarge(102, 83) <= 2; angryBirdLarge(102, 84) <= 2; angryBirdLarge(102, 85) <= 2; angryBirdLarge(102, 86) <= 2; angryBirdLarge(102, 87) <= 2; angryBirdLarge(102, 88) <= 2; angryBirdLarge(102, 89) <= 2; angryBirdLarge(102, 90) <= 5; angryBirdLarge(102, 91) <= 5; angryBirdLarge(102, 92) <= 5; angryBirdLarge(102, 93) <= 5; angryBirdLarge(102, 94) <= 5; angryBirdLarge(102, 95) <= 5; angryBirdLarge(102, 96) <= 3; angryBirdLarge(102, 97) <= 3; angryBirdLarge(102, 98) <= 3; angryBirdLarge(102, 99) <= 3; angryBirdLarge(102, 100) <= 3; angryBirdLarge(102, 101) <= 3; angryBirdLarge(102, 102) <= 5; angryBirdLarge(102, 103) <= 5; angryBirdLarge(102, 104) <= 5; angryBirdLarge(102, 105) <= 5; angryBirdLarge(102, 106) <= 5; angryBirdLarge(102, 107) <= 5; angryBirdLarge(102, 108) <= 5; angryBirdLarge(102, 109) <= 5; angryBirdLarge(102, 110) <= 5; angryBirdLarge(102, 111) <= 5; angryBirdLarge(102, 112) <= 5; angryBirdLarge(102, 113) <= 5; angryBirdLarge(102, 114) <= 3; angryBirdLarge(102, 115) <= 3; angryBirdLarge(102, 116) <= 3; angryBirdLarge(102, 117) <= 3; angryBirdLarge(102, 118) <= 3; angryBirdLarge(102, 119) <= 3; angryBirdLarge(102, 120) <= 3; angryBirdLarge(102, 121) <= 3; angryBirdLarge(102, 122) <= 3; angryBirdLarge(102, 123) <= 3; angryBirdLarge(102, 124) <= 3; angryBirdLarge(102, 125) <= 3; angryBirdLarge(102, 126) <= 3; angryBirdLarge(102, 127) <= 3; angryBirdLarge(102, 128) <= 3; angryBirdLarge(102, 129) <= 3; angryBirdLarge(102, 130) <= 3; angryBirdLarge(102, 131) <= 3; angryBirdLarge(102, 132) <= 3; angryBirdLarge(102, 133) <= 3; angryBirdLarge(102, 134) <= 3; angryBirdLarge(102, 135) <= 3; angryBirdLarge(102, 136) <= 3; angryBirdLarge(102, 137) <= 3; angryBirdLarge(102, 138) <= 5; angryBirdLarge(102, 139) <= 5; angryBirdLarge(102, 140) <= 5; angryBirdLarge(102, 141) <= 5; angryBirdLarge(102, 142) <= 5; angryBirdLarge(102, 143) <= 5; angryBirdLarge(102, 144) <= 5; angryBirdLarge(102, 145) <= 5; angryBirdLarge(102, 146) <= 5; angryBirdLarge(102, 147) <= 5; angryBirdLarge(102, 148) <= 5; angryBirdLarge(102, 149) <= 5; 
angryBirdLarge(103, 0) <= 0; angryBirdLarge(103, 1) <= 0; angryBirdLarge(103, 2) <= 0; angryBirdLarge(103, 3) <= 0; angryBirdLarge(103, 4) <= 0; angryBirdLarge(103, 5) <= 0; angryBirdLarge(103, 6) <= 0; angryBirdLarge(103, 7) <= 0; angryBirdLarge(103, 8) <= 0; angryBirdLarge(103, 9) <= 0; angryBirdLarge(103, 10) <= 0; angryBirdLarge(103, 11) <= 0; angryBirdLarge(103, 12) <= 0; angryBirdLarge(103, 13) <= 0; angryBirdLarge(103, 14) <= 0; angryBirdLarge(103, 15) <= 0; angryBirdLarge(103, 16) <= 0; angryBirdLarge(103, 17) <= 0; angryBirdLarge(103, 18) <= 0; angryBirdLarge(103, 19) <= 0; angryBirdLarge(103, 20) <= 0; angryBirdLarge(103, 21) <= 0; angryBirdLarge(103, 22) <= 0; angryBirdLarge(103, 23) <= 0; angryBirdLarge(103, 24) <= 5; angryBirdLarge(103, 25) <= 5; angryBirdLarge(103, 26) <= 5; angryBirdLarge(103, 27) <= 5; angryBirdLarge(103, 28) <= 5; angryBirdLarge(103, 29) <= 5; angryBirdLarge(103, 30) <= 4; angryBirdLarge(103, 31) <= 4; angryBirdLarge(103, 32) <= 4; angryBirdLarge(103, 33) <= 4; angryBirdLarge(103, 34) <= 4; angryBirdLarge(103, 35) <= 4; angryBirdLarge(103, 36) <= 4; angryBirdLarge(103, 37) <= 4; angryBirdLarge(103, 38) <= 4; angryBirdLarge(103, 39) <= 4; angryBirdLarge(103, 40) <= 4; angryBirdLarge(103, 41) <= 4; angryBirdLarge(103, 42) <= 4; angryBirdLarge(103, 43) <= 4; angryBirdLarge(103, 44) <= 4; angryBirdLarge(103, 45) <= 4; angryBirdLarge(103, 46) <= 4; angryBirdLarge(103, 47) <= 4; angryBirdLarge(103, 48) <= 4; angryBirdLarge(103, 49) <= 4; angryBirdLarge(103, 50) <= 4; angryBirdLarge(103, 51) <= 4; angryBirdLarge(103, 52) <= 4; angryBirdLarge(103, 53) <= 4; angryBirdLarge(103, 54) <= 4; angryBirdLarge(103, 55) <= 4; angryBirdLarge(103, 56) <= 4; angryBirdLarge(103, 57) <= 4; angryBirdLarge(103, 58) <= 4; angryBirdLarge(103, 59) <= 4; angryBirdLarge(103, 60) <= 4; angryBirdLarge(103, 61) <= 4; angryBirdLarge(103, 62) <= 4; angryBirdLarge(103, 63) <= 4; angryBirdLarge(103, 64) <= 4; angryBirdLarge(103, 65) <= 4; angryBirdLarge(103, 66) <= 2; angryBirdLarge(103, 67) <= 2; angryBirdLarge(103, 68) <= 2; angryBirdLarge(103, 69) <= 2; angryBirdLarge(103, 70) <= 2; angryBirdLarge(103, 71) <= 2; angryBirdLarge(103, 72) <= 2; angryBirdLarge(103, 73) <= 2; angryBirdLarge(103, 74) <= 2; angryBirdLarge(103, 75) <= 2; angryBirdLarge(103, 76) <= 2; angryBirdLarge(103, 77) <= 2; angryBirdLarge(103, 78) <= 2; angryBirdLarge(103, 79) <= 2; angryBirdLarge(103, 80) <= 2; angryBirdLarge(103, 81) <= 2; angryBirdLarge(103, 82) <= 2; angryBirdLarge(103, 83) <= 2; angryBirdLarge(103, 84) <= 2; angryBirdLarge(103, 85) <= 2; angryBirdLarge(103, 86) <= 2; angryBirdLarge(103, 87) <= 2; angryBirdLarge(103, 88) <= 2; angryBirdLarge(103, 89) <= 2; angryBirdLarge(103, 90) <= 5; angryBirdLarge(103, 91) <= 5; angryBirdLarge(103, 92) <= 5; angryBirdLarge(103, 93) <= 5; angryBirdLarge(103, 94) <= 5; angryBirdLarge(103, 95) <= 5; angryBirdLarge(103, 96) <= 3; angryBirdLarge(103, 97) <= 3; angryBirdLarge(103, 98) <= 3; angryBirdLarge(103, 99) <= 3; angryBirdLarge(103, 100) <= 3; angryBirdLarge(103, 101) <= 3; angryBirdLarge(103, 102) <= 5; angryBirdLarge(103, 103) <= 5; angryBirdLarge(103, 104) <= 5; angryBirdLarge(103, 105) <= 5; angryBirdLarge(103, 106) <= 5; angryBirdLarge(103, 107) <= 5; angryBirdLarge(103, 108) <= 5; angryBirdLarge(103, 109) <= 5; angryBirdLarge(103, 110) <= 5; angryBirdLarge(103, 111) <= 5; angryBirdLarge(103, 112) <= 5; angryBirdLarge(103, 113) <= 5; angryBirdLarge(103, 114) <= 3; angryBirdLarge(103, 115) <= 3; angryBirdLarge(103, 116) <= 3; angryBirdLarge(103, 117) <= 3; angryBirdLarge(103, 118) <= 3; angryBirdLarge(103, 119) <= 3; angryBirdLarge(103, 120) <= 3; angryBirdLarge(103, 121) <= 3; angryBirdLarge(103, 122) <= 3; angryBirdLarge(103, 123) <= 3; angryBirdLarge(103, 124) <= 3; angryBirdLarge(103, 125) <= 3; angryBirdLarge(103, 126) <= 3; angryBirdLarge(103, 127) <= 3; angryBirdLarge(103, 128) <= 3; angryBirdLarge(103, 129) <= 3; angryBirdLarge(103, 130) <= 3; angryBirdLarge(103, 131) <= 3; angryBirdLarge(103, 132) <= 3; angryBirdLarge(103, 133) <= 3; angryBirdLarge(103, 134) <= 3; angryBirdLarge(103, 135) <= 3; angryBirdLarge(103, 136) <= 3; angryBirdLarge(103, 137) <= 3; angryBirdLarge(103, 138) <= 5; angryBirdLarge(103, 139) <= 5; angryBirdLarge(103, 140) <= 5; angryBirdLarge(103, 141) <= 5; angryBirdLarge(103, 142) <= 5; angryBirdLarge(103, 143) <= 5; angryBirdLarge(103, 144) <= 5; angryBirdLarge(103, 145) <= 5; angryBirdLarge(103, 146) <= 5; angryBirdLarge(103, 147) <= 5; angryBirdLarge(103, 148) <= 5; angryBirdLarge(103, 149) <= 5; 
angryBirdLarge(104, 0) <= 0; angryBirdLarge(104, 1) <= 0; angryBirdLarge(104, 2) <= 0; angryBirdLarge(104, 3) <= 0; angryBirdLarge(104, 4) <= 0; angryBirdLarge(104, 5) <= 0; angryBirdLarge(104, 6) <= 0; angryBirdLarge(104, 7) <= 0; angryBirdLarge(104, 8) <= 0; angryBirdLarge(104, 9) <= 0; angryBirdLarge(104, 10) <= 0; angryBirdLarge(104, 11) <= 0; angryBirdLarge(104, 12) <= 0; angryBirdLarge(104, 13) <= 0; angryBirdLarge(104, 14) <= 0; angryBirdLarge(104, 15) <= 0; angryBirdLarge(104, 16) <= 0; angryBirdLarge(104, 17) <= 0; angryBirdLarge(104, 18) <= 0; angryBirdLarge(104, 19) <= 0; angryBirdLarge(104, 20) <= 0; angryBirdLarge(104, 21) <= 0; angryBirdLarge(104, 22) <= 0; angryBirdLarge(104, 23) <= 0; angryBirdLarge(104, 24) <= 5; angryBirdLarge(104, 25) <= 5; angryBirdLarge(104, 26) <= 5; angryBirdLarge(104, 27) <= 5; angryBirdLarge(104, 28) <= 5; angryBirdLarge(104, 29) <= 5; angryBirdLarge(104, 30) <= 4; angryBirdLarge(104, 31) <= 4; angryBirdLarge(104, 32) <= 4; angryBirdLarge(104, 33) <= 4; angryBirdLarge(104, 34) <= 4; angryBirdLarge(104, 35) <= 4; angryBirdLarge(104, 36) <= 4; angryBirdLarge(104, 37) <= 4; angryBirdLarge(104, 38) <= 4; angryBirdLarge(104, 39) <= 4; angryBirdLarge(104, 40) <= 4; angryBirdLarge(104, 41) <= 4; angryBirdLarge(104, 42) <= 4; angryBirdLarge(104, 43) <= 4; angryBirdLarge(104, 44) <= 4; angryBirdLarge(104, 45) <= 4; angryBirdLarge(104, 46) <= 4; angryBirdLarge(104, 47) <= 4; angryBirdLarge(104, 48) <= 4; angryBirdLarge(104, 49) <= 4; angryBirdLarge(104, 50) <= 4; angryBirdLarge(104, 51) <= 4; angryBirdLarge(104, 52) <= 4; angryBirdLarge(104, 53) <= 4; angryBirdLarge(104, 54) <= 4; angryBirdLarge(104, 55) <= 4; angryBirdLarge(104, 56) <= 4; angryBirdLarge(104, 57) <= 4; angryBirdLarge(104, 58) <= 4; angryBirdLarge(104, 59) <= 4; angryBirdLarge(104, 60) <= 4; angryBirdLarge(104, 61) <= 4; angryBirdLarge(104, 62) <= 4; angryBirdLarge(104, 63) <= 4; angryBirdLarge(104, 64) <= 4; angryBirdLarge(104, 65) <= 4; angryBirdLarge(104, 66) <= 2; angryBirdLarge(104, 67) <= 2; angryBirdLarge(104, 68) <= 2; angryBirdLarge(104, 69) <= 2; angryBirdLarge(104, 70) <= 2; angryBirdLarge(104, 71) <= 2; angryBirdLarge(104, 72) <= 2; angryBirdLarge(104, 73) <= 2; angryBirdLarge(104, 74) <= 2; angryBirdLarge(104, 75) <= 2; angryBirdLarge(104, 76) <= 2; angryBirdLarge(104, 77) <= 2; angryBirdLarge(104, 78) <= 2; angryBirdLarge(104, 79) <= 2; angryBirdLarge(104, 80) <= 2; angryBirdLarge(104, 81) <= 2; angryBirdLarge(104, 82) <= 2; angryBirdLarge(104, 83) <= 2; angryBirdLarge(104, 84) <= 2; angryBirdLarge(104, 85) <= 2; angryBirdLarge(104, 86) <= 2; angryBirdLarge(104, 87) <= 2; angryBirdLarge(104, 88) <= 2; angryBirdLarge(104, 89) <= 2; angryBirdLarge(104, 90) <= 5; angryBirdLarge(104, 91) <= 5; angryBirdLarge(104, 92) <= 5; angryBirdLarge(104, 93) <= 5; angryBirdLarge(104, 94) <= 5; angryBirdLarge(104, 95) <= 5; angryBirdLarge(104, 96) <= 3; angryBirdLarge(104, 97) <= 3; angryBirdLarge(104, 98) <= 3; angryBirdLarge(104, 99) <= 3; angryBirdLarge(104, 100) <= 3; angryBirdLarge(104, 101) <= 3; angryBirdLarge(104, 102) <= 5; angryBirdLarge(104, 103) <= 5; angryBirdLarge(104, 104) <= 5; angryBirdLarge(104, 105) <= 5; angryBirdLarge(104, 106) <= 5; angryBirdLarge(104, 107) <= 5; angryBirdLarge(104, 108) <= 5; angryBirdLarge(104, 109) <= 5; angryBirdLarge(104, 110) <= 5; angryBirdLarge(104, 111) <= 5; angryBirdLarge(104, 112) <= 5; angryBirdLarge(104, 113) <= 5; angryBirdLarge(104, 114) <= 3; angryBirdLarge(104, 115) <= 3; angryBirdLarge(104, 116) <= 3; angryBirdLarge(104, 117) <= 3; angryBirdLarge(104, 118) <= 3; angryBirdLarge(104, 119) <= 3; angryBirdLarge(104, 120) <= 3; angryBirdLarge(104, 121) <= 3; angryBirdLarge(104, 122) <= 3; angryBirdLarge(104, 123) <= 3; angryBirdLarge(104, 124) <= 3; angryBirdLarge(104, 125) <= 3; angryBirdLarge(104, 126) <= 3; angryBirdLarge(104, 127) <= 3; angryBirdLarge(104, 128) <= 3; angryBirdLarge(104, 129) <= 3; angryBirdLarge(104, 130) <= 3; angryBirdLarge(104, 131) <= 3; angryBirdLarge(104, 132) <= 3; angryBirdLarge(104, 133) <= 3; angryBirdLarge(104, 134) <= 3; angryBirdLarge(104, 135) <= 3; angryBirdLarge(104, 136) <= 3; angryBirdLarge(104, 137) <= 3; angryBirdLarge(104, 138) <= 5; angryBirdLarge(104, 139) <= 5; angryBirdLarge(104, 140) <= 5; angryBirdLarge(104, 141) <= 5; angryBirdLarge(104, 142) <= 5; angryBirdLarge(104, 143) <= 5; angryBirdLarge(104, 144) <= 5; angryBirdLarge(104, 145) <= 5; angryBirdLarge(104, 146) <= 5; angryBirdLarge(104, 147) <= 5; angryBirdLarge(104, 148) <= 5; angryBirdLarge(104, 149) <= 5; 
angryBirdLarge(105, 0) <= 0; angryBirdLarge(105, 1) <= 0; angryBirdLarge(105, 2) <= 0; angryBirdLarge(105, 3) <= 0; angryBirdLarge(105, 4) <= 0; angryBirdLarge(105, 5) <= 0; angryBirdLarge(105, 6) <= 0; angryBirdLarge(105, 7) <= 0; angryBirdLarge(105, 8) <= 0; angryBirdLarge(105, 9) <= 0; angryBirdLarge(105, 10) <= 0; angryBirdLarge(105, 11) <= 0; angryBirdLarge(105, 12) <= 0; angryBirdLarge(105, 13) <= 0; angryBirdLarge(105, 14) <= 0; angryBirdLarge(105, 15) <= 0; angryBirdLarge(105, 16) <= 0; angryBirdLarge(105, 17) <= 0; angryBirdLarge(105, 18) <= 0; angryBirdLarge(105, 19) <= 0; angryBirdLarge(105, 20) <= 0; angryBirdLarge(105, 21) <= 0; angryBirdLarge(105, 22) <= 0; angryBirdLarge(105, 23) <= 0; angryBirdLarge(105, 24) <= 5; angryBirdLarge(105, 25) <= 5; angryBirdLarge(105, 26) <= 5; angryBirdLarge(105, 27) <= 5; angryBirdLarge(105, 28) <= 5; angryBirdLarge(105, 29) <= 5; angryBirdLarge(105, 30) <= 4; angryBirdLarge(105, 31) <= 4; angryBirdLarge(105, 32) <= 4; angryBirdLarge(105, 33) <= 4; angryBirdLarge(105, 34) <= 4; angryBirdLarge(105, 35) <= 4; angryBirdLarge(105, 36) <= 4; angryBirdLarge(105, 37) <= 4; angryBirdLarge(105, 38) <= 4; angryBirdLarge(105, 39) <= 4; angryBirdLarge(105, 40) <= 4; angryBirdLarge(105, 41) <= 4; angryBirdLarge(105, 42) <= 4; angryBirdLarge(105, 43) <= 4; angryBirdLarge(105, 44) <= 4; angryBirdLarge(105, 45) <= 4; angryBirdLarge(105, 46) <= 4; angryBirdLarge(105, 47) <= 4; angryBirdLarge(105, 48) <= 4; angryBirdLarge(105, 49) <= 4; angryBirdLarge(105, 50) <= 4; angryBirdLarge(105, 51) <= 4; angryBirdLarge(105, 52) <= 4; angryBirdLarge(105, 53) <= 4; angryBirdLarge(105, 54) <= 4; angryBirdLarge(105, 55) <= 4; angryBirdLarge(105, 56) <= 4; angryBirdLarge(105, 57) <= 4; angryBirdLarge(105, 58) <= 4; angryBirdLarge(105, 59) <= 4; angryBirdLarge(105, 60) <= 4; angryBirdLarge(105, 61) <= 4; angryBirdLarge(105, 62) <= 4; angryBirdLarge(105, 63) <= 4; angryBirdLarge(105, 64) <= 4; angryBirdLarge(105, 65) <= 4; angryBirdLarge(105, 66) <= 2; angryBirdLarge(105, 67) <= 2; angryBirdLarge(105, 68) <= 2; angryBirdLarge(105, 69) <= 2; angryBirdLarge(105, 70) <= 2; angryBirdLarge(105, 71) <= 2; angryBirdLarge(105, 72) <= 2; angryBirdLarge(105, 73) <= 2; angryBirdLarge(105, 74) <= 2; angryBirdLarge(105, 75) <= 2; angryBirdLarge(105, 76) <= 2; angryBirdLarge(105, 77) <= 2; angryBirdLarge(105, 78) <= 2; angryBirdLarge(105, 79) <= 2; angryBirdLarge(105, 80) <= 2; angryBirdLarge(105, 81) <= 2; angryBirdLarge(105, 82) <= 2; angryBirdLarge(105, 83) <= 2; angryBirdLarge(105, 84) <= 2; angryBirdLarge(105, 85) <= 2; angryBirdLarge(105, 86) <= 2; angryBirdLarge(105, 87) <= 2; angryBirdLarge(105, 88) <= 2; angryBirdLarge(105, 89) <= 2; angryBirdLarge(105, 90) <= 5; angryBirdLarge(105, 91) <= 5; angryBirdLarge(105, 92) <= 5; angryBirdLarge(105, 93) <= 5; angryBirdLarge(105, 94) <= 5; angryBirdLarge(105, 95) <= 5; angryBirdLarge(105, 96) <= 3; angryBirdLarge(105, 97) <= 3; angryBirdLarge(105, 98) <= 3; angryBirdLarge(105, 99) <= 3; angryBirdLarge(105, 100) <= 3; angryBirdLarge(105, 101) <= 3; angryBirdLarge(105, 102) <= 5; angryBirdLarge(105, 103) <= 5; angryBirdLarge(105, 104) <= 5; angryBirdLarge(105, 105) <= 5; angryBirdLarge(105, 106) <= 5; angryBirdLarge(105, 107) <= 5; angryBirdLarge(105, 108) <= 5; angryBirdLarge(105, 109) <= 5; angryBirdLarge(105, 110) <= 5; angryBirdLarge(105, 111) <= 5; angryBirdLarge(105, 112) <= 5; angryBirdLarge(105, 113) <= 5; angryBirdLarge(105, 114) <= 3; angryBirdLarge(105, 115) <= 3; angryBirdLarge(105, 116) <= 3; angryBirdLarge(105, 117) <= 3; angryBirdLarge(105, 118) <= 3; angryBirdLarge(105, 119) <= 3; angryBirdLarge(105, 120) <= 3; angryBirdLarge(105, 121) <= 3; angryBirdLarge(105, 122) <= 3; angryBirdLarge(105, 123) <= 3; angryBirdLarge(105, 124) <= 3; angryBirdLarge(105, 125) <= 3; angryBirdLarge(105, 126) <= 3; angryBirdLarge(105, 127) <= 3; angryBirdLarge(105, 128) <= 3; angryBirdLarge(105, 129) <= 3; angryBirdLarge(105, 130) <= 3; angryBirdLarge(105, 131) <= 3; angryBirdLarge(105, 132) <= 3; angryBirdLarge(105, 133) <= 3; angryBirdLarge(105, 134) <= 3; angryBirdLarge(105, 135) <= 3; angryBirdLarge(105, 136) <= 3; angryBirdLarge(105, 137) <= 3; angryBirdLarge(105, 138) <= 5; angryBirdLarge(105, 139) <= 5; angryBirdLarge(105, 140) <= 5; angryBirdLarge(105, 141) <= 5; angryBirdLarge(105, 142) <= 5; angryBirdLarge(105, 143) <= 5; angryBirdLarge(105, 144) <= 5; angryBirdLarge(105, 145) <= 5; angryBirdLarge(105, 146) <= 5; angryBirdLarge(105, 147) <= 5; angryBirdLarge(105, 148) <= 5; angryBirdLarge(105, 149) <= 5; 
angryBirdLarge(106, 0) <= 0; angryBirdLarge(106, 1) <= 0; angryBirdLarge(106, 2) <= 0; angryBirdLarge(106, 3) <= 0; angryBirdLarge(106, 4) <= 0; angryBirdLarge(106, 5) <= 0; angryBirdLarge(106, 6) <= 0; angryBirdLarge(106, 7) <= 0; angryBirdLarge(106, 8) <= 0; angryBirdLarge(106, 9) <= 0; angryBirdLarge(106, 10) <= 0; angryBirdLarge(106, 11) <= 0; angryBirdLarge(106, 12) <= 0; angryBirdLarge(106, 13) <= 0; angryBirdLarge(106, 14) <= 0; angryBirdLarge(106, 15) <= 0; angryBirdLarge(106, 16) <= 0; angryBirdLarge(106, 17) <= 0; angryBirdLarge(106, 18) <= 0; angryBirdLarge(106, 19) <= 0; angryBirdLarge(106, 20) <= 0; angryBirdLarge(106, 21) <= 0; angryBirdLarge(106, 22) <= 0; angryBirdLarge(106, 23) <= 0; angryBirdLarge(106, 24) <= 5; angryBirdLarge(106, 25) <= 5; angryBirdLarge(106, 26) <= 5; angryBirdLarge(106, 27) <= 5; angryBirdLarge(106, 28) <= 5; angryBirdLarge(106, 29) <= 5; angryBirdLarge(106, 30) <= 4; angryBirdLarge(106, 31) <= 4; angryBirdLarge(106, 32) <= 4; angryBirdLarge(106, 33) <= 4; angryBirdLarge(106, 34) <= 4; angryBirdLarge(106, 35) <= 4; angryBirdLarge(106, 36) <= 4; angryBirdLarge(106, 37) <= 4; angryBirdLarge(106, 38) <= 4; angryBirdLarge(106, 39) <= 4; angryBirdLarge(106, 40) <= 4; angryBirdLarge(106, 41) <= 4; angryBirdLarge(106, 42) <= 4; angryBirdLarge(106, 43) <= 4; angryBirdLarge(106, 44) <= 4; angryBirdLarge(106, 45) <= 4; angryBirdLarge(106, 46) <= 4; angryBirdLarge(106, 47) <= 4; angryBirdLarge(106, 48) <= 4; angryBirdLarge(106, 49) <= 4; angryBirdLarge(106, 50) <= 4; angryBirdLarge(106, 51) <= 4; angryBirdLarge(106, 52) <= 4; angryBirdLarge(106, 53) <= 4; angryBirdLarge(106, 54) <= 4; angryBirdLarge(106, 55) <= 4; angryBirdLarge(106, 56) <= 4; angryBirdLarge(106, 57) <= 4; angryBirdLarge(106, 58) <= 4; angryBirdLarge(106, 59) <= 4; angryBirdLarge(106, 60) <= 4; angryBirdLarge(106, 61) <= 4; angryBirdLarge(106, 62) <= 4; angryBirdLarge(106, 63) <= 4; angryBirdLarge(106, 64) <= 4; angryBirdLarge(106, 65) <= 4; angryBirdLarge(106, 66) <= 2; angryBirdLarge(106, 67) <= 2; angryBirdLarge(106, 68) <= 2; angryBirdLarge(106, 69) <= 2; angryBirdLarge(106, 70) <= 2; angryBirdLarge(106, 71) <= 2; angryBirdLarge(106, 72) <= 2; angryBirdLarge(106, 73) <= 2; angryBirdLarge(106, 74) <= 2; angryBirdLarge(106, 75) <= 2; angryBirdLarge(106, 76) <= 2; angryBirdLarge(106, 77) <= 2; angryBirdLarge(106, 78) <= 2; angryBirdLarge(106, 79) <= 2; angryBirdLarge(106, 80) <= 2; angryBirdLarge(106, 81) <= 2; angryBirdLarge(106, 82) <= 2; angryBirdLarge(106, 83) <= 2; angryBirdLarge(106, 84) <= 2; angryBirdLarge(106, 85) <= 2; angryBirdLarge(106, 86) <= 2; angryBirdLarge(106, 87) <= 2; angryBirdLarge(106, 88) <= 2; angryBirdLarge(106, 89) <= 2; angryBirdLarge(106, 90) <= 5; angryBirdLarge(106, 91) <= 5; angryBirdLarge(106, 92) <= 5; angryBirdLarge(106, 93) <= 5; angryBirdLarge(106, 94) <= 5; angryBirdLarge(106, 95) <= 5; angryBirdLarge(106, 96) <= 3; angryBirdLarge(106, 97) <= 3; angryBirdLarge(106, 98) <= 3; angryBirdLarge(106, 99) <= 3; angryBirdLarge(106, 100) <= 3; angryBirdLarge(106, 101) <= 3; angryBirdLarge(106, 102) <= 5; angryBirdLarge(106, 103) <= 5; angryBirdLarge(106, 104) <= 5; angryBirdLarge(106, 105) <= 5; angryBirdLarge(106, 106) <= 5; angryBirdLarge(106, 107) <= 5; angryBirdLarge(106, 108) <= 5; angryBirdLarge(106, 109) <= 5; angryBirdLarge(106, 110) <= 5; angryBirdLarge(106, 111) <= 5; angryBirdLarge(106, 112) <= 5; angryBirdLarge(106, 113) <= 5; angryBirdLarge(106, 114) <= 3; angryBirdLarge(106, 115) <= 3; angryBirdLarge(106, 116) <= 3; angryBirdLarge(106, 117) <= 3; angryBirdLarge(106, 118) <= 3; angryBirdLarge(106, 119) <= 3; angryBirdLarge(106, 120) <= 3; angryBirdLarge(106, 121) <= 3; angryBirdLarge(106, 122) <= 3; angryBirdLarge(106, 123) <= 3; angryBirdLarge(106, 124) <= 3; angryBirdLarge(106, 125) <= 3; angryBirdLarge(106, 126) <= 3; angryBirdLarge(106, 127) <= 3; angryBirdLarge(106, 128) <= 3; angryBirdLarge(106, 129) <= 3; angryBirdLarge(106, 130) <= 3; angryBirdLarge(106, 131) <= 3; angryBirdLarge(106, 132) <= 3; angryBirdLarge(106, 133) <= 3; angryBirdLarge(106, 134) <= 3; angryBirdLarge(106, 135) <= 3; angryBirdLarge(106, 136) <= 3; angryBirdLarge(106, 137) <= 3; angryBirdLarge(106, 138) <= 5; angryBirdLarge(106, 139) <= 5; angryBirdLarge(106, 140) <= 5; angryBirdLarge(106, 141) <= 5; angryBirdLarge(106, 142) <= 5; angryBirdLarge(106, 143) <= 5; angryBirdLarge(106, 144) <= 5; angryBirdLarge(106, 145) <= 5; angryBirdLarge(106, 146) <= 5; angryBirdLarge(106, 147) <= 5; angryBirdLarge(106, 148) <= 5; angryBirdLarge(106, 149) <= 5; 
angryBirdLarge(107, 0) <= 0; angryBirdLarge(107, 1) <= 0; angryBirdLarge(107, 2) <= 0; angryBirdLarge(107, 3) <= 0; angryBirdLarge(107, 4) <= 0; angryBirdLarge(107, 5) <= 0; angryBirdLarge(107, 6) <= 0; angryBirdLarge(107, 7) <= 0; angryBirdLarge(107, 8) <= 0; angryBirdLarge(107, 9) <= 0; angryBirdLarge(107, 10) <= 0; angryBirdLarge(107, 11) <= 0; angryBirdLarge(107, 12) <= 0; angryBirdLarge(107, 13) <= 0; angryBirdLarge(107, 14) <= 0; angryBirdLarge(107, 15) <= 0; angryBirdLarge(107, 16) <= 0; angryBirdLarge(107, 17) <= 0; angryBirdLarge(107, 18) <= 0; angryBirdLarge(107, 19) <= 0; angryBirdLarge(107, 20) <= 0; angryBirdLarge(107, 21) <= 0; angryBirdLarge(107, 22) <= 0; angryBirdLarge(107, 23) <= 0; angryBirdLarge(107, 24) <= 5; angryBirdLarge(107, 25) <= 5; angryBirdLarge(107, 26) <= 5; angryBirdLarge(107, 27) <= 5; angryBirdLarge(107, 28) <= 5; angryBirdLarge(107, 29) <= 5; angryBirdLarge(107, 30) <= 4; angryBirdLarge(107, 31) <= 4; angryBirdLarge(107, 32) <= 4; angryBirdLarge(107, 33) <= 4; angryBirdLarge(107, 34) <= 4; angryBirdLarge(107, 35) <= 4; angryBirdLarge(107, 36) <= 4; angryBirdLarge(107, 37) <= 4; angryBirdLarge(107, 38) <= 4; angryBirdLarge(107, 39) <= 4; angryBirdLarge(107, 40) <= 4; angryBirdLarge(107, 41) <= 4; angryBirdLarge(107, 42) <= 4; angryBirdLarge(107, 43) <= 4; angryBirdLarge(107, 44) <= 4; angryBirdLarge(107, 45) <= 4; angryBirdLarge(107, 46) <= 4; angryBirdLarge(107, 47) <= 4; angryBirdLarge(107, 48) <= 4; angryBirdLarge(107, 49) <= 4; angryBirdLarge(107, 50) <= 4; angryBirdLarge(107, 51) <= 4; angryBirdLarge(107, 52) <= 4; angryBirdLarge(107, 53) <= 4; angryBirdLarge(107, 54) <= 4; angryBirdLarge(107, 55) <= 4; angryBirdLarge(107, 56) <= 4; angryBirdLarge(107, 57) <= 4; angryBirdLarge(107, 58) <= 4; angryBirdLarge(107, 59) <= 4; angryBirdLarge(107, 60) <= 4; angryBirdLarge(107, 61) <= 4; angryBirdLarge(107, 62) <= 4; angryBirdLarge(107, 63) <= 4; angryBirdLarge(107, 64) <= 4; angryBirdLarge(107, 65) <= 4; angryBirdLarge(107, 66) <= 2; angryBirdLarge(107, 67) <= 2; angryBirdLarge(107, 68) <= 2; angryBirdLarge(107, 69) <= 2; angryBirdLarge(107, 70) <= 2; angryBirdLarge(107, 71) <= 2; angryBirdLarge(107, 72) <= 2; angryBirdLarge(107, 73) <= 2; angryBirdLarge(107, 74) <= 2; angryBirdLarge(107, 75) <= 2; angryBirdLarge(107, 76) <= 2; angryBirdLarge(107, 77) <= 2; angryBirdLarge(107, 78) <= 2; angryBirdLarge(107, 79) <= 2; angryBirdLarge(107, 80) <= 2; angryBirdLarge(107, 81) <= 2; angryBirdLarge(107, 82) <= 2; angryBirdLarge(107, 83) <= 2; angryBirdLarge(107, 84) <= 2; angryBirdLarge(107, 85) <= 2; angryBirdLarge(107, 86) <= 2; angryBirdLarge(107, 87) <= 2; angryBirdLarge(107, 88) <= 2; angryBirdLarge(107, 89) <= 2; angryBirdLarge(107, 90) <= 5; angryBirdLarge(107, 91) <= 5; angryBirdLarge(107, 92) <= 5; angryBirdLarge(107, 93) <= 5; angryBirdLarge(107, 94) <= 5; angryBirdLarge(107, 95) <= 5; angryBirdLarge(107, 96) <= 3; angryBirdLarge(107, 97) <= 3; angryBirdLarge(107, 98) <= 3; angryBirdLarge(107, 99) <= 3; angryBirdLarge(107, 100) <= 3; angryBirdLarge(107, 101) <= 3; angryBirdLarge(107, 102) <= 5; angryBirdLarge(107, 103) <= 5; angryBirdLarge(107, 104) <= 5; angryBirdLarge(107, 105) <= 5; angryBirdLarge(107, 106) <= 5; angryBirdLarge(107, 107) <= 5; angryBirdLarge(107, 108) <= 5; angryBirdLarge(107, 109) <= 5; angryBirdLarge(107, 110) <= 5; angryBirdLarge(107, 111) <= 5; angryBirdLarge(107, 112) <= 5; angryBirdLarge(107, 113) <= 5; angryBirdLarge(107, 114) <= 3; angryBirdLarge(107, 115) <= 3; angryBirdLarge(107, 116) <= 3; angryBirdLarge(107, 117) <= 3; angryBirdLarge(107, 118) <= 3; angryBirdLarge(107, 119) <= 3; angryBirdLarge(107, 120) <= 3; angryBirdLarge(107, 121) <= 3; angryBirdLarge(107, 122) <= 3; angryBirdLarge(107, 123) <= 3; angryBirdLarge(107, 124) <= 3; angryBirdLarge(107, 125) <= 3; angryBirdLarge(107, 126) <= 3; angryBirdLarge(107, 127) <= 3; angryBirdLarge(107, 128) <= 3; angryBirdLarge(107, 129) <= 3; angryBirdLarge(107, 130) <= 3; angryBirdLarge(107, 131) <= 3; angryBirdLarge(107, 132) <= 3; angryBirdLarge(107, 133) <= 3; angryBirdLarge(107, 134) <= 3; angryBirdLarge(107, 135) <= 3; angryBirdLarge(107, 136) <= 3; angryBirdLarge(107, 137) <= 3; angryBirdLarge(107, 138) <= 5; angryBirdLarge(107, 139) <= 5; angryBirdLarge(107, 140) <= 5; angryBirdLarge(107, 141) <= 5; angryBirdLarge(107, 142) <= 5; angryBirdLarge(107, 143) <= 5; angryBirdLarge(107, 144) <= 5; angryBirdLarge(107, 145) <= 5; angryBirdLarge(107, 146) <= 5; angryBirdLarge(107, 147) <= 5; angryBirdLarge(107, 148) <= 5; angryBirdLarge(107, 149) <= 5; 
angryBirdLarge(108, 0) <= 0; angryBirdLarge(108, 1) <= 0; angryBirdLarge(108, 2) <= 0; angryBirdLarge(108, 3) <= 0; angryBirdLarge(108, 4) <= 0; angryBirdLarge(108, 5) <= 0; angryBirdLarge(108, 6) <= 0; angryBirdLarge(108, 7) <= 0; angryBirdLarge(108, 8) <= 0; angryBirdLarge(108, 9) <= 0; angryBirdLarge(108, 10) <= 0; angryBirdLarge(108, 11) <= 0; angryBirdLarge(108, 12) <= 0; angryBirdLarge(108, 13) <= 0; angryBirdLarge(108, 14) <= 0; angryBirdLarge(108, 15) <= 0; angryBirdLarge(108, 16) <= 0; angryBirdLarge(108, 17) <= 0; angryBirdLarge(108, 18) <= 0; angryBirdLarge(108, 19) <= 0; angryBirdLarge(108, 20) <= 0; angryBirdLarge(108, 21) <= 0; angryBirdLarge(108, 22) <= 0; angryBirdLarge(108, 23) <= 0; angryBirdLarge(108, 24) <= 0; angryBirdLarge(108, 25) <= 0; angryBirdLarge(108, 26) <= 0; angryBirdLarge(108, 27) <= 0; angryBirdLarge(108, 28) <= 0; angryBirdLarge(108, 29) <= 0; angryBirdLarge(108, 30) <= 5; angryBirdLarge(108, 31) <= 5; angryBirdLarge(108, 32) <= 5; angryBirdLarge(108, 33) <= 5; angryBirdLarge(108, 34) <= 5; angryBirdLarge(108, 35) <= 5; angryBirdLarge(108, 36) <= 4; angryBirdLarge(108, 37) <= 4; angryBirdLarge(108, 38) <= 4; angryBirdLarge(108, 39) <= 4; angryBirdLarge(108, 40) <= 4; angryBirdLarge(108, 41) <= 4; angryBirdLarge(108, 42) <= 4; angryBirdLarge(108, 43) <= 4; angryBirdLarge(108, 44) <= 4; angryBirdLarge(108, 45) <= 4; angryBirdLarge(108, 46) <= 4; angryBirdLarge(108, 47) <= 4; angryBirdLarge(108, 48) <= 4; angryBirdLarge(108, 49) <= 4; angryBirdLarge(108, 50) <= 4; angryBirdLarge(108, 51) <= 4; angryBirdLarge(108, 52) <= 4; angryBirdLarge(108, 53) <= 4; angryBirdLarge(108, 54) <= 4; angryBirdLarge(108, 55) <= 4; angryBirdLarge(108, 56) <= 4; angryBirdLarge(108, 57) <= 4; angryBirdLarge(108, 58) <= 4; angryBirdLarge(108, 59) <= 4; angryBirdLarge(108, 60) <= 2; angryBirdLarge(108, 61) <= 2; angryBirdLarge(108, 62) <= 2; angryBirdLarge(108, 63) <= 2; angryBirdLarge(108, 64) <= 2; angryBirdLarge(108, 65) <= 2; angryBirdLarge(108, 66) <= 2; angryBirdLarge(108, 67) <= 2; angryBirdLarge(108, 68) <= 2; angryBirdLarge(108, 69) <= 2; angryBirdLarge(108, 70) <= 2; angryBirdLarge(108, 71) <= 2; angryBirdLarge(108, 72) <= 2; angryBirdLarge(108, 73) <= 2; angryBirdLarge(108, 74) <= 2; angryBirdLarge(108, 75) <= 2; angryBirdLarge(108, 76) <= 2; angryBirdLarge(108, 77) <= 2; angryBirdLarge(108, 78) <= 2; angryBirdLarge(108, 79) <= 2; angryBirdLarge(108, 80) <= 2; angryBirdLarge(108, 81) <= 2; angryBirdLarge(108, 82) <= 2; angryBirdLarge(108, 83) <= 2; angryBirdLarge(108, 84) <= 2; angryBirdLarge(108, 85) <= 2; angryBirdLarge(108, 86) <= 2; angryBirdLarge(108, 87) <= 2; angryBirdLarge(108, 88) <= 2; angryBirdLarge(108, 89) <= 2; angryBirdLarge(108, 90) <= 2; angryBirdLarge(108, 91) <= 2; angryBirdLarge(108, 92) <= 2; angryBirdLarge(108, 93) <= 2; angryBirdLarge(108, 94) <= 2; angryBirdLarge(108, 95) <= 2; angryBirdLarge(108, 96) <= 5; angryBirdLarge(108, 97) <= 5; angryBirdLarge(108, 98) <= 5; angryBirdLarge(108, 99) <= 5; angryBirdLarge(108, 100) <= 5; angryBirdLarge(108, 101) <= 5; angryBirdLarge(108, 102) <= 3; angryBirdLarge(108, 103) <= 3; angryBirdLarge(108, 104) <= 3; angryBirdLarge(108, 105) <= 3; angryBirdLarge(108, 106) <= 3; angryBirdLarge(108, 107) <= 3; angryBirdLarge(108, 108) <= 3; angryBirdLarge(108, 109) <= 3; angryBirdLarge(108, 110) <= 3; angryBirdLarge(108, 111) <= 3; angryBirdLarge(108, 112) <= 3; angryBirdLarge(108, 113) <= 3; angryBirdLarge(108, 114) <= 5; angryBirdLarge(108, 115) <= 5; angryBirdLarge(108, 116) <= 5; angryBirdLarge(108, 117) <= 5; angryBirdLarge(108, 118) <= 5; angryBirdLarge(108, 119) <= 5; angryBirdLarge(108, 120) <= 5; angryBirdLarge(108, 121) <= 5; angryBirdLarge(108, 122) <= 5; angryBirdLarge(108, 123) <= 5; angryBirdLarge(108, 124) <= 5; angryBirdLarge(108, 125) <= 5; angryBirdLarge(108, 126) <= 5; angryBirdLarge(108, 127) <= 5; angryBirdLarge(108, 128) <= 5; angryBirdLarge(108, 129) <= 5; angryBirdLarge(108, 130) <= 5; angryBirdLarge(108, 131) <= 5; angryBirdLarge(108, 132) <= 5; angryBirdLarge(108, 133) <= 5; angryBirdLarge(108, 134) <= 5; angryBirdLarge(108, 135) <= 5; angryBirdLarge(108, 136) <= 5; angryBirdLarge(108, 137) <= 5; angryBirdLarge(108, 138) <= 4; angryBirdLarge(108, 139) <= 4; angryBirdLarge(108, 140) <= 4; angryBirdLarge(108, 141) <= 4; angryBirdLarge(108, 142) <= 4; angryBirdLarge(108, 143) <= 4; angryBirdLarge(108, 144) <= 5; angryBirdLarge(108, 145) <= 5; angryBirdLarge(108, 146) <= 5; angryBirdLarge(108, 147) <= 5; angryBirdLarge(108, 148) <= 5; angryBirdLarge(108, 149) <= 5; 
angryBirdLarge(109, 0) <= 0; angryBirdLarge(109, 1) <= 0; angryBirdLarge(109, 2) <= 0; angryBirdLarge(109, 3) <= 0; angryBirdLarge(109, 4) <= 0; angryBirdLarge(109, 5) <= 0; angryBirdLarge(109, 6) <= 0; angryBirdLarge(109, 7) <= 0; angryBirdLarge(109, 8) <= 0; angryBirdLarge(109, 9) <= 0; angryBirdLarge(109, 10) <= 0; angryBirdLarge(109, 11) <= 0; angryBirdLarge(109, 12) <= 0; angryBirdLarge(109, 13) <= 0; angryBirdLarge(109, 14) <= 0; angryBirdLarge(109, 15) <= 0; angryBirdLarge(109, 16) <= 0; angryBirdLarge(109, 17) <= 0; angryBirdLarge(109, 18) <= 0; angryBirdLarge(109, 19) <= 0; angryBirdLarge(109, 20) <= 0; angryBirdLarge(109, 21) <= 0; angryBirdLarge(109, 22) <= 0; angryBirdLarge(109, 23) <= 0; angryBirdLarge(109, 24) <= 0; angryBirdLarge(109, 25) <= 0; angryBirdLarge(109, 26) <= 0; angryBirdLarge(109, 27) <= 0; angryBirdLarge(109, 28) <= 0; angryBirdLarge(109, 29) <= 0; angryBirdLarge(109, 30) <= 5; angryBirdLarge(109, 31) <= 5; angryBirdLarge(109, 32) <= 5; angryBirdLarge(109, 33) <= 5; angryBirdLarge(109, 34) <= 5; angryBirdLarge(109, 35) <= 5; angryBirdLarge(109, 36) <= 4; angryBirdLarge(109, 37) <= 4; angryBirdLarge(109, 38) <= 4; angryBirdLarge(109, 39) <= 4; angryBirdLarge(109, 40) <= 4; angryBirdLarge(109, 41) <= 4; angryBirdLarge(109, 42) <= 4; angryBirdLarge(109, 43) <= 4; angryBirdLarge(109, 44) <= 4; angryBirdLarge(109, 45) <= 4; angryBirdLarge(109, 46) <= 4; angryBirdLarge(109, 47) <= 4; angryBirdLarge(109, 48) <= 4; angryBirdLarge(109, 49) <= 4; angryBirdLarge(109, 50) <= 4; angryBirdLarge(109, 51) <= 4; angryBirdLarge(109, 52) <= 4; angryBirdLarge(109, 53) <= 4; angryBirdLarge(109, 54) <= 4; angryBirdLarge(109, 55) <= 4; angryBirdLarge(109, 56) <= 4; angryBirdLarge(109, 57) <= 4; angryBirdLarge(109, 58) <= 4; angryBirdLarge(109, 59) <= 4; angryBirdLarge(109, 60) <= 2; angryBirdLarge(109, 61) <= 2; angryBirdLarge(109, 62) <= 2; angryBirdLarge(109, 63) <= 2; angryBirdLarge(109, 64) <= 2; angryBirdLarge(109, 65) <= 2; angryBirdLarge(109, 66) <= 2; angryBirdLarge(109, 67) <= 2; angryBirdLarge(109, 68) <= 2; angryBirdLarge(109, 69) <= 2; angryBirdLarge(109, 70) <= 2; angryBirdLarge(109, 71) <= 2; angryBirdLarge(109, 72) <= 2; angryBirdLarge(109, 73) <= 2; angryBirdLarge(109, 74) <= 2; angryBirdLarge(109, 75) <= 2; angryBirdLarge(109, 76) <= 2; angryBirdLarge(109, 77) <= 2; angryBirdLarge(109, 78) <= 2; angryBirdLarge(109, 79) <= 2; angryBirdLarge(109, 80) <= 2; angryBirdLarge(109, 81) <= 2; angryBirdLarge(109, 82) <= 2; angryBirdLarge(109, 83) <= 2; angryBirdLarge(109, 84) <= 2; angryBirdLarge(109, 85) <= 2; angryBirdLarge(109, 86) <= 2; angryBirdLarge(109, 87) <= 2; angryBirdLarge(109, 88) <= 2; angryBirdLarge(109, 89) <= 2; angryBirdLarge(109, 90) <= 2; angryBirdLarge(109, 91) <= 2; angryBirdLarge(109, 92) <= 2; angryBirdLarge(109, 93) <= 2; angryBirdLarge(109, 94) <= 2; angryBirdLarge(109, 95) <= 2; angryBirdLarge(109, 96) <= 5; angryBirdLarge(109, 97) <= 5; angryBirdLarge(109, 98) <= 5; angryBirdLarge(109, 99) <= 5; angryBirdLarge(109, 100) <= 5; angryBirdLarge(109, 101) <= 5; angryBirdLarge(109, 102) <= 3; angryBirdLarge(109, 103) <= 3; angryBirdLarge(109, 104) <= 3; angryBirdLarge(109, 105) <= 3; angryBirdLarge(109, 106) <= 3; angryBirdLarge(109, 107) <= 3; angryBirdLarge(109, 108) <= 3; angryBirdLarge(109, 109) <= 3; angryBirdLarge(109, 110) <= 3; angryBirdLarge(109, 111) <= 3; angryBirdLarge(109, 112) <= 3; angryBirdLarge(109, 113) <= 3; angryBirdLarge(109, 114) <= 5; angryBirdLarge(109, 115) <= 5; angryBirdLarge(109, 116) <= 5; angryBirdLarge(109, 117) <= 5; angryBirdLarge(109, 118) <= 5; angryBirdLarge(109, 119) <= 5; angryBirdLarge(109, 120) <= 5; angryBirdLarge(109, 121) <= 5; angryBirdLarge(109, 122) <= 5; angryBirdLarge(109, 123) <= 5; angryBirdLarge(109, 124) <= 5; angryBirdLarge(109, 125) <= 5; angryBirdLarge(109, 126) <= 5; angryBirdLarge(109, 127) <= 5; angryBirdLarge(109, 128) <= 5; angryBirdLarge(109, 129) <= 5; angryBirdLarge(109, 130) <= 5; angryBirdLarge(109, 131) <= 5; angryBirdLarge(109, 132) <= 5; angryBirdLarge(109, 133) <= 5; angryBirdLarge(109, 134) <= 5; angryBirdLarge(109, 135) <= 5; angryBirdLarge(109, 136) <= 5; angryBirdLarge(109, 137) <= 5; angryBirdLarge(109, 138) <= 4; angryBirdLarge(109, 139) <= 4; angryBirdLarge(109, 140) <= 4; angryBirdLarge(109, 141) <= 4; angryBirdLarge(109, 142) <= 4; angryBirdLarge(109, 143) <= 4; angryBirdLarge(109, 144) <= 5; angryBirdLarge(109, 145) <= 5; angryBirdLarge(109, 146) <= 5; angryBirdLarge(109, 147) <= 5; angryBirdLarge(109, 148) <= 5; angryBirdLarge(109, 149) <= 5; 
angryBirdLarge(110, 0) <= 0; angryBirdLarge(110, 1) <= 0; angryBirdLarge(110, 2) <= 0; angryBirdLarge(110, 3) <= 0; angryBirdLarge(110, 4) <= 0; angryBirdLarge(110, 5) <= 0; angryBirdLarge(110, 6) <= 0; angryBirdLarge(110, 7) <= 0; angryBirdLarge(110, 8) <= 0; angryBirdLarge(110, 9) <= 0; angryBirdLarge(110, 10) <= 0; angryBirdLarge(110, 11) <= 0; angryBirdLarge(110, 12) <= 0; angryBirdLarge(110, 13) <= 0; angryBirdLarge(110, 14) <= 0; angryBirdLarge(110, 15) <= 0; angryBirdLarge(110, 16) <= 0; angryBirdLarge(110, 17) <= 0; angryBirdLarge(110, 18) <= 0; angryBirdLarge(110, 19) <= 0; angryBirdLarge(110, 20) <= 0; angryBirdLarge(110, 21) <= 0; angryBirdLarge(110, 22) <= 0; angryBirdLarge(110, 23) <= 0; angryBirdLarge(110, 24) <= 0; angryBirdLarge(110, 25) <= 0; angryBirdLarge(110, 26) <= 0; angryBirdLarge(110, 27) <= 0; angryBirdLarge(110, 28) <= 0; angryBirdLarge(110, 29) <= 0; angryBirdLarge(110, 30) <= 5; angryBirdLarge(110, 31) <= 5; angryBirdLarge(110, 32) <= 5; angryBirdLarge(110, 33) <= 5; angryBirdLarge(110, 34) <= 5; angryBirdLarge(110, 35) <= 5; angryBirdLarge(110, 36) <= 4; angryBirdLarge(110, 37) <= 4; angryBirdLarge(110, 38) <= 4; angryBirdLarge(110, 39) <= 4; angryBirdLarge(110, 40) <= 4; angryBirdLarge(110, 41) <= 4; angryBirdLarge(110, 42) <= 4; angryBirdLarge(110, 43) <= 4; angryBirdLarge(110, 44) <= 4; angryBirdLarge(110, 45) <= 4; angryBirdLarge(110, 46) <= 4; angryBirdLarge(110, 47) <= 4; angryBirdLarge(110, 48) <= 4; angryBirdLarge(110, 49) <= 4; angryBirdLarge(110, 50) <= 4; angryBirdLarge(110, 51) <= 4; angryBirdLarge(110, 52) <= 4; angryBirdLarge(110, 53) <= 4; angryBirdLarge(110, 54) <= 4; angryBirdLarge(110, 55) <= 4; angryBirdLarge(110, 56) <= 4; angryBirdLarge(110, 57) <= 4; angryBirdLarge(110, 58) <= 4; angryBirdLarge(110, 59) <= 4; angryBirdLarge(110, 60) <= 2; angryBirdLarge(110, 61) <= 2; angryBirdLarge(110, 62) <= 2; angryBirdLarge(110, 63) <= 2; angryBirdLarge(110, 64) <= 2; angryBirdLarge(110, 65) <= 2; angryBirdLarge(110, 66) <= 2; angryBirdLarge(110, 67) <= 2; angryBirdLarge(110, 68) <= 2; angryBirdLarge(110, 69) <= 2; angryBirdLarge(110, 70) <= 2; angryBirdLarge(110, 71) <= 2; angryBirdLarge(110, 72) <= 2; angryBirdLarge(110, 73) <= 2; angryBirdLarge(110, 74) <= 2; angryBirdLarge(110, 75) <= 2; angryBirdLarge(110, 76) <= 2; angryBirdLarge(110, 77) <= 2; angryBirdLarge(110, 78) <= 2; angryBirdLarge(110, 79) <= 2; angryBirdLarge(110, 80) <= 2; angryBirdLarge(110, 81) <= 2; angryBirdLarge(110, 82) <= 2; angryBirdLarge(110, 83) <= 2; angryBirdLarge(110, 84) <= 2; angryBirdLarge(110, 85) <= 2; angryBirdLarge(110, 86) <= 2; angryBirdLarge(110, 87) <= 2; angryBirdLarge(110, 88) <= 2; angryBirdLarge(110, 89) <= 2; angryBirdLarge(110, 90) <= 2; angryBirdLarge(110, 91) <= 2; angryBirdLarge(110, 92) <= 2; angryBirdLarge(110, 93) <= 2; angryBirdLarge(110, 94) <= 2; angryBirdLarge(110, 95) <= 2; angryBirdLarge(110, 96) <= 5; angryBirdLarge(110, 97) <= 5; angryBirdLarge(110, 98) <= 5; angryBirdLarge(110, 99) <= 5; angryBirdLarge(110, 100) <= 5; angryBirdLarge(110, 101) <= 5; angryBirdLarge(110, 102) <= 3; angryBirdLarge(110, 103) <= 3; angryBirdLarge(110, 104) <= 3; angryBirdLarge(110, 105) <= 3; angryBirdLarge(110, 106) <= 3; angryBirdLarge(110, 107) <= 3; angryBirdLarge(110, 108) <= 3; angryBirdLarge(110, 109) <= 3; angryBirdLarge(110, 110) <= 3; angryBirdLarge(110, 111) <= 3; angryBirdLarge(110, 112) <= 3; angryBirdLarge(110, 113) <= 3; angryBirdLarge(110, 114) <= 5; angryBirdLarge(110, 115) <= 5; angryBirdLarge(110, 116) <= 5; angryBirdLarge(110, 117) <= 5; angryBirdLarge(110, 118) <= 5; angryBirdLarge(110, 119) <= 5; angryBirdLarge(110, 120) <= 5; angryBirdLarge(110, 121) <= 5; angryBirdLarge(110, 122) <= 5; angryBirdLarge(110, 123) <= 5; angryBirdLarge(110, 124) <= 5; angryBirdLarge(110, 125) <= 5; angryBirdLarge(110, 126) <= 5; angryBirdLarge(110, 127) <= 5; angryBirdLarge(110, 128) <= 5; angryBirdLarge(110, 129) <= 5; angryBirdLarge(110, 130) <= 5; angryBirdLarge(110, 131) <= 5; angryBirdLarge(110, 132) <= 5; angryBirdLarge(110, 133) <= 5; angryBirdLarge(110, 134) <= 5; angryBirdLarge(110, 135) <= 5; angryBirdLarge(110, 136) <= 5; angryBirdLarge(110, 137) <= 5; angryBirdLarge(110, 138) <= 4; angryBirdLarge(110, 139) <= 4; angryBirdLarge(110, 140) <= 4; angryBirdLarge(110, 141) <= 4; angryBirdLarge(110, 142) <= 4; angryBirdLarge(110, 143) <= 4; angryBirdLarge(110, 144) <= 5; angryBirdLarge(110, 145) <= 5; angryBirdLarge(110, 146) <= 5; angryBirdLarge(110, 147) <= 5; angryBirdLarge(110, 148) <= 5; angryBirdLarge(110, 149) <= 5; 
angryBirdLarge(111, 0) <= 0; angryBirdLarge(111, 1) <= 0; angryBirdLarge(111, 2) <= 0; angryBirdLarge(111, 3) <= 0; angryBirdLarge(111, 4) <= 0; angryBirdLarge(111, 5) <= 0; angryBirdLarge(111, 6) <= 0; angryBirdLarge(111, 7) <= 0; angryBirdLarge(111, 8) <= 0; angryBirdLarge(111, 9) <= 0; angryBirdLarge(111, 10) <= 0; angryBirdLarge(111, 11) <= 0; angryBirdLarge(111, 12) <= 0; angryBirdLarge(111, 13) <= 0; angryBirdLarge(111, 14) <= 0; angryBirdLarge(111, 15) <= 0; angryBirdLarge(111, 16) <= 0; angryBirdLarge(111, 17) <= 0; angryBirdLarge(111, 18) <= 0; angryBirdLarge(111, 19) <= 0; angryBirdLarge(111, 20) <= 0; angryBirdLarge(111, 21) <= 0; angryBirdLarge(111, 22) <= 0; angryBirdLarge(111, 23) <= 0; angryBirdLarge(111, 24) <= 0; angryBirdLarge(111, 25) <= 0; angryBirdLarge(111, 26) <= 0; angryBirdLarge(111, 27) <= 0; angryBirdLarge(111, 28) <= 0; angryBirdLarge(111, 29) <= 0; angryBirdLarge(111, 30) <= 5; angryBirdLarge(111, 31) <= 5; angryBirdLarge(111, 32) <= 5; angryBirdLarge(111, 33) <= 5; angryBirdLarge(111, 34) <= 5; angryBirdLarge(111, 35) <= 5; angryBirdLarge(111, 36) <= 4; angryBirdLarge(111, 37) <= 4; angryBirdLarge(111, 38) <= 4; angryBirdLarge(111, 39) <= 4; angryBirdLarge(111, 40) <= 4; angryBirdLarge(111, 41) <= 4; angryBirdLarge(111, 42) <= 4; angryBirdLarge(111, 43) <= 4; angryBirdLarge(111, 44) <= 4; angryBirdLarge(111, 45) <= 4; angryBirdLarge(111, 46) <= 4; angryBirdLarge(111, 47) <= 4; angryBirdLarge(111, 48) <= 4; angryBirdLarge(111, 49) <= 4; angryBirdLarge(111, 50) <= 4; angryBirdLarge(111, 51) <= 4; angryBirdLarge(111, 52) <= 4; angryBirdLarge(111, 53) <= 4; angryBirdLarge(111, 54) <= 4; angryBirdLarge(111, 55) <= 4; angryBirdLarge(111, 56) <= 4; angryBirdLarge(111, 57) <= 4; angryBirdLarge(111, 58) <= 4; angryBirdLarge(111, 59) <= 4; angryBirdLarge(111, 60) <= 2; angryBirdLarge(111, 61) <= 2; angryBirdLarge(111, 62) <= 2; angryBirdLarge(111, 63) <= 2; angryBirdLarge(111, 64) <= 2; angryBirdLarge(111, 65) <= 2; angryBirdLarge(111, 66) <= 2; angryBirdLarge(111, 67) <= 2; angryBirdLarge(111, 68) <= 2; angryBirdLarge(111, 69) <= 2; angryBirdLarge(111, 70) <= 2; angryBirdLarge(111, 71) <= 2; angryBirdLarge(111, 72) <= 2; angryBirdLarge(111, 73) <= 2; angryBirdLarge(111, 74) <= 2; angryBirdLarge(111, 75) <= 2; angryBirdLarge(111, 76) <= 2; angryBirdLarge(111, 77) <= 2; angryBirdLarge(111, 78) <= 2; angryBirdLarge(111, 79) <= 2; angryBirdLarge(111, 80) <= 2; angryBirdLarge(111, 81) <= 2; angryBirdLarge(111, 82) <= 2; angryBirdLarge(111, 83) <= 2; angryBirdLarge(111, 84) <= 2; angryBirdLarge(111, 85) <= 2; angryBirdLarge(111, 86) <= 2; angryBirdLarge(111, 87) <= 2; angryBirdLarge(111, 88) <= 2; angryBirdLarge(111, 89) <= 2; angryBirdLarge(111, 90) <= 2; angryBirdLarge(111, 91) <= 2; angryBirdLarge(111, 92) <= 2; angryBirdLarge(111, 93) <= 2; angryBirdLarge(111, 94) <= 2; angryBirdLarge(111, 95) <= 2; angryBirdLarge(111, 96) <= 5; angryBirdLarge(111, 97) <= 5; angryBirdLarge(111, 98) <= 5; angryBirdLarge(111, 99) <= 5; angryBirdLarge(111, 100) <= 5; angryBirdLarge(111, 101) <= 5; angryBirdLarge(111, 102) <= 3; angryBirdLarge(111, 103) <= 3; angryBirdLarge(111, 104) <= 3; angryBirdLarge(111, 105) <= 3; angryBirdLarge(111, 106) <= 3; angryBirdLarge(111, 107) <= 3; angryBirdLarge(111, 108) <= 3; angryBirdLarge(111, 109) <= 3; angryBirdLarge(111, 110) <= 3; angryBirdLarge(111, 111) <= 3; angryBirdLarge(111, 112) <= 3; angryBirdLarge(111, 113) <= 3; angryBirdLarge(111, 114) <= 5; angryBirdLarge(111, 115) <= 5; angryBirdLarge(111, 116) <= 5; angryBirdLarge(111, 117) <= 5; angryBirdLarge(111, 118) <= 5; angryBirdLarge(111, 119) <= 5; angryBirdLarge(111, 120) <= 5; angryBirdLarge(111, 121) <= 5; angryBirdLarge(111, 122) <= 5; angryBirdLarge(111, 123) <= 5; angryBirdLarge(111, 124) <= 5; angryBirdLarge(111, 125) <= 5; angryBirdLarge(111, 126) <= 5; angryBirdLarge(111, 127) <= 5; angryBirdLarge(111, 128) <= 5; angryBirdLarge(111, 129) <= 5; angryBirdLarge(111, 130) <= 5; angryBirdLarge(111, 131) <= 5; angryBirdLarge(111, 132) <= 5; angryBirdLarge(111, 133) <= 5; angryBirdLarge(111, 134) <= 5; angryBirdLarge(111, 135) <= 5; angryBirdLarge(111, 136) <= 5; angryBirdLarge(111, 137) <= 5; angryBirdLarge(111, 138) <= 4; angryBirdLarge(111, 139) <= 4; angryBirdLarge(111, 140) <= 4; angryBirdLarge(111, 141) <= 4; angryBirdLarge(111, 142) <= 4; angryBirdLarge(111, 143) <= 4; angryBirdLarge(111, 144) <= 5; angryBirdLarge(111, 145) <= 5; angryBirdLarge(111, 146) <= 5; angryBirdLarge(111, 147) <= 5; angryBirdLarge(111, 148) <= 5; angryBirdLarge(111, 149) <= 5; 
angryBirdLarge(112, 0) <= 0; angryBirdLarge(112, 1) <= 0; angryBirdLarge(112, 2) <= 0; angryBirdLarge(112, 3) <= 0; angryBirdLarge(112, 4) <= 0; angryBirdLarge(112, 5) <= 0; angryBirdLarge(112, 6) <= 0; angryBirdLarge(112, 7) <= 0; angryBirdLarge(112, 8) <= 0; angryBirdLarge(112, 9) <= 0; angryBirdLarge(112, 10) <= 0; angryBirdLarge(112, 11) <= 0; angryBirdLarge(112, 12) <= 0; angryBirdLarge(112, 13) <= 0; angryBirdLarge(112, 14) <= 0; angryBirdLarge(112, 15) <= 0; angryBirdLarge(112, 16) <= 0; angryBirdLarge(112, 17) <= 0; angryBirdLarge(112, 18) <= 0; angryBirdLarge(112, 19) <= 0; angryBirdLarge(112, 20) <= 0; angryBirdLarge(112, 21) <= 0; angryBirdLarge(112, 22) <= 0; angryBirdLarge(112, 23) <= 0; angryBirdLarge(112, 24) <= 0; angryBirdLarge(112, 25) <= 0; angryBirdLarge(112, 26) <= 0; angryBirdLarge(112, 27) <= 0; angryBirdLarge(112, 28) <= 0; angryBirdLarge(112, 29) <= 0; angryBirdLarge(112, 30) <= 5; angryBirdLarge(112, 31) <= 5; angryBirdLarge(112, 32) <= 5; angryBirdLarge(112, 33) <= 5; angryBirdLarge(112, 34) <= 5; angryBirdLarge(112, 35) <= 5; angryBirdLarge(112, 36) <= 4; angryBirdLarge(112, 37) <= 4; angryBirdLarge(112, 38) <= 4; angryBirdLarge(112, 39) <= 4; angryBirdLarge(112, 40) <= 4; angryBirdLarge(112, 41) <= 4; angryBirdLarge(112, 42) <= 4; angryBirdLarge(112, 43) <= 4; angryBirdLarge(112, 44) <= 4; angryBirdLarge(112, 45) <= 4; angryBirdLarge(112, 46) <= 4; angryBirdLarge(112, 47) <= 4; angryBirdLarge(112, 48) <= 4; angryBirdLarge(112, 49) <= 4; angryBirdLarge(112, 50) <= 4; angryBirdLarge(112, 51) <= 4; angryBirdLarge(112, 52) <= 4; angryBirdLarge(112, 53) <= 4; angryBirdLarge(112, 54) <= 4; angryBirdLarge(112, 55) <= 4; angryBirdLarge(112, 56) <= 4; angryBirdLarge(112, 57) <= 4; angryBirdLarge(112, 58) <= 4; angryBirdLarge(112, 59) <= 4; angryBirdLarge(112, 60) <= 2; angryBirdLarge(112, 61) <= 2; angryBirdLarge(112, 62) <= 2; angryBirdLarge(112, 63) <= 2; angryBirdLarge(112, 64) <= 2; angryBirdLarge(112, 65) <= 2; angryBirdLarge(112, 66) <= 2; angryBirdLarge(112, 67) <= 2; angryBirdLarge(112, 68) <= 2; angryBirdLarge(112, 69) <= 2; angryBirdLarge(112, 70) <= 2; angryBirdLarge(112, 71) <= 2; angryBirdLarge(112, 72) <= 2; angryBirdLarge(112, 73) <= 2; angryBirdLarge(112, 74) <= 2; angryBirdLarge(112, 75) <= 2; angryBirdLarge(112, 76) <= 2; angryBirdLarge(112, 77) <= 2; angryBirdLarge(112, 78) <= 2; angryBirdLarge(112, 79) <= 2; angryBirdLarge(112, 80) <= 2; angryBirdLarge(112, 81) <= 2; angryBirdLarge(112, 82) <= 2; angryBirdLarge(112, 83) <= 2; angryBirdLarge(112, 84) <= 2; angryBirdLarge(112, 85) <= 2; angryBirdLarge(112, 86) <= 2; angryBirdLarge(112, 87) <= 2; angryBirdLarge(112, 88) <= 2; angryBirdLarge(112, 89) <= 2; angryBirdLarge(112, 90) <= 2; angryBirdLarge(112, 91) <= 2; angryBirdLarge(112, 92) <= 2; angryBirdLarge(112, 93) <= 2; angryBirdLarge(112, 94) <= 2; angryBirdLarge(112, 95) <= 2; angryBirdLarge(112, 96) <= 5; angryBirdLarge(112, 97) <= 5; angryBirdLarge(112, 98) <= 5; angryBirdLarge(112, 99) <= 5; angryBirdLarge(112, 100) <= 5; angryBirdLarge(112, 101) <= 5; angryBirdLarge(112, 102) <= 3; angryBirdLarge(112, 103) <= 3; angryBirdLarge(112, 104) <= 3; angryBirdLarge(112, 105) <= 3; angryBirdLarge(112, 106) <= 3; angryBirdLarge(112, 107) <= 3; angryBirdLarge(112, 108) <= 3; angryBirdLarge(112, 109) <= 3; angryBirdLarge(112, 110) <= 3; angryBirdLarge(112, 111) <= 3; angryBirdLarge(112, 112) <= 3; angryBirdLarge(112, 113) <= 3; angryBirdLarge(112, 114) <= 5; angryBirdLarge(112, 115) <= 5; angryBirdLarge(112, 116) <= 5; angryBirdLarge(112, 117) <= 5; angryBirdLarge(112, 118) <= 5; angryBirdLarge(112, 119) <= 5; angryBirdLarge(112, 120) <= 5; angryBirdLarge(112, 121) <= 5; angryBirdLarge(112, 122) <= 5; angryBirdLarge(112, 123) <= 5; angryBirdLarge(112, 124) <= 5; angryBirdLarge(112, 125) <= 5; angryBirdLarge(112, 126) <= 5; angryBirdLarge(112, 127) <= 5; angryBirdLarge(112, 128) <= 5; angryBirdLarge(112, 129) <= 5; angryBirdLarge(112, 130) <= 5; angryBirdLarge(112, 131) <= 5; angryBirdLarge(112, 132) <= 5; angryBirdLarge(112, 133) <= 5; angryBirdLarge(112, 134) <= 5; angryBirdLarge(112, 135) <= 5; angryBirdLarge(112, 136) <= 5; angryBirdLarge(112, 137) <= 5; angryBirdLarge(112, 138) <= 4; angryBirdLarge(112, 139) <= 4; angryBirdLarge(112, 140) <= 4; angryBirdLarge(112, 141) <= 4; angryBirdLarge(112, 142) <= 4; angryBirdLarge(112, 143) <= 4; angryBirdLarge(112, 144) <= 5; angryBirdLarge(112, 145) <= 5; angryBirdLarge(112, 146) <= 5; angryBirdLarge(112, 147) <= 5; angryBirdLarge(112, 148) <= 5; angryBirdLarge(112, 149) <= 5; 
angryBirdLarge(113, 0) <= 0; angryBirdLarge(113, 1) <= 0; angryBirdLarge(113, 2) <= 0; angryBirdLarge(113, 3) <= 0; angryBirdLarge(113, 4) <= 0; angryBirdLarge(113, 5) <= 0; angryBirdLarge(113, 6) <= 0; angryBirdLarge(113, 7) <= 0; angryBirdLarge(113, 8) <= 0; angryBirdLarge(113, 9) <= 0; angryBirdLarge(113, 10) <= 0; angryBirdLarge(113, 11) <= 0; angryBirdLarge(113, 12) <= 0; angryBirdLarge(113, 13) <= 0; angryBirdLarge(113, 14) <= 0; angryBirdLarge(113, 15) <= 0; angryBirdLarge(113, 16) <= 0; angryBirdLarge(113, 17) <= 0; angryBirdLarge(113, 18) <= 0; angryBirdLarge(113, 19) <= 0; angryBirdLarge(113, 20) <= 0; angryBirdLarge(113, 21) <= 0; angryBirdLarge(113, 22) <= 0; angryBirdLarge(113, 23) <= 0; angryBirdLarge(113, 24) <= 0; angryBirdLarge(113, 25) <= 0; angryBirdLarge(113, 26) <= 0; angryBirdLarge(113, 27) <= 0; angryBirdLarge(113, 28) <= 0; angryBirdLarge(113, 29) <= 0; angryBirdLarge(113, 30) <= 5; angryBirdLarge(113, 31) <= 5; angryBirdLarge(113, 32) <= 5; angryBirdLarge(113, 33) <= 5; angryBirdLarge(113, 34) <= 5; angryBirdLarge(113, 35) <= 5; angryBirdLarge(113, 36) <= 4; angryBirdLarge(113, 37) <= 4; angryBirdLarge(113, 38) <= 4; angryBirdLarge(113, 39) <= 4; angryBirdLarge(113, 40) <= 4; angryBirdLarge(113, 41) <= 4; angryBirdLarge(113, 42) <= 4; angryBirdLarge(113, 43) <= 4; angryBirdLarge(113, 44) <= 4; angryBirdLarge(113, 45) <= 4; angryBirdLarge(113, 46) <= 4; angryBirdLarge(113, 47) <= 4; angryBirdLarge(113, 48) <= 4; angryBirdLarge(113, 49) <= 4; angryBirdLarge(113, 50) <= 4; angryBirdLarge(113, 51) <= 4; angryBirdLarge(113, 52) <= 4; angryBirdLarge(113, 53) <= 4; angryBirdLarge(113, 54) <= 4; angryBirdLarge(113, 55) <= 4; angryBirdLarge(113, 56) <= 4; angryBirdLarge(113, 57) <= 4; angryBirdLarge(113, 58) <= 4; angryBirdLarge(113, 59) <= 4; angryBirdLarge(113, 60) <= 2; angryBirdLarge(113, 61) <= 2; angryBirdLarge(113, 62) <= 2; angryBirdLarge(113, 63) <= 2; angryBirdLarge(113, 64) <= 2; angryBirdLarge(113, 65) <= 2; angryBirdLarge(113, 66) <= 2; angryBirdLarge(113, 67) <= 2; angryBirdLarge(113, 68) <= 2; angryBirdLarge(113, 69) <= 2; angryBirdLarge(113, 70) <= 2; angryBirdLarge(113, 71) <= 2; angryBirdLarge(113, 72) <= 2; angryBirdLarge(113, 73) <= 2; angryBirdLarge(113, 74) <= 2; angryBirdLarge(113, 75) <= 2; angryBirdLarge(113, 76) <= 2; angryBirdLarge(113, 77) <= 2; angryBirdLarge(113, 78) <= 2; angryBirdLarge(113, 79) <= 2; angryBirdLarge(113, 80) <= 2; angryBirdLarge(113, 81) <= 2; angryBirdLarge(113, 82) <= 2; angryBirdLarge(113, 83) <= 2; angryBirdLarge(113, 84) <= 2; angryBirdLarge(113, 85) <= 2; angryBirdLarge(113, 86) <= 2; angryBirdLarge(113, 87) <= 2; angryBirdLarge(113, 88) <= 2; angryBirdLarge(113, 89) <= 2; angryBirdLarge(113, 90) <= 2; angryBirdLarge(113, 91) <= 2; angryBirdLarge(113, 92) <= 2; angryBirdLarge(113, 93) <= 2; angryBirdLarge(113, 94) <= 2; angryBirdLarge(113, 95) <= 2; angryBirdLarge(113, 96) <= 5; angryBirdLarge(113, 97) <= 5; angryBirdLarge(113, 98) <= 5; angryBirdLarge(113, 99) <= 5; angryBirdLarge(113, 100) <= 5; angryBirdLarge(113, 101) <= 5; angryBirdLarge(113, 102) <= 3; angryBirdLarge(113, 103) <= 3; angryBirdLarge(113, 104) <= 3; angryBirdLarge(113, 105) <= 3; angryBirdLarge(113, 106) <= 3; angryBirdLarge(113, 107) <= 3; angryBirdLarge(113, 108) <= 3; angryBirdLarge(113, 109) <= 3; angryBirdLarge(113, 110) <= 3; angryBirdLarge(113, 111) <= 3; angryBirdLarge(113, 112) <= 3; angryBirdLarge(113, 113) <= 3; angryBirdLarge(113, 114) <= 5; angryBirdLarge(113, 115) <= 5; angryBirdLarge(113, 116) <= 5; angryBirdLarge(113, 117) <= 5; angryBirdLarge(113, 118) <= 5; angryBirdLarge(113, 119) <= 5; angryBirdLarge(113, 120) <= 5; angryBirdLarge(113, 121) <= 5; angryBirdLarge(113, 122) <= 5; angryBirdLarge(113, 123) <= 5; angryBirdLarge(113, 124) <= 5; angryBirdLarge(113, 125) <= 5; angryBirdLarge(113, 126) <= 5; angryBirdLarge(113, 127) <= 5; angryBirdLarge(113, 128) <= 5; angryBirdLarge(113, 129) <= 5; angryBirdLarge(113, 130) <= 5; angryBirdLarge(113, 131) <= 5; angryBirdLarge(113, 132) <= 5; angryBirdLarge(113, 133) <= 5; angryBirdLarge(113, 134) <= 5; angryBirdLarge(113, 135) <= 5; angryBirdLarge(113, 136) <= 5; angryBirdLarge(113, 137) <= 5; angryBirdLarge(113, 138) <= 4; angryBirdLarge(113, 139) <= 4; angryBirdLarge(113, 140) <= 4; angryBirdLarge(113, 141) <= 4; angryBirdLarge(113, 142) <= 4; angryBirdLarge(113, 143) <= 4; angryBirdLarge(113, 144) <= 5; angryBirdLarge(113, 145) <= 5; angryBirdLarge(113, 146) <= 5; angryBirdLarge(113, 147) <= 5; angryBirdLarge(113, 148) <= 5; angryBirdLarge(113, 149) <= 5; 
angryBirdLarge(114, 0) <= 0; angryBirdLarge(114, 1) <= 0; angryBirdLarge(114, 2) <= 0; angryBirdLarge(114, 3) <= 0; angryBirdLarge(114, 4) <= 0; angryBirdLarge(114, 5) <= 0; angryBirdLarge(114, 6) <= 0; angryBirdLarge(114, 7) <= 0; angryBirdLarge(114, 8) <= 0; angryBirdLarge(114, 9) <= 0; angryBirdLarge(114, 10) <= 0; angryBirdLarge(114, 11) <= 0; angryBirdLarge(114, 12) <= 0; angryBirdLarge(114, 13) <= 0; angryBirdLarge(114, 14) <= 0; angryBirdLarge(114, 15) <= 0; angryBirdLarge(114, 16) <= 0; angryBirdLarge(114, 17) <= 0; angryBirdLarge(114, 18) <= 0; angryBirdLarge(114, 19) <= 0; angryBirdLarge(114, 20) <= 0; angryBirdLarge(114, 21) <= 0; angryBirdLarge(114, 22) <= 0; angryBirdLarge(114, 23) <= 0; angryBirdLarge(114, 24) <= 0; angryBirdLarge(114, 25) <= 0; angryBirdLarge(114, 26) <= 0; angryBirdLarge(114, 27) <= 0; angryBirdLarge(114, 28) <= 0; angryBirdLarge(114, 29) <= 0; angryBirdLarge(114, 30) <= 0; angryBirdLarge(114, 31) <= 0; angryBirdLarge(114, 32) <= 0; angryBirdLarge(114, 33) <= 0; angryBirdLarge(114, 34) <= 0; angryBirdLarge(114, 35) <= 0; angryBirdLarge(114, 36) <= 5; angryBirdLarge(114, 37) <= 5; angryBirdLarge(114, 38) <= 5; angryBirdLarge(114, 39) <= 5; angryBirdLarge(114, 40) <= 5; angryBirdLarge(114, 41) <= 5; angryBirdLarge(114, 42) <= 4; angryBirdLarge(114, 43) <= 4; angryBirdLarge(114, 44) <= 4; angryBirdLarge(114, 45) <= 4; angryBirdLarge(114, 46) <= 4; angryBirdLarge(114, 47) <= 4; angryBirdLarge(114, 48) <= 4; angryBirdLarge(114, 49) <= 4; angryBirdLarge(114, 50) <= 4; angryBirdLarge(114, 51) <= 4; angryBirdLarge(114, 52) <= 4; angryBirdLarge(114, 53) <= 4; angryBirdLarge(114, 54) <= 2; angryBirdLarge(114, 55) <= 2; angryBirdLarge(114, 56) <= 2; angryBirdLarge(114, 57) <= 2; angryBirdLarge(114, 58) <= 2; angryBirdLarge(114, 59) <= 2; angryBirdLarge(114, 60) <= 2; angryBirdLarge(114, 61) <= 2; angryBirdLarge(114, 62) <= 2; angryBirdLarge(114, 63) <= 2; angryBirdLarge(114, 64) <= 2; angryBirdLarge(114, 65) <= 2; angryBirdLarge(114, 66) <= 2; angryBirdLarge(114, 67) <= 2; angryBirdLarge(114, 68) <= 2; angryBirdLarge(114, 69) <= 2; angryBirdLarge(114, 70) <= 2; angryBirdLarge(114, 71) <= 2; angryBirdLarge(114, 72) <= 2; angryBirdLarge(114, 73) <= 2; angryBirdLarge(114, 74) <= 2; angryBirdLarge(114, 75) <= 2; angryBirdLarge(114, 76) <= 2; angryBirdLarge(114, 77) <= 2; angryBirdLarge(114, 78) <= 2; angryBirdLarge(114, 79) <= 2; angryBirdLarge(114, 80) <= 2; angryBirdLarge(114, 81) <= 2; angryBirdLarge(114, 82) <= 2; angryBirdLarge(114, 83) <= 2; angryBirdLarge(114, 84) <= 2; angryBirdLarge(114, 85) <= 2; angryBirdLarge(114, 86) <= 2; angryBirdLarge(114, 87) <= 2; angryBirdLarge(114, 88) <= 2; angryBirdLarge(114, 89) <= 2; angryBirdLarge(114, 90) <= 2; angryBirdLarge(114, 91) <= 2; angryBirdLarge(114, 92) <= 2; angryBirdLarge(114, 93) <= 2; angryBirdLarge(114, 94) <= 2; angryBirdLarge(114, 95) <= 2; angryBirdLarge(114, 96) <= 2; angryBirdLarge(114, 97) <= 2; angryBirdLarge(114, 98) <= 2; angryBirdLarge(114, 99) <= 2; angryBirdLarge(114, 100) <= 2; angryBirdLarge(114, 101) <= 2; angryBirdLarge(114, 102) <= 5; angryBirdLarge(114, 103) <= 5; angryBirdLarge(114, 104) <= 5; angryBirdLarge(114, 105) <= 5; angryBirdLarge(114, 106) <= 5; angryBirdLarge(114, 107) <= 5; angryBirdLarge(114, 108) <= 5; angryBirdLarge(114, 109) <= 5; angryBirdLarge(114, 110) <= 5; angryBirdLarge(114, 111) <= 5; angryBirdLarge(114, 112) <= 5; angryBirdLarge(114, 113) <= 5; angryBirdLarge(114, 114) <= 5; angryBirdLarge(114, 115) <= 5; angryBirdLarge(114, 116) <= 5; angryBirdLarge(114, 117) <= 5; angryBirdLarge(114, 118) <= 5; angryBirdLarge(114, 119) <= 5; angryBirdLarge(114, 120) <= 2; angryBirdLarge(114, 121) <= 2; angryBirdLarge(114, 122) <= 2; angryBirdLarge(114, 123) <= 2; angryBirdLarge(114, 124) <= 2; angryBirdLarge(114, 125) <= 2; angryBirdLarge(114, 126) <= 2; angryBirdLarge(114, 127) <= 2; angryBirdLarge(114, 128) <= 2; angryBirdLarge(114, 129) <= 2; angryBirdLarge(114, 130) <= 2; angryBirdLarge(114, 131) <= 2; angryBirdLarge(114, 132) <= 4; angryBirdLarge(114, 133) <= 4; angryBirdLarge(114, 134) <= 4; angryBirdLarge(114, 135) <= 4; angryBirdLarge(114, 136) <= 4; angryBirdLarge(114, 137) <= 4; angryBirdLarge(114, 138) <= 5; angryBirdLarge(114, 139) <= 5; angryBirdLarge(114, 140) <= 5; angryBirdLarge(114, 141) <= 5; angryBirdLarge(114, 142) <= 5; angryBirdLarge(114, 143) <= 5; angryBirdLarge(114, 144) <= 0; angryBirdLarge(114, 145) <= 0; angryBirdLarge(114, 146) <= 0; angryBirdLarge(114, 147) <= 0; angryBirdLarge(114, 148) <= 0; angryBirdLarge(114, 149) <= 0; 
angryBirdLarge(115, 0) <= 0; angryBirdLarge(115, 1) <= 0; angryBirdLarge(115, 2) <= 0; angryBirdLarge(115, 3) <= 0; angryBirdLarge(115, 4) <= 0; angryBirdLarge(115, 5) <= 0; angryBirdLarge(115, 6) <= 0; angryBirdLarge(115, 7) <= 0; angryBirdLarge(115, 8) <= 0; angryBirdLarge(115, 9) <= 0; angryBirdLarge(115, 10) <= 0; angryBirdLarge(115, 11) <= 0; angryBirdLarge(115, 12) <= 0; angryBirdLarge(115, 13) <= 0; angryBirdLarge(115, 14) <= 0; angryBirdLarge(115, 15) <= 0; angryBirdLarge(115, 16) <= 0; angryBirdLarge(115, 17) <= 0; angryBirdLarge(115, 18) <= 0; angryBirdLarge(115, 19) <= 0; angryBirdLarge(115, 20) <= 0; angryBirdLarge(115, 21) <= 0; angryBirdLarge(115, 22) <= 0; angryBirdLarge(115, 23) <= 0; angryBirdLarge(115, 24) <= 0; angryBirdLarge(115, 25) <= 0; angryBirdLarge(115, 26) <= 0; angryBirdLarge(115, 27) <= 0; angryBirdLarge(115, 28) <= 0; angryBirdLarge(115, 29) <= 0; angryBirdLarge(115, 30) <= 0; angryBirdLarge(115, 31) <= 0; angryBirdLarge(115, 32) <= 0; angryBirdLarge(115, 33) <= 0; angryBirdLarge(115, 34) <= 0; angryBirdLarge(115, 35) <= 0; angryBirdLarge(115, 36) <= 5; angryBirdLarge(115, 37) <= 5; angryBirdLarge(115, 38) <= 5; angryBirdLarge(115, 39) <= 5; angryBirdLarge(115, 40) <= 5; angryBirdLarge(115, 41) <= 5; angryBirdLarge(115, 42) <= 4; angryBirdLarge(115, 43) <= 4; angryBirdLarge(115, 44) <= 4; angryBirdLarge(115, 45) <= 4; angryBirdLarge(115, 46) <= 4; angryBirdLarge(115, 47) <= 4; angryBirdLarge(115, 48) <= 4; angryBirdLarge(115, 49) <= 4; angryBirdLarge(115, 50) <= 4; angryBirdLarge(115, 51) <= 4; angryBirdLarge(115, 52) <= 4; angryBirdLarge(115, 53) <= 4; angryBirdLarge(115, 54) <= 2; angryBirdLarge(115, 55) <= 2; angryBirdLarge(115, 56) <= 2; angryBirdLarge(115, 57) <= 2; angryBirdLarge(115, 58) <= 2; angryBirdLarge(115, 59) <= 2; angryBirdLarge(115, 60) <= 2; angryBirdLarge(115, 61) <= 2; angryBirdLarge(115, 62) <= 2; angryBirdLarge(115, 63) <= 2; angryBirdLarge(115, 64) <= 2; angryBirdLarge(115, 65) <= 2; angryBirdLarge(115, 66) <= 2; angryBirdLarge(115, 67) <= 2; angryBirdLarge(115, 68) <= 2; angryBirdLarge(115, 69) <= 2; angryBirdLarge(115, 70) <= 2; angryBirdLarge(115, 71) <= 2; angryBirdLarge(115, 72) <= 2; angryBirdLarge(115, 73) <= 2; angryBirdLarge(115, 74) <= 2; angryBirdLarge(115, 75) <= 2; angryBirdLarge(115, 76) <= 2; angryBirdLarge(115, 77) <= 2; angryBirdLarge(115, 78) <= 2; angryBirdLarge(115, 79) <= 2; angryBirdLarge(115, 80) <= 2; angryBirdLarge(115, 81) <= 2; angryBirdLarge(115, 82) <= 2; angryBirdLarge(115, 83) <= 2; angryBirdLarge(115, 84) <= 2; angryBirdLarge(115, 85) <= 2; angryBirdLarge(115, 86) <= 2; angryBirdLarge(115, 87) <= 2; angryBirdLarge(115, 88) <= 2; angryBirdLarge(115, 89) <= 2; angryBirdLarge(115, 90) <= 2; angryBirdLarge(115, 91) <= 2; angryBirdLarge(115, 92) <= 2; angryBirdLarge(115, 93) <= 2; angryBirdLarge(115, 94) <= 2; angryBirdLarge(115, 95) <= 2; angryBirdLarge(115, 96) <= 2; angryBirdLarge(115, 97) <= 2; angryBirdLarge(115, 98) <= 2; angryBirdLarge(115, 99) <= 2; angryBirdLarge(115, 100) <= 2; angryBirdLarge(115, 101) <= 2; angryBirdLarge(115, 102) <= 5; angryBirdLarge(115, 103) <= 5; angryBirdLarge(115, 104) <= 5; angryBirdLarge(115, 105) <= 5; angryBirdLarge(115, 106) <= 5; angryBirdLarge(115, 107) <= 5; angryBirdLarge(115, 108) <= 5; angryBirdLarge(115, 109) <= 5; angryBirdLarge(115, 110) <= 5; angryBirdLarge(115, 111) <= 5; angryBirdLarge(115, 112) <= 5; angryBirdLarge(115, 113) <= 5; angryBirdLarge(115, 114) <= 5; angryBirdLarge(115, 115) <= 5; angryBirdLarge(115, 116) <= 5; angryBirdLarge(115, 117) <= 5; angryBirdLarge(115, 118) <= 5; angryBirdLarge(115, 119) <= 5; angryBirdLarge(115, 120) <= 2; angryBirdLarge(115, 121) <= 2; angryBirdLarge(115, 122) <= 2; angryBirdLarge(115, 123) <= 2; angryBirdLarge(115, 124) <= 2; angryBirdLarge(115, 125) <= 2; angryBirdLarge(115, 126) <= 2; angryBirdLarge(115, 127) <= 2; angryBirdLarge(115, 128) <= 2; angryBirdLarge(115, 129) <= 2; angryBirdLarge(115, 130) <= 2; angryBirdLarge(115, 131) <= 2; angryBirdLarge(115, 132) <= 4; angryBirdLarge(115, 133) <= 4; angryBirdLarge(115, 134) <= 4; angryBirdLarge(115, 135) <= 4; angryBirdLarge(115, 136) <= 4; angryBirdLarge(115, 137) <= 4; angryBirdLarge(115, 138) <= 5; angryBirdLarge(115, 139) <= 5; angryBirdLarge(115, 140) <= 5; angryBirdLarge(115, 141) <= 5; angryBirdLarge(115, 142) <= 5; angryBirdLarge(115, 143) <= 5; angryBirdLarge(115, 144) <= 0; angryBirdLarge(115, 145) <= 0; angryBirdLarge(115, 146) <= 0; angryBirdLarge(115, 147) <= 0; angryBirdLarge(115, 148) <= 0; angryBirdLarge(115, 149) <= 0; 
angryBirdLarge(116, 0) <= 0; angryBirdLarge(116, 1) <= 0; angryBirdLarge(116, 2) <= 0; angryBirdLarge(116, 3) <= 0; angryBirdLarge(116, 4) <= 0; angryBirdLarge(116, 5) <= 0; angryBirdLarge(116, 6) <= 0; angryBirdLarge(116, 7) <= 0; angryBirdLarge(116, 8) <= 0; angryBirdLarge(116, 9) <= 0; angryBirdLarge(116, 10) <= 0; angryBirdLarge(116, 11) <= 0; angryBirdLarge(116, 12) <= 0; angryBirdLarge(116, 13) <= 0; angryBirdLarge(116, 14) <= 0; angryBirdLarge(116, 15) <= 0; angryBirdLarge(116, 16) <= 0; angryBirdLarge(116, 17) <= 0; angryBirdLarge(116, 18) <= 0; angryBirdLarge(116, 19) <= 0; angryBirdLarge(116, 20) <= 0; angryBirdLarge(116, 21) <= 0; angryBirdLarge(116, 22) <= 0; angryBirdLarge(116, 23) <= 0; angryBirdLarge(116, 24) <= 0; angryBirdLarge(116, 25) <= 0; angryBirdLarge(116, 26) <= 0; angryBirdLarge(116, 27) <= 0; angryBirdLarge(116, 28) <= 0; angryBirdLarge(116, 29) <= 0; angryBirdLarge(116, 30) <= 0; angryBirdLarge(116, 31) <= 0; angryBirdLarge(116, 32) <= 0; angryBirdLarge(116, 33) <= 0; angryBirdLarge(116, 34) <= 0; angryBirdLarge(116, 35) <= 0; angryBirdLarge(116, 36) <= 5; angryBirdLarge(116, 37) <= 5; angryBirdLarge(116, 38) <= 5; angryBirdLarge(116, 39) <= 5; angryBirdLarge(116, 40) <= 5; angryBirdLarge(116, 41) <= 5; angryBirdLarge(116, 42) <= 4; angryBirdLarge(116, 43) <= 4; angryBirdLarge(116, 44) <= 4; angryBirdLarge(116, 45) <= 4; angryBirdLarge(116, 46) <= 4; angryBirdLarge(116, 47) <= 4; angryBirdLarge(116, 48) <= 4; angryBirdLarge(116, 49) <= 4; angryBirdLarge(116, 50) <= 4; angryBirdLarge(116, 51) <= 4; angryBirdLarge(116, 52) <= 4; angryBirdLarge(116, 53) <= 4; angryBirdLarge(116, 54) <= 2; angryBirdLarge(116, 55) <= 2; angryBirdLarge(116, 56) <= 2; angryBirdLarge(116, 57) <= 2; angryBirdLarge(116, 58) <= 2; angryBirdLarge(116, 59) <= 2; angryBirdLarge(116, 60) <= 2; angryBirdLarge(116, 61) <= 2; angryBirdLarge(116, 62) <= 2; angryBirdLarge(116, 63) <= 2; angryBirdLarge(116, 64) <= 2; angryBirdLarge(116, 65) <= 2; angryBirdLarge(116, 66) <= 2; angryBirdLarge(116, 67) <= 2; angryBirdLarge(116, 68) <= 2; angryBirdLarge(116, 69) <= 2; angryBirdLarge(116, 70) <= 2; angryBirdLarge(116, 71) <= 2; angryBirdLarge(116, 72) <= 2; angryBirdLarge(116, 73) <= 2; angryBirdLarge(116, 74) <= 2; angryBirdLarge(116, 75) <= 2; angryBirdLarge(116, 76) <= 2; angryBirdLarge(116, 77) <= 2; angryBirdLarge(116, 78) <= 2; angryBirdLarge(116, 79) <= 2; angryBirdLarge(116, 80) <= 2; angryBirdLarge(116, 81) <= 2; angryBirdLarge(116, 82) <= 2; angryBirdLarge(116, 83) <= 2; angryBirdLarge(116, 84) <= 2; angryBirdLarge(116, 85) <= 2; angryBirdLarge(116, 86) <= 2; angryBirdLarge(116, 87) <= 2; angryBirdLarge(116, 88) <= 2; angryBirdLarge(116, 89) <= 2; angryBirdLarge(116, 90) <= 2; angryBirdLarge(116, 91) <= 2; angryBirdLarge(116, 92) <= 2; angryBirdLarge(116, 93) <= 2; angryBirdLarge(116, 94) <= 2; angryBirdLarge(116, 95) <= 2; angryBirdLarge(116, 96) <= 2; angryBirdLarge(116, 97) <= 2; angryBirdLarge(116, 98) <= 2; angryBirdLarge(116, 99) <= 2; angryBirdLarge(116, 100) <= 2; angryBirdLarge(116, 101) <= 2; angryBirdLarge(116, 102) <= 5; angryBirdLarge(116, 103) <= 5; angryBirdLarge(116, 104) <= 5; angryBirdLarge(116, 105) <= 5; angryBirdLarge(116, 106) <= 5; angryBirdLarge(116, 107) <= 5; angryBirdLarge(116, 108) <= 5; angryBirdLarge(116, 109) <= 5; angryBirdLarge(116, 110) <= 5; angryBirdLarge(116, 111) <= 5; angryBirdLarge(116, 112) <= 5; angryBirdLarge(116, 113) <= 5; angryBirdLarge(116, 114) <= 5; angryBirdLarge(116, 115) <= 5; angryBirdLarge(116, 116) <= 5; angryBirdLarge(116, 117) <= 5; angryBirdLarge(116, 118) <= 5; angryBirdLarge(116, 119) <= 5; angryBirdLarge(116, 120) <= 2; angryBirdLarge(116, 121) <= 2; angryBirdLarge(116, 122) <= 2; angryBirdLarge(116, 123) <= 2; angryBirdLarge(116, 124) <= 2; angryBirdLarge(116, 125) <= 2; angryBirdLarge(116, 126) <= 2; angryBirdLarge(116, 127) <= 2; angryBirdLarge(116, 128) <= 2; angryBirdLarge(116, 129) <= 2; angryBirdLarge(116, 130) <= 2; angryBirdLarge(116, 131) <= 2; angryBirdLarge(116, 132) <= 4; angryBirdLarge(116, 133) <= 4; angryBirdLarge(116, 134) <= 4; angryBirdLarge(116, 135) <= 4; angryBirdLarge(116, 136) <= 4; angryBirdLarge(116, 137) <= 4; angryBirdLarge(116, 138) <= 5; angryBirdLarge(116, 139) <= 5; angryBirdLarge(116, 140) <= 5; angryBirdLarge(116, 141) <= 5; angryBirdLarge(116, 142) <= 5; angryBirdLarge(116, 143) <= 5; angryBirdLarge(116, 144) <= 0; angryBirdLarge(116, 145) <= 0; angryBirdLarge(116, 146) <= 0; angryBirdLarge(116, 147) <= 0; angryBirdLarge(116, 148) <= 0; angryBirdLarge(116, 149) <= 0; 
angryBirdLarge(117, 0) <= 0; angryBirdLarge(117, 1) <= 0; angryBirdLarge(117, 2) <= 0; angryBirdLarge(117, 3) <= 0; angryBirdLarge(117, 4) <= 0; angryBirdLarge(117, 5) <= 0; angryBirdLarge(117, 6) <= 0; angryBirdLarge(117, 7) <= 0; angryBirdLarge(117, 8) <= 0; angryBirdLarge(117, 9) <= 0; angryBirdLarge(117, 10) <= 0; angryBirdLarge(117, 11) <= 0; angryBirdLarge(117, 12) <= 0; angryBirdLarge(117, 13) <= 0; angryBirdLarge(117, 14) <= 0; angryBirdLarge(117, 15) <= 0; angryBirdLarge(117, 16) <= 0; angryBirdLarge(117, 17) <= 0; angryBirdLarge(117, 18) <= 0; angryBirdLarge(117, 19) <= 0; angryBirdLarge(117, 20) <= 0; angryBirdLarge(117, 21) <= 0; angryBirdLarge(117, 22) <= 0; angryBirdLarge(117, 23) <= 0; angryBirdLarge(117, 24) <= 0; angryBirdLarge(117, 25) <= 0; angryBirdLarge(117, 26) <= 0; angryBirdLarge(117, 27) <= 0; angryBirdLarge(117, 28) <= 0; angryBirdLarge(117, 29) <= 0; angryBirdLarge(117, 30) <= 0; angryBirdLarge(117, 31) <= 0; angryBirdLarge(117, 32) <= 0; angryBirdLarge(117, 33) <= 0; angryBirdLarge(117, 34) <= 0; angryBirdLarge(117, 35) <= 0; angryBirdLarge(117, 36) <= 5; angryBirdLarge(117, 37) <= 5; angryBirdLarge(117, 38) <= 5; angryBirdLarge(117, 39) <= 5; angryBirdLarge(117, 40) <= 5; angryBirdLarge(117, 41) <= 5; angryBirdLarge(117, 42) <= 4; angryBirdLarge(117, 43) <= 4; angryBirdLarge(117, 44) <= 4; angryBirdLarge(117, 45) <= 4; angryBirdLarge(117, 46) <= 4; angryBirdLarge(117, 47) <= 4; angryBirdLarge(117, 48) <= 4; angryBirdLarge(117, 49) <= 4; angryBirdLarge(117, 50) <= 4; angryBirdLarge(117, 51) <= 4; angryBirdLarge(117, 52) <= 4; angryBirdLarge(117, 53) <= 4; angryBirdLarge(117, 54) <= 2; angryBirdLarge(117, 55) <= 2; angryBirdLarge(117, 56) <= 2; angryBirdLarge(117, 57) <= 2; angryBirdLarge(117, 58) <= 2; angryBirdLarge(117, 59) <= 2; angryBirdLarge(117, 60) <= 2; angryBirdLarge(117, 61) <= 2; angryBirdLarge(117, 62) <= 2; angryBirdLarge(117, 63) <= 2; angryBirdLarge(117, 64) <= 2; angryBirdLarge(117, 65) <= 2; angryBirdLarge(117, 66) <= 2; angryBirdLarge(117, 67) <= 2; angryBirdLarge(117, 68) <= 2; angryBirdLarge(117, 69) <= 2; angryBirdLarge(117, 70) <= 2; angryBirdLarge(117, 71) <= 2; angryBirdLarge(117, 72) <= 2; angryBirdLarge(117, 73) <= 2; angryBirdLarge(117, 74) <= 2; angryBirdLarge(117, 75) <= 2; angryBirdLarge(117, 76) <= 2; angryBirdLarge(117, 77) <= 2; angryBirdLarge(117, 78) <= 2; angryBirdLarge(117, 79) <= 2; angryBirdLarge(117, 80) <= 2; angryBirdLarge(117, 81) <= 2; angryBirdLarge(117, 82) <= 2; angryBirdLarge(117, 83) <= 2; angryBirdLarge(117, 84) <= 2; angryBirdLarge(117, 85) <= 2; angryBirdLarge(117, 86) <= 2; angryBirdLarge(117, 87) <= 2; angryBirdLarge(117, 88) <= 2; angryBirdLarge(117, 89) <= 2; angryBirdLarge(117, 90) <= 2; angryBirdLarge(117, 91) <= 2; angryBirdLarge(117, 92) <= 2; angryBirdLarge(117, 93) <= 2; angryBirdLarge(117, 94) <= 2; angryBirdLarge(117, 95) <= 2; angryBirdLarge(117, 96) <= 2; angryBirdLarge(117, 97) <= 2; angryBirdLarge(117, 98) <= 2; angryBirdLarge(117, 99) <= 2; angryBirdLarge(117, 100) <= 2; angryBirdLarge(117, 101) <= 2; angryBirdLarge(117, 102) <= 5; angryBirdLarge(117, 103) <= 5; angryBirdLarge(117, 104) <= 5; angryBirdLarge(117, 105) <= 5; angryBirdLarge(117, 106) <= 5; angryBirdLarge(117, 107) <= 5; angryBirdLarge(117, 108) <= 5; angryBirdLarge(117, 109) <= 5; angryBirdLarge(117, 110) <= 5; angryBirdLarge(117, 111) <= 5; angryBirdLarge(117, 112) <= 5; angryBirdLarge(117, 113) <= 5; angryBirdLarge(117, 114) <= 5; angryBirdLarge(117, 115) <= 5; angryBirdLarge(117, 116) <= 5; angryBirdLarge(117, 117) <= 5; angryBirdLarge(117, 118) <= 5; angryBirdLarge(117, 119) <= 5; angryBirdLarge(117, 120) <= 2; angryBirdLarge(117, 121) <= 2; angryBirdLarge(117, 122) <= 2; angryBirdLarge(117, 123) <= 2; angryBirdLarge(117, 124) <= 2; angryBirdLarge(117, 125) <= 2; angryBirdLarge(117, 126) <= 2; angryBirdLarge(117, 127) <= 2; angryBirdLarge(117, 128) <= 2; angryBirdLarge(117, 129) <= 2; angryBirdLarge(117, 130) <= 2; angryBirdLarge(117, 131) <= 2; angryBirdLarge(117, 132) <= 4; angryBirdLarge(117, 133) <= 4; angryBirdLarge(117, 134) <= 4; angryBirdLarge(117, 135) <= 4; angryBirdLarge(117, 136) <= 4; angryBirdLarge(117, 137) <= 4; angryBirdLarge(117, 138) <= 5; angryBirdLarge(117, 139) <= 5; angryBirdLarge(117, 140) <= 5; angryBirdLarge(117, 141) <= 5; angryBirdLarge(117, 142) <= 5; angryBirdLarge(117, 143) <= 5; angryBirdLarge(117, 144) <= 0; angryBirdLarge(117, 145) <= 0; angryBirdLarge(117, 146) <= 0; angryBirdLarge(117, 147) <= 0; angryBirdLarge(117, 148) <= 0; angryBirdLarge(117, 149) <= 0; 
angryBirdLarge(118, 0) <= 0; angryBirdLarge(118, 1) <= 0; angryBirdLarge(118, 2) <= 0; angryBirdLarge(118, 3) <= 0; angryBirdLarge(118, 4) <= 0; angryBirdLarge(118, 5) <= 0; angryBirdLarge(118, 6) <= 0; angryBirdLarge(118, 7) <= 0; angryBirdLarge(118, 8) <= 0; angryBirdLarge(118, 9) <= 0; angryBirdLarge(118, 10) <= 0; angryBirdLarge(118, 11) <= 0; angryBirdLarge(118, 12) <= 0; angryBirdLarge(118, 13) <= 0; angryBirdLarge(118, 14) <= 0; angryBirdLarge(118, 15) <= 0; angryBirdLarge(118, 16) <= 0; angryBirdLarge(118, 17) <= 0; angryBirdLarge(118, 18) <= 0; angryBirdLarge(118, 19) <= 0; angryBirdLarge(118, 20) <= 0; angryBirdLarge(118, 21) <= 0; angryBirdLarge(118, 22) <= 0; angryBirdLarge(118, 23) <= 0; angryBirdLarge(118, 24) <= 0; angryBirdLarge(118, 25) <= 0; angryBirdLarge(118, 26) <= 0; angryBirdLarge(118, 27) <= 0; angryBirdLarge(118, 28) <= 0; angryBirdLarge(118, 29) <= 0; angryBirdLarge(118, 30) <= 0; angryBirdLarge(118, 31) <= 0; angryBirdLarge(118, 32) <= 0; angryBirdLarge(118, 33) <= 0; angryBirdLarge(118, 34) <= 0; angryBirdLarge(118, 35) <= 0; angryBirdLarge(118, 36) <= 5; angryBirdLarge(118, 37) <= 5; angryBirdLarge(118, 38) <= 5; angryBirdLarge(118, 39) <= 5; angryBirdLarge(118, 40) <= 5; angryBirdLarge(118, 41) <= 5; angryBirdLarge(118, 42) <= 4; angryBirdLarge(118, 43) <= 4; angryBirdLarge(118, 44) <= 4; angryBirdLarge(118, 45) <= 4; angryBirdLarge(118, 46) <= 4; angryBirdLarge(118, 47) <= 4; angryBirdLarge(118, 48) <= 4; angryBirdLarge(118, 49) <= 4; angryBirdLarge(118, 50) <= 4; angryBirdLarge(118, 51) <= 4; angryBirdLarge(118, 52) <= 4; angryBirdLarge(118, 53) <= 4; angryBirdLarge(118, 54) <= 2; angryBirdLarge(118, 55) <= 2; angryBirdLarge(118, 56) <= 2; angryBirdLarge(118, 57) <= 2; angryBirdLarge(118, 58) <= 2; angryBirdLarge(118, 59) <= 2; angryBirdLarge(118, 60) <= 2; angryBirdLarge(118, 61) <= 2; angryBirdLarge(118, 62) <= 2; angryBirdLarge(118, 63) <= 2; angryBirdLarge(118, 64) <= 2; angryBirdLarge(118, 65) <= 2; angryBirdLarge(118, 66) <= 2; angryBirdLarge(118, 67) <= 2; angryBirdLarge(118, 68) <= 2; angryBirdLarge(118, 69) <= 2; angryBirdLarge(118, 70) <= 2; angryBirdLarge(118, 71) <= 2; angryBirdLarge(118, 72) <= 2; angryBirdLarge(118, 73) <= 2; angryBirdLarge(118, 74) <= 2; angryBirdLarge(118, 75) <= 2; angryBirdLarge(118, 76) <= 2; angryBirdLarge(118, 77) <= 2; angryBirdLarge(118, 78) <= 2; angryBirdLarge(118, 79) <= 2; angryBirdLarge(118, 80) <= 2; angryBirdLarge(118, 81) <= 2; angryBirdLarge(118, 82) <= 2; angryBirdLarge(118, 83) <= 2; angryBirdLarge(118, 84) <= 2; angryBirdLarge(118, 85) <= 2; angryBirdLarge(118, 86) <= 2; angryBirdLarge(118, 87) <= 2; angryBirdLarge(118, 88) <= 2; angryBirdLarge(118, 89) <= 2; angryBirdLarge(118, 90) <= 2; angryBirdLarge(118, 91) <= 2; angryBirdLarge(118, 92) <= 2; angryBirdLarge(118, 93) <= 2; angryBirdLarge(118, 94) <= 2; angryBirdLarge(118, 95) <= 2; angryBirdLarge(118, 96) <= 2; angryBirdLarge(118, 97) <= 2; angryBirdLarge(118, 98) <= 2; angryBirdLarge(118, 99) <= 2; angryBirdLarge(118, 100) <= 2; angryBirdLarge(118, 101) <= 2; angryBirdLarge(118, 102) <= 5; angryBirdLarge(118, 103) <= 5; angryBirdLarge(118, 104) <= 5; angryBirdLarge(118, 105) <= 5; angryBirdLarge(118, 106) <= 5; angryBirdLarge(118, 107) <= 5; angryBirdLarge(118, 108) <= 5; angryBirdLarge(118, 109) <= 5; angryBirdLarge(118, 110) <= 5; angryBirdLarge(118, 111) <= 5; angryBirdLarge(118, 112) <= 5; angryBirdLarge(118, 113) <= 5; angryBirdLarge(118, 114) <= 5; angryBirdLarge(118, 115) <= 5; angryBirdLarge(118, 116) <= 5; angryBirdLarge(118, 117) <= 5; angryBirdLarge(118, 118) <= 5; angryBirdLarge(118, 119) <= 5; angryBirdLarge(118, 120) <= 2; angryBirdLarge(118, 121) <= 2; angryBirdLarge(118, 122) <= 2; angryBirdLarge(118, 123) <= 2; angryBirdLarge(118, 124) <= 2; angryBirdLarge(118, 125) <= 2; angryBirdLarge(118, 126) <= 2; angryBirdLarge(118, 127) <= 2; angryBirdLarge(118, 128) <= 2; angryBirdLarge(118, 129) <= 2; angryBirdLarge(118, 130) <= 2; angryBirdLarge(118, 131) <= 2; angryBirdLarge(118, 132) <= 4; angryBirdLarge(118, 133) <= 4; angryBirdLarge(118, 134) <= 4; angryBirdLarge(118, 135) <= 4; angryBirdLarge(118, 136) <= 4; angryBirdLarge(118, 137) <= 4; angryBirdLarge(118, 138) <= 5; angryBirdLarge(118, 139) <= 5; angryBirdLarge(118, 140) <= 5; angryBirdLarge(118, 141) <= 5; angryBirdLarge(118, 142) <= 5; angryBirdLarge(118, 143) <= 5; angryBirdLarge(118, 144) <= 0; angryBirdLarge(118, 145) <= 0; angryBirdLarge(118, 146) <= 0; angryBirdLarge(118, 147) <= 0; angryBirdLarge(118, 148) <= 0; angryBirdLarge(118, 149) <= 0; 
angryBirdLarge(119, 0) <= 0; angryBirdLarge(119, 1) <= 0; angryBirdLarge(119, 2) <= 0; angryBirdLarge(119, 3) <= 0; angryBirdLarge(119, 4) <= 0; angryBirdLarge(119, 5) <= 0; angryBirdLarge(119, 6) <= 0; angryBirdLarge(119, 7) <= 0; angryBirdLarge(119, 8) <= 0; angryBirdLarge(119, 9) <= 0; angryBirdLarge(119, 10) <= 0; angryBirdLarge(119, 11) <= 0; angryBirdLarge(119, 12) <= 0; angryBirdLarge(119, 13) <= 0; angryBirdLarge(119, 14) <= 0; angryBirdLarge(119, 15) <= 0; angryBirdLarge(119, 16) <= 0; angryBirdLarge(119, 17) <= 0; angryBirdLarge(119, 18) <= 0; angryBirdLarge(119, 19) <= 0; angryBirdLarge(119, 20) <= 0; angryBirdLarge(119, 21) <= 0; angryBirdLarge(119, 22) <= 0; angryBirdLarge(119, 23) <= 0; angryBirdLarge(119, 24) <= 0; angryBirdLarge(119, 25) <= 0; angryBirdLarge(119, 26) <= 0; angryBirdLarge(119, 27) <= 0; angryBirdLarge(119, 28) <= 0; angryBirdLarge(119, 29) <= 0; angryBirdLarge(119, 30) <= 0; angryBirdLarge(119, 31) <= 0; angryBirdLarge(119, 32) <= 0; angryBirdLarge(119, 33) <= 0; angryBirdLarge(119, 34) <= 0; angryBirdLarge(119, 35) <= 0; angryBirdLarge(119, 36) <= 5; angryBirdLarge(119, 37) <= 5; angryBirdLarge(119, 38) <= 5; angryBirdLarge(119, 39) <= 5; angryBirdLarge(119, 40) <= 5; angryBirdLarge(119, 41) <= 5; angryBirdLarge(119, 42) <= 4; angryBirdLarge(119, 43) <= 4; angryBirdLarge(119, 44) <= 4; angryBirdLarge(119, 45) <= 4; angryBirdLarge(119, 46) <= 4; angryBirdLarge(119, 47) <= 4; angryBirdLarge(119, 48) <= 4; angryBirdLarge(119, 49) <= 4; angryBirdLarge(119, 50) <= 4; angryBirdLarge(119, 51) <= 4; angryBirdLarge(119, 52) <= 4; angryBirdLarge(119, 53) <= 4; angryBirdLarge(119, 54) <= 2; angryBirdLarge(119, 55) <= 2; angryBirdLarge(119, 56) <= 2; angryBirdLarge(119, 57) <= 2; angryBirdLarge(119, 58) <= 2; angryBirdLarge(119, 59) <= 2; angryBirdLarge(119, 60) <= 2; angryBirdLarge(119, 61) <= 2; angryBirdLarge(119, 62) <= 2; angryBirdLarge(119, 63) <= 2; angryBirdLarge(119, 64) <= 2; angryBirdLarge(119, 65) <= 2; angryBirdLarge(119, 66) <= 2; angryBirdLarge(119, 67) <= 2; angryBirdLarge(119, 68) <= 2; angryBirdLarge(119, 69) <= 2; angryBirdLarge(119, 70) <= 2; angryBirdLarge(119, 71) <= 2; angryBirdLarge(119, 72) <= 2; angryBirdLarge(119, 73) <= 2; angryBirdLarge(119, 74) <= 2; angryBirdLarge(119, 75) <= 2; angryBirdLarge(119, 76) <= 2; angryBirdLarge(119, 77) <= 2; angryBirdLarge(119, 78) <= 2; angryBirdLarge(119, 79) <= 2; angryBirdLarge(119, 80) <= 2; angryBirdLarge(119, 81) <= 2; angryBirdLarge(119, 82) <= 2; angryBirdLarge(119, 83) <= 2; angryBirdLarge(119, 84) <= 2; angryBirdLarge(119, 85) <= 2; angryBirdLarge(119, 86) <= 2; angryBirdLarge(119, 87) <= 2; angryBirdLarge(119, 88) <= 2; angryBirdLarge(119, 89) <= 2; angryBirdLarge(119, 90) <= 2; angryBirdLarge(119, 91) <= 2; angryBirdLarge(119, 92) <= 2; angryBirdLarge(119, 93) <= 2; angryBirdLarge(119, 94) <= 2; angryBirdLarge(119, 95) <= 2; angryBirdLarge(119, 96) <= 2; angryBirdLarge(119, 97) <= 2; angryBirdLarge(119, 98) <= 2; angryBirdLarge(119, 99) <= 2; angryBirdLarge(119, 100) <= 2; angryBirdLarge(119, 101) <= 2; angryBirdLarge(119, 102) <= 5; angryBirdLarge(119, 103) <= 5; angryBirdLarge(119, 104) <= 5; angryBirdLarge(119, 105) <= 5; angryBirdLarge(119, 106) <= 5; angryBirdLarge(119, 107) <= 5; angryBirdLarge(119, 108) <= 5; angryBirdLarge(119, 109) <= 5; angryBirdLarge(119, 110) <= 5; angryBirdLarge(119, 111) <= 5; angryBirdLarge(119, 112) <= 5; angryBirdLarge(119, 113) <= 5; angryBirdLarge(119, 114) <= 5; angryBirdLarge(119, 115) <= 5; angryBirdLarge(119, 116) <= 5; angryBirdLarge(119, 117) <= 5; angryBirdLarge(119, 118) <= 5; angryBirdLarge(119, 119) <= 5; angryBirdLarge(119, 120) <= 2; angryBirdLarge(119, 121) <= 2; angryBirdLarge(119, 122) <= 2; angryBirdLarge(119, 123) <= 2; angryBirdLarge(119, 124) <= 2; angryBirdLarge(119, 125) <= 2; angryBirdLarge(119, 126) <= 2; angryBirdLarge(119, 127) <= 2; angryBirdLarge(119, 128) <= 2; angryBirdLarge(119, 129) <= 2; angryBirdLarge(119, 130) <= 2; angryBirdLarge(119, 131) <= 2; angryBirdLarge(119, 132) <= 4; angryBirdLarge(119, 133) <= 4; angryBirdLarge(119, 134) <= 4; angryBirdLarge(119, 135) <= 4; angryBirdLarge(119, 136) <= 4; angryBirdLarge(119, 137) <= 4; angryBirdLarge(119, 138) <= 5; angryBirdLarge(119, 139) <= 5; angryBirdLarge(119, 140) <= 5; angryBirdLarge(119, 141) <= 5; angryBirdLarge(119, 142) <= 5; angryBirdLarge(119, 143) <= 5; angryBirdLarge(119, 144) <= 0; angryBirdLarge(119, 145) <= 0; angryBirdLarge(119, 146) <= 0; angryBirdLarge(119, 147) <= 0; angryBirdLarge(119, 148) <= 0; angryBirdLarge(119, 149) <= 0; 
angryBirdLarge(120, 0) <= 0; angryBirdLarge(120, 1) <= 0; angryBirdLarge(120, 2) <= 0; angryBirdLarge(120, 3) <= 0; angryBirdLarge(120, 4) <= 0; angryBirdLarge(120, 5) <= 0; angryBirdLarge(120, 6) <= 0; angryBirdLarge(120, 7) <= 0; angryBirdLarge(120, 8) <= 0; angryBirdLarge(120, 9) <= 0; angryBirdLarge(120, 10) <= 0; angryBirdLarge(120, 11) <= 0; angryBirdLarge(120, 12) <= 0; angryBirdLarge(120, 13) <= 0; angryBirdLarge(120, 14) <= 0; angryBirdLarge(120, 15) <= 0; angryBirdLarge(120, 16) <= 0; angryBirdLarge(120, 17) <= 0; angryBirdLarge(120, 18) <= 0; angryBirdLarge(120, 19) <= 0; angryBirdLarge(120, 20) <= 0; angryBirdLarge(120, 21) <= 0; angryBirdLarge(120, 22) <= 0; angryBirdLarge(120, 23) <= 0; angryBirdLarge(120, 24) <= 0; angryBirdLarge(120, 25) <= 0; angryBirdLarge(120, 26) <= 0; angryBirdLarge(120, 27) <= 0; angryBirdLarge(120, 28) <= 0; angryBirdLarge(120, 29) <= 0; angryBirdLarge(120, 30) <= 0; angryBirdLarge(120, 31) <= 0; angryBirdLarge(120, 32) <= 0; angryBirdLarge(120, 33) <= 0; angryBirdLarge(120, 34) <= 0; angryBirdLarge(120, 35) <= 0; angryBirdLarge(120, 36) <= 0; angryBirdLarge(120, 37) <= 0; angryBirdLarge(120, 38) <= 0; angryBirdLarge(120, 39) <= 0; angryBirdLarge(120, 40) <= 0; angryBirdLarge(120, 41) <= 0; angryBirdLarge(120, 42) <= 5; angryBirdLarge(120, 43) <= 5; angryBirdLarge(120, 44) <= 5; angryBirdLarge(120, 45) <= 5; angryBirdLarge(120, 46) <= 5; angryBirdLarge(120, 47) <= 5; angryBirdLarge(120, 48) <= 2; angryBirdLarge(120, 49) <= 2; angryBirdLarge(120, 50) <= 2; angryBirdLarge(120, 51) <= 2; angryBirdLarge(120, 52) <= 2; angryBirdLarge(120, 53) <= 2; angryBirdLarge(120, 54) <= 2; angryBirdLarge(120, 55) <= 2; angryBirdLarge(120, 56) <= 2; angryBirdLarge(120, 57) <= 2; angryBirdLarge(120, 58) <= 2; angryBirdLarge(120, 59) <= 2; angryBirdLarge(120, 60) <= 2; angryBirdLarge(120, 61) <= 2; angryBirdLarge(120, 62) <= 2; angryBirdLarge(120, 63) <= 2; angryBirdLarge(120, 64) <= 2; angryBirdLarge(120, 65) <= 2; angryBirdLarge(120, 66) <= 2; angryBirdLarge(120, 67) <= 2; angryBirdLarge(120, 68) <= 2; angryBirdLarge(120, 69) <= 2; angryBirdLarge(120, 70) <= 2; angryBirdLarge(120, 71) <= 2; angryBirdLarge(120, 72) <= 2; angryBirdLarge(120, 73) <= 2; angryBirdLarge(120, 74) <= 2; angryBirdLarge(120, 75) <= 2; angryBirdLarge(120, 76) <= 2; angryBirdLarge(120, 77) <= 2; angryBirdLarge(120, 78) <= 2; angryBirdLarge(120, 79) <= 2; angryBirdLarge(120, 80) <= 2; angryBirdLarge(120, 81) <= 2; angryBirdLarge(120, 82) <= 2; angryBirdLarge(120, 83) <= 2; angryBirdLarge(120, 84) <= 2; angryBirdLarge(120, 85) <= 2; angryBirdLarge(120, 86) <= 2; angryBirdLarge(120, 87) <= 2; angryBirdLarge(120, 88) <= 2; angryBirdLarge(120, 89) <= 2; angryBirdLarge(120, 90) <= 2; angryBirdLarge(120, 91) <= 2; angryBirdLarge(120, 92) <= 2; angryBirdLarge(120, 93) <= 2; angryBirdLarge(120, 94) <= 2; angryBirdLarge(120, 95) <= 2; angryBirdLarge(120, 96) <= 2; angryBirdLarge(120, 97) <= 2; angryBirdLarge(120, 98) <= 2; angryBirdLarge(120, 99) <= 2; angryBirdLarge(120, 100) <= 2; angryBirdLarge(120, 101) <= 2; angryBirdLarge(120, 102) <= 2; angryBirdLarge(120, 103) <= 2; angryBirdLarge(120, 104) <= 2; angryBirdLarge(120, 105) <= 2; angryBirdLarge(120, 106) <= 2; angryBirdLarge(120, 107) <= 2; angryBirdLarge(120, 108) <= 2; angryBirdLarge(120, 109) <= 2; angryBirdLarge(120, 110) <= 2; angryBirdLarge(120, 111) <= 2; angryBirdLarge(120, 112) <= 2; angryBirdLarge(120, 113) <= 2; angryBirdLarge(120, 114) <= 2; angryBirdLarge(120, 115) <= 2; angryBirdLarge(120, 116) <= 2; angryBirdLarge(120, 117) <= 2; angryBirdLarge(120, 118) <= 2; angryBirdLarge(120, 119) <= 2; angryBirdLarge(120, 120) <= 2; angryBirdLarge(120, 121) <= 2; angryBirdLarge(120, 122) <= 2; angryBirdLarge(120, 123) <= 2; angryBirdLarge(120, 124) <= 2; angryBirdLarge(120, 125) <= 2; angryBirdLarge(120, 126) <= 2; angryBirdLarge(120, 127) <= 2; angryBirdLarge(120, 128) <= 2; angryBirdLarge(120, 129) <= 2; angryBirdLarge(120, 130) <= 2; angryBirdLarge(120, 131) <= 2; angryBirdLarge(120, 132) <= 5; angryBirdLarge(120, 133) <= 5; angryBirdLarge(120, 134) <= 5; angryBirdLarge(120, 135) <= 5; angryBirdLarge(120, 136) <= 5; angryBirdLarge(120, 137) <= 5; angryBirdLarge(120, 138) <= 0; angryBirdLarge(120, 139) <= 0; angryBirdLarge(120, 140) <= 0; angryBirdLarge(120, 141) <= 0; angryBirdLarge(120, 142) <= 0; angryBirdLarge(120, 143) <= 0; angryBirdLarge(120, 144) <= 0; angryBirdLarge(120, 145) <= 0; angryBirdLarge(120, 146) <= 0; angryBirdLarge(120, 147) <= 0; angryBirdLarge(120, 148) <= 0; angryBirdLarge(120, 149) <= 0; 
angryBirdLarge(121, 0) <= 0; angryBirdLarge(121, 1) <= 0; angryBirdLarge(121, 2) <= 0; angryBirdLarge(121, 3) <= 0; angryBirdLarge(121, 4) <= 0; angryBirdLarge(121, 5) <= 0; angryBirdLarge(121, 6) <= 0; angryBirdLarge(121, 7) <= 0; angryBirdLarge(121, 8) <= 0; angryBirdLarge(121, 9) <= 0; angryBirdLarge(121, 10) <= 0; angryBirdLarge(121, 11) <= 0; angryBirdLarge(121, 12) <= 0; angryBirdLarge(121, 13) <= 0; angryBirdLarge(121, 14) <= 0; angryBirdLarge(121, 15) <= 0; angryBirdLarge(121, 16) <= 0; angryBirdLarge(121, 17) <= 0; angryBirdLarge(121, 18) <= 0; angryBirdLarge(121, 19) <= 0; angryBirdLarge(121, 20) <= 0; angryBirdLarge(121, 21) <= 0; angryBirdLarge(121, 22) <= 0; angryBirdLarge(121, 23) <= 0; angryBirdLarge(121, 24) <= 0; angryBirdLarge(121, 25) <= 0; angryBirdLarge(121, 26) <= 0; angryBirdLarge(121, 27) <= 0; angryBirdLarge(121, 28) <= 0; angryBirdLarge(121, 29) <= 0; angryBirdLarge(121, 30) <= 0; angryBirdLarge(121, 31) <= 0; angryBirdLarge(121, 32) <= 0; angryBirdLarge(121, 33) <= 0; angryBirdLarge(121, 34) <= 0; angryBirdLarge(121, 35) <= 0; angryBirdLarge(121, 36) <= 0; angryBirdLarge(121, 37) <= 0; angryBirdLarge(121, 38) <= 0; angryBirdLarge(121, 39) <= 0; angryBirdLarge(121, 40) <= 0; angryBirdLarge(121, 41) <= 0; angryBirdLarge(121, 42) <= 5; angryBirdLarge(121, 43) <= 5; angryBirdLarge(121, 44) <= 5; angryBirdLarge(121, 45) <= 5; angryBirdLarge(121, 46) <= 5; angryBirdLarge(121, 47) <= 5; angryBirdLarge(121, 48) <= 2; angryBirdLarge(121, 49) <= 2; angryBirdLarge(121, 50) <= 2; angryBirdLarge(121, 51) <= 2; angryBirdLarge(121, 52) <= 2; angryBirdLarge(121, 53) <= 2; angryBirdLarge(121, 54) <= 2; angryBirdLarge(121, 55) <= 2; angryBirdLarge(121, 56) <= 2; angryBirdLarge(121, 57) <= 2; angryBirdLarge(121, 58) <= 2; angryBirdLarge(121, 59) <= 2; angryBirdLarge(121, 60) <= 2; angryBirdLarge(121, 61) <= 2; angryBirdLarge(121, 62) <= 2; angryBirdLarge(121, 63) <= 2; angryBirdLarge(121, 64) <= 2; angryBirdLarge(121, 65) <= 2; angryBirdLarge(121, 66) <= 2; angryBirdLarge(121, 67) <= 2; angryBirdLarge(121, 68) <= 2; angryBirdLarge(121, 69) <= 2; angryBirdLarge(121, 70) <= 2; angryBirdLarge(121, 71) <= 2; angryBirdLarge(121, 72) <= 2; angryBirdLarge(121, 73) <= 2; angryBirdLarge(121, 74) <= 2; angryBirdLarge(121, 75) <= 2; angryBirdLarge(121, 76) <= 2; angryBirdLarge(121, 77) <= 2; angryBirdLarge(121, 78) <= 2; angryBirdLarge(121, 79) <= 2; angryBirdLarge(121, 80) <= 2; angryBirdLarge(121, 81) <= 2; angryBirdLarge(121, 82) <= 2; angryBirdLarge(121, 83) <= 2; angryBirdLarge(121, 84) <= 2; angryBirdLarge(121, 85) <= 2; angryBirdLarge(121, 86) <= 2; angryBirdLarge(121, 87) <= 2; angryBirdLarge(121, 88) <= 2; angryBirdLarge(121, 89) <= 2; angryBirdLarge(121, 90) <= 2; angryBirdLarge(121, 91) <= 2; angryBirdLarge(121, 92) <= 2; angryBirdLarge(121, 93) <= 2; angryBirdLarge(121, 94) <= 2; angryBirdLarge(121, 95) <= 2; angryBirdLarge(121, 96) <= 2; angryBirdLarge(121, 97) <= 2; angryBirdLarge(121, 98) <= 2; angryBirdLarge(121, 99) <= 2; angryBirdLarge(121, 100) <= 2; angryBirdLarge(121, 101) <= 2; angryBirdLarge(121, 102) <= 2; angryBirdLarge(121, 103) <= 2; angryBirdLarge(121, 104) <= 2; angryBirdLarge(121, 105) <= 2; angryBirdLarge(121, 106) <= 2; angryBirdLarge(121, 107) <= 2; angryBirdLarge(121, 108) <= 2; angryBirdLarge(121, 109) <= 2; angryBirdLarge(121, 110) <= 2; angryBirdLarge(121, 111) <= 2; angryBirdLarge(121, 112) <= 2; angryBirdLarge(121, 113) <= 2; angryBirdLarge(121, 114) <= 2; angryBirdLarge(121, 115) <= 2; angryBirdLarge(121, 116) <= 2; angryBirdLarge(121, 117) <= 2; angryBirdLarge(121, 118) <= 2; angryBirdLarge(121, 119) <= 2; angryBirdLarge(121, 120) <= 2; angryBirdLarge(121, 121) <= 2; angryBirdLarge(121, 122) <= 2; angryBirdLarge(121, 123) <= 2; angryBirdLarge(121, 124) <= 2; angryBirdLarge(121, 125) <= 2; angryBirdLarge(121, 126) <= 2; angryBirdLarge(121, 127) <= 2; angryBirdLarge(121, 128) <= 2; angryBirdLarge(121, 129) <= 2; angryBirdLarge(121, 130) <= 2; angryBirdLarge(121, 131) <= 2; angryBirdLarge(121, 132) <= 5; angryBirdLarge(121, 133) <= 5; angryBirdLarge(121, 134) <= 5; angryBirdLarge(121, 135) <= 5; angryBirdLarge(121, 136) <= 5; angryBirdLarge(121, 137) <= 5; angryBirdLarge(121, 138) <= 0; angryBirdLarge(121, 139) <= 0; angryBirdLarge(121, 140) <= 0; angryBirdLarge(121, 141) <= 0; angryBirdLarge(121, 142) <= 0; angryBirdLarge(121, 143) <= 0; angryBirdLarge(121, 144) <= 0; angryBirdLarge(121, 145) <= 0; angryBirdLarge(121, 146) <= 0; angryBirdLarge(121, 147) <= 0; angryBirdLarge(121, 148) <= 0; angryBirdLarge(121, 149) <= 0; 
angryBirdLarge(122, 0) <= 0; angryBirdLarge(122, 1) <= 0; angryBirdLarge(122, 2) <= 0; angryBirdLarge(122, 3) <= 0; angryBirdLarge(122, 4) <= 0; angryBirdLarge(122, 5) <= 0; angryBirdLarge(122, 6) <= 0; angryBirdLarge(122, 7) <= 0; angryBirdLarge(122, 8) <= 0; angryBirdLarge(122, 9) <= 0; angryBirdLarge(122, 10) <= 0; angryBirdLarge(122, 11) <= 0; angryBirdLarge(122, 12) <= 0; angryBirdLarge(122, 13) <= 0; angryBirdLarge(122, 14) <= 0; angryBirdLarge(122, 15) <= 0; angryBirdLarge(122, 16) <= 0; angryBirdLarge(122, 17) <= 0; angryBirdLarge(122, 18) <= 0; angryBirdLarge(122, 19) <= 0; angryBirdLarge(122, 20) <= 0; angryBirdLarge(122, 21) <= 0; angryBirdLarge(122, 22) <= 0; angryBirdLarge(122, 23) <= 0; angryBirdLarge(122, 24) <= 0; angryBirdLarge(122, 25) <= 0; angryBirdLarge(122, 26) <= 0; angryBirdLarge(122, 27) <= 0; angryBirdLarge(122, 28) <= 0; angryBirdLarge(122, 29) <= 0; angryBirdLarge(122, 30) <= 0; angryBirdLarge(122, 31) <= 0; angryBirdLarge(122, 32) <= 0; angryBirdLarge(122, 33) <= 0; angryBirdLarge(122, 34) <= 0; angryBirdLarge(122, 35) <= 0; angryBirdLarge(122, 36) <= 0; angryBirdLarge(122, 37) <= 0; angryBirdLarge(122, 38) <= 0; angryBirdLarge(122, 39) <= 0; angryBirdLarge(122, 40) <= 0; angryBirdLarge(122, 41) <= 0; angryBirdLarge(122, 42) <= 5; angryBirdLarge(122, 43) <= 5; angryBirdLarge(122, 44) <= 5; angryBirdLarge(122, 45) <= 5; angryBirdLarge(122, 46) <= 5; angryBirdLarge(122, 47) <= 5; angryBirdLarge(122, 48) <= 2; angryBirdLarge(122, 49) <= 2; angryBirdLarge(122, 50) <= 2; angryBirdLarge(122, 51) <= 2; angryBirdLarge(122, 52) <= 2; angryBirdLarge(122, 53) <= 2; angryBirdLarge(122, 54) <= 2; angryBirdLarge(122, 55) <= 2; angryBirdLarge(122, 56) <= 2; angryBirdLarge(122, 57) <= 2; angryBirdLarge(122, 58) <= 2; angryBirdLarge(122, 59) <= 2; angryBirdLarge(122, 60) <= 2; angryBirdLarge(122, 61) <= 2; angryBirdLarge(122, 62) <= 2; angryBirdLarge(122, 63) <= 2; angryBirdLarge(122, 64) <= 2; angryBirdLarge(122, 65) <= 2; angryBirdLarge(122, 66) <= 2; angryBirdLarge(122, 67) <= 2; angryBirdLarge(122, 68) <= 2; angryBirdLarge(122, 69) <= 2; angryBirdLarge(122, 70) <= 2; angryBirdLarge(122, 71) <= 2; angryBirdLarge(122, 72) <= 2; angryBirdLarge(122, 73) <= 2; angryBirdLarge(122, 74) <= 2; angryBirdLarge(122, 75) <= 2; angryBirdLarge(122, 76) <= 2; angryBirdLarge(122, 77) <= 2; angryBirdLarge(122, 78) <= 2; angryBirdLarge(122, 79) <= 2; angryBirdLarge(122, 80) <= 2; angryBirdLarge(122, 81) <= 2; angryBirdLarge(122, 82) <= 2; angryBirdLarge(122, 83) <= 2; angryBirdLarge(122, 84) <= 2; angryBirdLarge(122, 85) <= 2; angryBirdLarge(122, 86) <= 2; angryBirdLarge(122, 87) <= 2; angryBirdLarge(122, 88) <= 2; angryBirdLarge(122, 89) <= 2; angryBirdLarge(122, 90) <= 2; angryBirdLarge(122, 91) <= 2; angryBirdLarge(122, 92) <= 2; angryBirdLarge(122, 93) <= 2; angryBirdLarge(122, 94) <= 2; angryBirdLarge(122, 95) <= 2; angryBirdLarge(122, 96) <= 2; angryBirdLarge(122, 97) <= 2; angryBirdLarge(122, 98) <= 2; angryBirdLarge(122, 99) <= 2; angryBirdLarge(122, 100) <= 2; angryBirdLarge(122, 101) <= 2; angryBirdLarge(122, 102) <= 2; angryBirdLarge(122, 103) <= 2; angryBirdLarge(122, 104) <= 2; angryBirdLarge(122, 105) <= 2; angryBirdLarge(122, 106) <= 2; angryBirdLarge(122, 107) <= 2; angryBirdLarge(122, 108) <= 2; angryBirdLarge(122, 109) <= 2; angryBirdLarge(122, 110) <= 2; angryBirdLarge(122, 111) <= 2; angryBirdLarge(122, 112) <= 2; angryBirdLarge(122, 113) <= 2; angryBirdLarge(122, 114) <= 2; angryBirdLarge(122, 115) <= 2; angryBirdLarge(122, 116) <= 2; angryBirdLarge(122, 117) <= 2; angryBirdLarge(122, 118) <= 2; angryBirdLarge(122, 119) <= 2; angryBirdLarge(122, 120) <= 2; angryBirdLarge(122, 121) <= 2; angryBirdLarge(122, 122) <= 2; angryBirdLarge(122, 123) <= 2; angryBirdLarge(122, 124) <= 2; angryBirdLarge(122, 125) <= 2; angryBirdLarge(122, 126) <= 2; angryBirdLarge(122, 127) <= 2; angryBirdLarge(122, 128) <= 2; angryBirdLarge(122, 129) <= 2; angryBirdLarge(122, 130) <= 2; angryBirdLarge(122, 131) <= 2; angryBirdLarge(122, 132) <= 5; angryBirdLarge(122, 133) <= 5; angryBirdLarge(122, 134) <= 5; angryBirdLarge(122, 135) <= 5; angryBirdLarge(122, 136) <= 5; angryBirdLarge(122, 137) <= 5; angryBirdLarge(122, 138) <= 0; angryBirdLarge(122, 139) <= 0; angryBirdLarge(122, 140) <= 0; angryBirdLarge(122, 141) <= 0; angryBirdLarge(122, 142) <= 0; angryBirdLarge(122, 143) <= 0; angryBirdLarge(122, 144) <= 0; angryBirdLarge(122, 145) <= 0; angryBirdLarge(122, 146) <= 0; angryBirdLarge(122, 147) <= 0; angryBirdLarge(122, 148) <= 0; angryBirdLarge(122, 149) <= 0; 
angryBirdLarge(123, 0) <= 0; angryBirdLarge(123, 1) <= 0; angryBirdLarge(123, 2) <= 0; angryBirdLarge(123, 3) <= 0; angryBirdLarge(123, 4) <= 0; angryBirdLarge(123, 5) <= 0; angryBirdLarge(123, 6) <= 0; angryBirdLarge(123, 7) <= 0; angryBirdLarge(123, 8) <= 0; angryBirdLarge(123, 9) <= 0; angryBirdLarge(123, 10) <= 0; angryBirdLarge(123, 11) <= 0; angryBirdLarge(123, 12) <= 0; angryBirdLarge(123, 13) <= 0; angryBirdLarge(123, 14) <= 0; angryBirdLarge(123, 15) <= 0; angryBirdLarge(123, 16) <= 0; angryBirdLarge(123, 17) <= 0; angryBirdLarge(123, 18) <= 0; angryBirdLarge(123, 19) <= 0; angryBirdLarge(123, 20) <= 0; angryBirdLarge(123, 21) <= 0; angryBirdLarge(123, 22) <= 0; angryBirdLarge(123, 23) <= 0; angryBirdLarge(123, 24) <= 0; angryBirdLarge(123, 25) <= 0; angryBirdLarge(123, 26) <= 0; angryBirdLarge(123, 27) <= 0; angryBirdLarge(123, 28) <= 0; angryBirdLarge(123, 29) <= 0; angryBirdLarge(123, 30) <= 0; angryBirdLarge(123, 31) <= 0; angryBirdLarge(123, 32) <= 0; angryBirdLarge(123, 33) <= 0; angryBirdLarge(123, 34) <= 0; angryBirdLarge(123, 35) <= 0; angryBirdLarge(123, 36) <= 0; angryBirdLarge(123, 37) <= 0; angryBirdLarge(123, 38) <= 0; angryBirdLarge(123, 39) <= 0; angryBirdLarge(123, 40) <= 0; angryBirdLarge(123, 41) <= 0; angryBirdLarge(123, 42) <= 5; angryBirdLarge(123, 43) <= 5; angryBirdLarge(123, 44) <= 5; angryBirdLarge(123, 45) <= 5; angryBirdLarge(123, 46) <= 5; angryBirdLarge(123, 47) <= 5; angryBirdLarge(123, 48) <= 2; angryBirdLarge(123, 49) <= 2; angryBirdLarge(123, 50) <= 2; angryBirdLarge(123, 51) <= 2; angryBirdLarge(123, 52) <= 2; angryBirdLarge(123, 53) <= 2; angryBirdLarge(123, 54) <= 2; angryBirdLarge(123, 55) <= 2; angryBirdLarge(123, 56) <= 2; angryBirdLarge(123, 57) <= 2; angryBirdLarge(123, 58) <= 2; angryBirdLarge(123, 59) <= 2; angryBirdLarge(123, 60) <= 2; angryBirdLarge(123, 61) <= 2; angryBirdLarge(123, 62) <= 2; angryBirdLarge(123, 63) <= 2; angryBirdLarge(123, 64) <= 2; angryBirdLarge(123, 65) <= 2; angryBirdLarge(123, 66) <= 2; angryBirdLarge(123, 67) <= 2; angryBirdLarge(123, 68) <= 2; angryBirdLarge(123, 69) <= 2; angryBirdLarge(123, 70) <= 2; angryBirdLarge(123, 71) <= 2; angryBirdLarge(123, 72) <= 2; angryBirdLarge(123, 73) <= 2; angryBirdLarge(123, 74) <= 2; angryBirdLarge(123, 75) <= 2; angryBirdLarge(123, 76) <= 2; angryBirdLarge(123, 77) <= 2; angryBirdLarge(123, 78) <= 2; angryBirdLarge(123, 79) <= 2; angryBirdLarge(123, 80) <= 2; angryBirdLarge(123, 81) <= 2; angryBirdLarge(123, 82) <= 2; angryBirdLarge(123, 83) <= 2; angryBirdLarge(123, 84) <= 2; angryBirdLarge(123, 85) <= 2; angryBirdLarge(123, 86) <= 2; angryBirdLarge(123, 87) <= 2; angryBirdLarge(123, 88) <= 2; angryBirdLarge(123, 89) <= 2; angryBirdLarge(123, 90) <= 2; angryBirdLarge(123, 91) <= 2; angryBirdLarge(123, 92) <= 2; angryBirdLarge(123, 93) <= 2; angryBirdLarge(123, 94) <= 2; angryBirdLarge(123, 95) <= 2; angryBirdLarge(123, 96) <= 2; angryBirdLarge(123, 97) <= 2; angryBirdLarge(123, 98) <= 2; angryBirdLarge(123, 99) <= 2; angryBirdLarge(123, 100) <= 2; angryBirdLarge(123, 101) <= 2; angryBirdLarge(123, 102) <= 2; angryBirdLarge(123, 103) <= 2; angryBirdLarge(123, 104) <= 2; angryBirdLarge(123, 105) <= 2; angryBirdLarge(123, 106) <= 2; angryBirdLarge(123, 107) <= 2; angryBirdLarge(123, 108) <= 2; angryBirdLarge(123, 109) <= 2; angryBirdLarge(123, 110) <= 2; angryBirdLarge(123, 111) <= 2; angryBirdLarge(123, 112) <= 2; angryBirdLarge(123, 113) <= 2; angryBirdLarge(123, 114) <= 2; angryBirdLarge(123, 115) <= 2; angryBirdLarge(123, 116) <= 2; angryBirdLarge(123, 117) <= 2; angryBirdLarge(123, 118) <= 2; angryBirdLarge(123, 119) <= 2; angryBirdLarge(123, 120) <= 2; angryBirdLarge(123, 121) <= 2; angryBirdLarge(123, 122) <= 2; angryBirdLarge(123, 123) <= 2; angryBirdLarge(123, 124) <= 2; angryBirdLarge(123, 125) <= 2; angryBirdLarge(123, 126) <= 2; angryBirdLarge(123, 127) <= 2; angryBirdLarge(123, 128) <= 2; angryBirdLarge(123, 129) <= 2; angryBirdLarge(123, 130) <= 2; angryBirdLarge(123, 131) <= 2; angryBirdLarge(123, 132) <= 5; angryBirdLarge(123, 133) <= 5; angryBirdLarge(123, 134) <= 5; angryBirdLarge(123, 135) <= 5; angryBirdLarge(123, 136) <= 5; angryBirdLarge(123, 137) <= 5; angryBirdLarge(123, 138) <= 0; angryBirdLarge(123, 139) <= 0; angryBirdLarge(123, 140) <= 0; angryBirdLarge(123, 141) <= 0; angryBirdLarge(123, 142) <= 0; angryBirdLarge(123, 143) <= 0; angryBirdLarge(123, 144) <= 0; angryBirdLarge(123, 145) <= 0; angryBirdLarge(123, 146) <= 0; angryBirdLarge(123, 147) <= 0; angryBirdLarge(123, 148) <= 0; angryBirdLarge(123, 149) <= 0; 
angryBirdLarge(124, 0) <= 0; angryBirdLarge(124, 1) <= 0; angryBirdLarge(124, 2) <= 0; angryBirdLarge(124, 3) <= 0; angryBirdLarge(124, 4) <= 0; angryBirdLarge(124, 5) <= 0; angryBirdLarge(124, 6) <= 0; angryBirdLarge(124, 7) <= 0; angryBirdLarge(124, 8) <= 0; angryBirdLarge(124, 9) <= 0; angryBirdLarge(124, 10) <= 0; angryBirdLarge(124, 11) <= 0; angryBirdLarge(124, 12) <= 0; angryBirdLarge(124, 13) <= 0; angryBirdLarge(124, 14) <= 0; angryBirdLarge(124, 15) <= 0; angryBirdLarge(124, 16) <= 0; angryBirdLarge(124, 17) <= 0; angryBirdLarge(124, 18) <= 0; angryBirdLarge(124, 19) <= 0; angryBirdLarge(124, 20) <= 0; angryBirdLarge(124, 21) <= 0; angryBirdLarge(124, 22) <= 0; angryBirdLarge(124, 23) <= 0; angryBirdLarge(124, 24) <= 0; angryBirdLarge(124, 25) <= 0; angryBirdLarge(124, 26) <= 0; angryBirdLarge(124, 27) <= 0; angryBirdLarge(124, 28) <= 0; angryBirdLarge(124, 29) <= 0; angryBirdLarge(124, 30) <= 0; angryBirdLarge(124, 31) <= 0; angryBirdLarge(124, 32) <= 0; angryBirdLarge(124, 33) <= 0; angryBirdLarge(124, 34) <= 0; angryBirdLarge(124, 35) <= 0; angryBirdLarge(124, 36) <= 0; angryBirdLarge(124, 37) <= 0; angryBirdLarge(124, 38) <= 0; angryBirdLarge(124, 39) <= 0; angryBirdLarge(124, 40) <= 0; angryBirdLarge(124, 41) <= 0; angryBirdLarge(124, 42) <= 5; angryBirdLarge(124, 43) <= 5; angryBirdLarge(124, 44) <= 5; angryBirdLarge(124, 45) <= 5; angryBirdLarge(124, 46) <= 5; angryBirdLarge(124, 47) <= 5; angryBirdLarge(124, 48) <= 2; angryBirdLarge(124, 49) <= 2; angryBirdLarge(124, 50) <= 2; angryBirdLarge(124, 51) <= 2; angryBirdLarge(124, 52) <= 2; angryBirdLarge(124, 53) <= 2; angryBirdLarge(124, 54) <= 2; angryBirdLarge(124, 55) <= 2; angryBirdLarge(124, 56) <= 2; angryBirdLarge(124, 57) <= 2; angryBirdLarge(124, 58) <= 2; angryBirdLarge(124, 59) <= 2; angryBirdLarge(124, 60) <= 2; angryBirdLarge(124, 61) <= 2; angryBirdLarge(124, 62) <= 2; angryBirdLarge(124, 63) <= 2; angryBirdLarge(124, 64) <= 2; angryBirdLarge(124, 65) <= 2; angryBirdLarge(124, 66) <= 2; angryBirdLarge(124, 67) <= 2; angryBirdLarge(124, 68) <= 2; angryBirdLarge(124, 69) <= 2; angryBirdLarge(124, 70) <= 2; angryBirdLarge(124, 71) <= 2; angryBirdLarge(124, 72) <= 2; angryBirdLarge(124, 73) <= 2; angryBirdLarge(124, 74) <= 2; angryBirdLarge(124, 75) <= 2; angryBirdLarge(124, 76) <= 2; angryBirdLarge(124, 77) <= 2; angryBirdLarge(124, 78) <= 2; angryBirdLarge(124, 79) <= 2; angryBirdLarge(124, 80) <= 2; angryBirdLarge(124, 81) <= 2; angryBirdLarge(124, 82) <= 2; angryBirdLarge(124, 83) <= 2; angryBirdLarge(124, 84) <= 2; angryBirdLarge(124, 85) <= 2; angryBirdLarge(124, 86) <= 2; angryBirdLarge(124, 87) <= 2; angryBirdLarge(124, 88) <= 2; angryBirdLarge(124, 89) <= 2; angryBirdLarge(124, 90) <= 2; angryBirdLarge(124, 91) <= 2; angryBirdLarge(124, 92) <= 2; angryBirdLarge(124, 93) <= 2; angryBirdLarge(124, 94) <= 2; angryBirdLarge(124, 95) <= 2; angryBirdLarge(124, 96) <= 2; angryBirdLarge(124, 97) <= 2; angryBirdLarge(124, 98) <= 2; angryBirdLarge(124, 99) <= 2; angryBirdLarge(124, 100) <= 2; angryBirdLarge(124, 101) <= 2; angryBirdLarge(124, 102) <= 2; angryBirdLarge(124, 103) <= 2; angryBirdLarge(124, 104) <= 2; angryBirdLarge(124, 105) <= 2; angryBirdLarge(124, 106) <= 2; angryBirdLarge(124, 107) <= 2; angryBirdLarge(124, 108) <= 2; angryBirdLarge(124, 109) <= 2; angryBirdLarge(124, 110) <= 2; angryBirdLarge(124, 111) <= 2; angryBirdLarge(124, 112) <= 2; angryBirdLarge(124, 113) <= 2; angryBirdLarge(124, 114) <= 2; angryBirdLarge(124, 115) <= 2; angryBirdLarge(124, 116) <= 2; angryBirdLarge(124, 117) <= 2; angryBirdLarge(124, 118) <= 2; angryBirdLarge(124, 119) <= 2; angryBirdLarge(124, 120) <= 2; angryBirdLarge(124, 121) <= 2; angryBirdLarge(124, 122) <= 2; angryBirdLarge(124, 123) <= 2; angryBirdLarge(124, 124) <= 2; angryBirdLarge(124, 125) <= 2; angryBirdLarge(124, 126) <= 2; angryBirdLarge(124, 127) <= 2; angryBirdLarge(124, 128) <= 2; angryBirdLarge(124, 129) <= 2; angryBirdLarge(124, 130) <= 2; angryBirdLarge(124, 131) <= 2; angryBirdLarge(124, 132) <= 5; angryBirdLarge(124, 133) <= 5; angryBirdLarge(124, 134) <= 5; angryBirdLarge(124, 135) <= 5; angryBirdLarge(124, 136) <= 5; angryBirdLarge(124, 137) <= 5; angryBirdLarge(124, 138) <= 0; angryBirdLarge(124, 139) <= 0; angryBirdLarge(124, 140) <= 0; angryBirdLarge(124, 141) <= 0; angryBirdLarge(124, 142) <= 0; angryBirdLarge(124, 143) <= 0; angryBirdLarge(124, 144) <= 0; angryBirdLarge(124, 145) <= 0; angryBirdLarge(124, 146) <= 0; angryBirdLarge(124, 147) <= 0; angryBirdLarge(124, 148) <= 0; angryBirdLarge(124, 149) <= 0; 
angryBirdLarge(125, 0) <= 0; angryBirdLarge(125, 1) <= 0; angryBirdLarge(125, 2) <= 0; angryBirdLarge(125, 3) <= 0; angryBirdLarge(125, 4) <= 0; angryBirdLarge(125, 5) <= 0; angryBirdLarge(125, 6) <= 0; angryBirdLarge(125, 7) <= 0; angryBirdLarge(125, 8) <= 0; angryBirdLarge(125, 9) <= 0; angryBirdLarge(125, 10) <= 0; angryBirdLarge(125, 11) <= 0; angryBirdLarge(125, 12) <= 0; angryBirdLarge(125, 13) <= 0; angryBirdLarge(125, 14) <= 0; angryBirdLarge(125, 15) <= 0; angryBirdLarge(125, 16) <= 0; angryBirdLarge(125, 17) <= 0; angryBirdLarge(125, 18) <= 0; angryBirdLarge(125, 19) <= 0; angryBirdLarge(125, 20) <= 0; angryBirdLarge(125, 21) <= 0; angryBirdLarge(125, 22) <= 0; angryBirdLarge(125, 23) <= 0; angryBirdLarge(125, 24) <= 0; angryBirdLarge(125, 25) <= 0; angryBirdLarge(125, 26) <= 0; angryBirdLarge(125, 27) <= 0; angryBirdLarge(125, 28) <= 0; angryBirdLarge(125, 29) <= 0; angryBirdLarge(125, 30) <= 0; angryBirdLarge(125, 31) <= 0; angryBirdLarge(125, 32) <= 0; angryBirdLarge(125, 33) <= 0; angryBirdLarge(125, 34) <= 0; angryBirdLarge(125, 35) <= 0; angryBirdLarge(125, 36) <= 0; angryBirdLarge(125, 37) <= 0; angryBirdLarge(125, 38) <= 0; angryBirdLarge(125, 39) <= 0; angryBirdLarge(125, 40) <= 0; angryBirdLarge(125, 41) <= 0; angryBirdLarge(125, 42) <= 5; angryBirdLarge(125, 43) <= 5; angryBirdLarge(125, 44) <= 5; angryBirdLarge(125, 45) <= 5; angryBirdLarge(125, 46) <= 5; angryBirdLarge(125, 47) <= 5; angryBirdLarge(125, 48) <= 2; angryBirdLarge(125, 49) <= 2; angryBirdLarge(125, 50) <= 2; angryBirdLarge(125, 51) <= 2; angryBirdLarge(125, 52) <= 2; angryBirdLarge(125, 53) <= 2; angryBirdLarge(125, 54) <= 2; angryBirdLarge(125, 55) <= 2; angryBirdLarge(125, 56) <= 2; angryBirdLarge(125, 57) <= 2; angryBirdLarge(125, 58) <= 2; angryBirdLarge(125, 59) <= 2; angryBirdLarge(125, 60) <= 2; angryBirdLarge(125, 61) <= 2; angryBirdLarge(125, 62) <= 2; angryBirdLarge(125, 63) <= 2; angryBirdLarge(125, 64) <= 2; angryBirdLarge(125, 65) <= 2; angryBirdLarge(125, 66) <= 2; angryBirdLarge(125, 67) <= 2; angryBirdLarge(125, 68) <= 2; angryBirdLarge(125, 69) <= 2; angryBirdLarge(125, 70) <= 2; angryBirdLarge(125, 71) <= 2; angryBirdLarge(125, 72) <= 2; angryBirdLarge(125, 73) <= 2; angryBirdLarge(125, 74) <= 2; angryBirdLarge(125, 75) <= 2; angryBirdLarge(125, 76) <= 2; angryBirdLarge(125, 77) <= 2; angryBirdLarge(125, 78) <= 2; angryBirdLarge(125, 79) <= 2; angryBirdLarge(125, 80) <= 2; angryBirdLarge(125, 81) <= 2; angryBirdLarge(125, 82) <= 2; angryBirdLarge(125, 83) <= 2; angryBirdLarge(125, 84) <= 2; angryBirdLarge(125, 85) <= 2; angryBirdLarge(125, 86) <= 2; angryBirdLarge(125, 87) <= 2; angryBirdLarge(125, 88) <= 2; angryBirdLarge(125, 89) <= 2; angryBirdLarge(125, 90) <= 2; angryBirdLarge(125, 91) <= 2; angryBirdLarge(125, 92) <= 2; angryBirdLarge(125, 93) <= 2; angryBirdLarge(125, 94) <= 2; angryBirdLarge(125, 95) <= 2; angryBirdLarge(125, 96) <= 2; angryBirdLarge(125, 97) <= 2; angryBirdLarge(125, 98) <= 2; angryBirdLarge(125, 99) <= 2; angryBirdLarge(125, 100) <= 2; angryBirdLarge(125, 101) <= 2; angryBirdLarge(125, 102) <= 2; angryBirdLarge(125, 103) <= 2; angryBirdLarge(125, 104) <= 2; angryBirdLarge(125, 105) <= 2; angryBirdLarge(125, 106) <= 2; angryBirdLarge(125, 107) <= 2; angryBirdLarge(125, 108) <= 2; angryBirdLarge(125, 109) <= 2; angryBirdLarge(125, 110) <= 2; angryBirdLarge(125, 111) <= 2; angryBirdLarge(125, 112) <= 2; angryBirdLarge(125, 113) <= 2; angryBirdLarge(125, 114) <= 2; angryBirdLarge(125, 115) <= 2; angryBirdLarge(125, 116) <= 2; angryBirdLarge(125, 117) <= 2; angryBirdLarge(125, 118) <= 2; angryBirdLarge(125, 119) <= 2; angryBirdLarge(125, 120) <= 2; angryBirdLarge(125, 121) <= 2; angryBirdLarge(125, 122) <= 2; angryBirdLarge(125, 123) <= 2; angryBirdLarge(125, 124) <= 2; angryBirdLarge(125, 125) <= 2; angryBirdLarge(125, 126) <= 2; angryBirdLarge(125, 127) <= 2; angryBirdLarge(125, 128) <= 2; angryBirdLarge(125, 129) <= 2; angryBirdLarge(125, 130) <= 2; angryBirdLarge(125, 131) <= 2; angryBirdLarge(125, 132) <= 5; angryBirdLarge(125, 133) <= 5; angryBirdLarge(125, 134) <= 5; angryBirdLarge(125, 135) <= 5; angryBirdLarge(125, 136) <= 5; angryBirdLarge(125, 137) <= 5; angryBirdLarge(125, 138) <= 0; angryBirdLarge(125, 139) <= 0; angryBirdLarge(125, 140) <= 0; angryBirdLarge(125, 141) <= 0; angryBirdLarge(125, 142) <= 0; angryBirdLarge(125, 143) <= 0; angryBirdLarge(125, 144) <= 0; angryBirdLarge(125, 145) <= 0; angryBirdLarge(125, 146) <= 0; angryBirdLarge(125, 147) <= 0; angryBirdLarge(125, 148) <= 0; angryBirdLarge(125, 149) <= 0; 
angryBirdLarge(126, 0) <= 0; angryBirdLarge(126, 1) <= 0; angryBirdLarge(126, 2) <= 0; angryBirdLarge(126, 3) <= 0; angryBirdLarge(126, 4) <= 0; angryBirdLarge(126, 5) <= 0; angryBirdLarge(126, 6) <= 0; angryBirdLarge(126, 7) <= 0; angryBirdLarge(126, 8) <= 0; angryBirdLarge(126, 9) <= 0; angryBirdLarge(126, 10) <= 0; angryBirdLarge(126, 11) <= 0; angryBirdLarge(126, 12) <= 0; angryBirdLarge(126, 13) <= 0; angryBirdLarge(126, 14) <= 0; angryBirdLarge(126, 15) <= 0; angryBirdLarge(126, 16) <= 0; angryBirdLarge(126, 17) <= 0; angryBirdLarge(126, 18) <= 0; angryBirdLarge(126, 19) <= 0; angryBirdLarge(126, 20) <= 0; angryBirdLarge(126, 21) <= 0; angryBirdLarge(126, 22) <= 0; angryBirdLarge(126, 23) <= 0; angryBirdLarge(126, 24) <= 0; angryBirdLarge(126, 25) <= 0; angryBirdLarge(126, 26) <= 0; angryBirdLarge(126, 27) <= 0; angryBirdLarge(126, 28) <= 0; angryBirdLarge(126, 29) <= 0; angryBirdLarge(126, 30) <= 0; angryBirdLarge(126, 31) <= 0; angryBirdLarge(126, 32) <= 0; angryBirdLarge(126, 33) <= 0; angryBirdLarge(126, 34) <= 0; angryBirdLarge(126, 35) <= 0; angryBirdLarge(126, 36) <= 0; angryBirdLarge(126, 37) <= 0; angryBirdLarge(126, 38) <= 0; angryBirdLarge(126, 39) <= 0; angryBirdLarge(126, 40) <= 0; angryBirdLarge(126, 41) <= 0; angryBirdLarge(126, 42) <= 0; angryBirdLarge(126, 43) <= 0; angryBirdLarge(126, 44) <= 0; angryBirdLarge(126, 45) <= 0; angryBirdLarge(126, 46) <= 0; angryBirdLarge(126, 47) <= 0; angryBirdLarge(126, 48) <= 5; angryBirdLarge(126, 49) <= 5; angryBirdLarge(126, 50) <= 5; angryBirdLarge(126, 51) <= 5; angryBirdLarge(126, 52) <= 5; angryBirdLarge(126, 53) <= 5; angryBirdLarge(126, 54) <= 5; angryBirdLarge(126, 55) <= 5; angryBirdLarge(126, 56) <= 5; angryBirdLarge(126, 57) <= 5; angryBirdLarge(126, 58) <= 5; angryBirdLarge(126, 59) <= 5; angryBirdLarge(126, 60) <= 2; angryBirdLarge(126, 61) <= 2; angryBirdLarge(126, 62) <= 2; angryBirdLarge(126, 63) <= 2; angryBirdLarge(126, 64) <= 2; angryBirdLarge(126, 65) <= 2; angryBirdLarge(126, 66) <= 2; angryBirdLarge(126, 67) <= 2; angryBirdLarge(126, 68) <= 2; angryBirdLarge(126, 69) <= 2; angryBirdLarge(126, 70) <= 2; angryBirdLarge(126, 71) <= 2; angryBirdLarge(126, 72) <= 2; angryBirdLarge(126, 73) <= 2; angryBirdLarge(126, 74) <= 2; angryBirdLarge(126, 75) <= 2; angryBirdLarge(126, 76) <= 2; angryBirdLarge(126, 77) <= 2; angryBirdLarge(126, 78) <= 2; angryBirdLarge(126, 79) <= 2; angryBirdLarge(126, 80) <= 2; angryBirdLarge(126, 81) <= 2; angryBirdLarge(126, 82) <= 2; angryBirdLarge(126, 83) <= 2; angryBirdLarge(126, 84) <= 2; angryBirdLarge(126, 85) <= 2; angryBirdLarge(126, 86) <= 2; angryBirdLarge(126, 87) <= 2; angryBirdLarge(126, 88) <= 2; angryBirdLarge(126, 89) <= 2; angryBirdLarge(126, 90) <= 2; angryBirdLarge(126, 91) <= 2; angryBirdLarge(126, 92) <= 2; angryBirdLarge(126, 93) <= 2; angryBirdLarge(126, 94) <= 2; angryBirdLarge(126, 95) <= 2; angryBirdLarge(126, 96) <= 2; angryBirdLarge(126, 97) <= 2; angryBirdLarge(126, 98) <= 2; angryBirdLarge(126, 99) <= 2; angryBirdLarge(126, 100) <= 2; angryBirdLarge(126, 101) <= 2; angryBirdLarge(126, 102) <= 2; angryBirdLarge(126, 103) <= 2; angryBirdLarge(126, 104) <= 2; angryBirdLarge(126, 105) <= 2; angryBirdLarge(126, 106) <= 2; angryBirdLarge(126, 107) <= 2; angryBirdLarge(126, 108) <= 2; angryBirdLarge(126, 109) <= 2; angryBirdLarge(126, 110) <= 2; angryBirdLarge(126, 111) <= 2; angryBirdLarge(126, 112) <= 2; angryBirdLarge(126, 113) <= 2; angryBirdLarge(126, 114) <= 2; angryBirdLarge(126, 115) <= 2; angryBirdLarge(126, 116) <= 2; angryBirdLarge(126, 117) <= 2; angryBirdLarge(126, 118) <= 2; angryBirdLarge(126, 119) <= 2; angryBirdLarge(126, 120) <= 2; angryBirdLarge(126, 121) <= 2; angryBirdLarge(126, 122) <= 2; angryBirdLarge(126, 123) <= 2; angryBirdLarge(126, 124) <= 2; angryBirdLarge(126, 125) <= 2; angryBirdLarge(126, 126) <= 5; angryBirdLarge(126, 127) <= 5; angryBirdLarge(126, 128) <= 5; angryBirdLarge(126, 129) <= 5; angryBirdLarge(126, 130) <= 5; angryBirdLarge(126, 131) <= 5; angryBirdLarge(126, 132) <= 0; angryBirdLarge(126, 133) <= 0; angryBirdLarge(126, 134) <= 0; angryBirdLarge(126, 135) <= 0; angryBirdLarge(126, 136) <= 0; angryBirdLarge(126, 137) <= 0; angryBirdLarge(126, 138) <= 0; angryBirdLarge(126, 139) <= 0; angryBirdLarge(126, 140) <= 0; angryBirdLarge(126, 141) <= 0; angryBirdLarge(126, 142) <= 0; angryBirdLarge(126, 143) <= 0; angryBirdLarge(126, 144) <= 0; angryBirdLarge(126, 145) <= 0; angryBirdLarge(126, 146) <= 0; angryBirdLarge(126, 147) <= 0; angryBirdLarge(126, 148) <= 0; angryBirdLarge(126, 149) <= 0; 
angryBirdLarge(127, 0) <= 0; angryBirdLarge(127, 1) <= 0; angryBirdLarge(127, 2) <= 0; angryBirdLarge(127, 3) <= 0; angryBirdLarge(127, 4) <= 0; angryBirdLarge(127, 5) <= 0; angryBirdLarge(127, 6) <= 0; angryBirdLarge(127, 7) <= 0; angryBirdLarge(127, 8) <= 0; angryBirdLarge(127, 9) <= 0; angryBirdLarge(127, 10) <= 0; angryBirdLarge(127, 11) <= 0; angryBirdLarge(127, 12) <= 0; angryBirdLarge(127, 13) <= 0; angryBirdLarge(127, 14) <= 0; angryBirdLarge(127, 15) <= 0; angryBirdLarge(127, 16) <= 0; angryBirdLarge(127, 17) <= 0; angryBirdLarge(127, 18) <= 0; angryBirdLarge(127, 19) <= 0; angryBirdLarge(127, 20) <= 0; angryBirdLarge(127, 21) <= 0; angryBirdLarge(127, 22) <= 0; angryBirdLarge(127, 23) <= 0; angryBirdLarge(127, 24) <= 0; angryBirdLarge(127, 25) <= 0; angryBirdLarge(127, 26) <= 0; angryBirdLarge(127, 27) <= 0; angryBirdLarge(127, 28) <= 0; angryBirdLarge(127, 29) <= 0; angryBirdLarge(127, 30) <= 0; angryBirdLarge(127, 31) <= 0; angryBirdLarge(127, 32) <= 0; angryBirdLarge(127, 33) <= 0; angryBirdLarge(127, 34) <= 0; angryBirdLarge(127, 35) <= 0; angryBirdLarge(127, 36) <= 0; angryBirdLarge(127, 37) <= 0; angryBirdLarge(127, 38) <= 0; angryBirdLarge(127, 39) <= 0; angryBirdLarge(127, 40) <= 0; angryBirdLarge(127, 41) <= 0; angryBirdLarge(127, 42) <= 0; angryBirdLarge(127, 43) <= 0; angryBirdLarge(127, 44) <= 0; angryBirdLarge(127, 45) <= 0; angryBirdLarge(127, 46) <= 0; angryBirdLarge(127, 47) <= 0; angryBirdLarge(127, 48) <= 5; angryBirdLarge(127, 49) <= 5; angryBirdLarge(127, 50) <= 5; angryBirdLarge(127, 51) <= 5; angryBirdLarge(127, 52) <= 5; angryBirdLarge(127, 53) <= 5; angryBirdLarge(127, 54) <= 5; angryBirdLarge(127, 55) <= 5; angryBirdLarge(127, 56) <= 5; angryBirdLarge(127, 57) <= 5; angryBirdLarge(127, 58) <= 5; angryBirdLarge(127, 59) <= 5; angryBirdLarge(127, 60) <= 2; angryBirdLarge(127, 61) <= 2; angryBirdLarge(127, 62) <= 2; angryBirdLarge(127, 63) <= 2; angryBirdLarge(127, 64) <= 2; angryBirdLarge(127, 65) <= 2; angryBirdLarge(127, 66) <= 2; angryBirdLarge(127, 67) <= 2; angryBirdLarge(127, 68) <= 2; angryBirdLarge(127, 69) <= 2; angryBirdLarge(127, 70) <= 2; angryBirdLarge(127, 71) <= 2; angryBirdLarge(127, 72) <= 2; angryBirdLarge(127, 73) <= 2; angryBirdLarge(127, 74) <= 2; angryBirdLarge(127, 75) <= 2; angryBirdLarge(127, 76) <= 2; angryBirdLarge(127, 77) <= 2; angryBirdLarge(127, 78) <= 2; angryBirdLarge(127, 79) <= 2; angryBirdLarge(127, 80) <= 2; angryBirdLarge(127, 81) <= 2; angryBirdLarge(127, 82) <= 2; angryBirdLarge(127, 83) <= 2; angryBirdLarge(127, 84) <= 2; angryBirdLarge(127, 85) <= 2; angryBirdLarge(127, 86) <= 2; angryBirdLarge(127, 87) <= 2; angryBirdLarge(127, 88) <= 2; angryBirdLarge(127, 89) <= 2; angryBirdLarge(127, 90) <= 2; angryBirdLarge(127, 91) <= 2; angryBirdLarge(127, 92) <= 2; angryBirdLarge(127, 93) <= 2; angryBirdLarge(127, 94) <= 2; angryBirdLarge(127, 95) <= 2; angryBirdLarge(127, 96) <= 2; angryBirdLarge(127, 97) <= 2; angryBirdLarge(127, 98) <= 2; angryBirdLarge(127, 99) <= 2; angryBirdLarge(127, 100) <= 2; angryBirdLarge(127, 101) <= 2; angryBirdLarge(127, 102) <= 2; angryBirdLarge(127, 103) <= 2; angryBirdLarge(127, 104) <= 2; angryBirdLarge(127, 105) <= 2; angryBirdLarge(127, 106) <= 2; angryBirdLarge(127, 107) <= 2; angryBirdLarge(127, 108) <= 2; angryBirdLarge(127, 109) <= 2; angryBirdLarge(127, 110) <= 2; angryBirdLarge(127, 111) <= 2; angryBirdLarge(127, 112) <= 2; angryBirdLarge(127, 113) <= 2; angryBirdLarge(127, 114) <= 2; angryBirdLarge(127, 115) <= 2; angryBirdLarge(127, 116) <= 2; angryBirdLarge(127, 117) <= 2; angryBirdLarge(127, 118) <= 2; angryBirdLarge(127, 119) <= 2; angryBirdLarge(127, 120) <= 2; angryBirdLarge(127, 121) <= 2; angryBirdLarge(127, 122) <= 2; angryBirdLarge(127, 123) <= 2; angryBirdLarge(127, 124) <= 2; angryBirdLarge(127, 125) <= 2; angryBirdLarge(127, 126) <= 5; angryBirdLarge(127, 127) <= 5; angryBirdLarge(127, 128) <= 5; angryBirdLarge(127, 129) <= 5; angryBirdLarge(127, 130) <= 5; angryBirdLarge(127, 131) <= 5; angryBirdLarge(127, 132) <= 0; angryBirdLarge(127, 133) <= 0; angryBirdLarge(127, 134) <= 0; angryBirdLarge(127, 135) <= 0; angryBirdLarge(127, 136) <= 0; angryBirdLarge(127, 137) <= 0; angryBirdLarge(127, 138) <= 0; angryBirdLarge(127, 139) <= 0; angryBirdLarge(127, 140) <= 0; angryBirdLarge(127, 141) <= 0; angryBirdLarge(127, 142) <= 0; angryBirdLarge(127, 143) <= 0; angryBirdLarge(127, 144) <= 0; angryBirdLarge(127, 145) <= 0; angryBirdLarge(127, 146) <= 0; angryBirdLarge(127, 147) <= 0; angryBirdLarge(127, 148) <= 0; angryBirdLarge(127, 149) <= 0; 
angryBirdLarge(128, 0) <= 0; angryBirdLarge(128, 1) <= 0; angryBirdLarge(128, 2) <= 0; angryBirdLarge(128, 3) <= 0; angryBirdLarge(128, 4) <= 0; angryBirdLarge(128, 5) <= 0; angryBirdLarge(128, 6) <= 0; angryBirdLarge(128, 7) <= 0; angryBirdLarge(128, 8) <= 0; angryBirdLarge(128, 9) <= 0; angryBirdLarge(128, 10) <= 0; angryBirdLarge(128, 11) <= 0; angryBirdLarge(128, 12) <= 0; angryBirdLarge(128, 13) <= 0; angryBirdLarge(128, 14) <= 0; angryBirdLarge(128, 15) <= 0; angryBirdLarge(128, 16) <= 0; angryBirdLarge(128, 17) <= 0; angryBirdLarge(128, 18) <= 0; angryBirdLarge(128, 19) <= 0; angryBirdLarge(128, 20) <= 0; angryBirdLarge(128, 21) <= 0; angryBirdLarge(128, 22) <= 0; angryBirdLarge(128, 23) <= 0; angryBirdLarge(128, 24) <= 0; angryBirdLarge(128, 25) <= 0; angryBirdLarge(128, 26) <= 0; angryBirdLarge(128, 27) <= 0; angryBirdLarge(128, 28) <= 0; angryBirdLarge(128, 29) <= 0; angryBirdLarge(128, 30) <= 0; angryBirdLarge(128, 31) <= 0; angryBirdLarge(128, 32) <= 0; angryBirdLarge(128, 33) <= 0; angryBirdLarge(128, 34) <= 0; angryBirdLarge(128, 35) <= 0; angryBirdLarge(128, 36) <= 0; angryBirdLarge(128, 37) <= 0; angryBirdLarge(128, 38) <= 0; angryBirdLarge(128, 39) <= 0; angryBirdLarge(128, 40) <= 0; angryBirdLarge(128, 41) <= 0; angryBirdLarge(128, 42) <= 0; angryBirdLarge(128, 43) <= 0; angryBirdLarge(128, 44) <= 0; angryBirdLarge(128, 45) <= 0; angryBirdLarge(128, 46) <= 0; angryBirdLarge(128, 47) <= 0; angryBirdLarge(128, 48) <= 5; angryBirdLarge(128, 49) <= 5; angryBirdLarge(128, 50) <= 5; angryBirdLarge(128, 51) <= 5; angryBirdLarge(128, 52) <= 5; angryBirdLarge(128, 53) <= 5; angryBirdLarge(128, 54) <= 5; angryBirdLarge(128, 55) <= 5; angryBirdLarge(128, 56) <= 5; angryBirdLarge(128, 57) <= 5; angryBirdLarge(128, 58) <= 5; angryBirdLarge(128, 59) <= 5; angryBirdLarge(128, 60) <= 2; angryBirdLarge(128, 61) <= 2; angryBirdLarge(128, 62) <= 2; angryBirdLarge(128, 63) <= 2; angryBirdLarge(128, 64) <= 2; angryBirdLarge(128, 65) <= 2; angryBirdLarge(128, 66) <= 2; angryBirdLarge(128, 67) <= 2; angryBirdLarge(128, 68) <= 2; angryBirdLarge(128, 69) <= 2; angryBirdLarge(128, 70) <= 2; angryBirdLarge(128, 71) <= 2; angryBirdLarge(128, 72) <= 2; angryBirdLarge(128, 73) <= 2; angryBirdLarge(128, 74) <= 2; angryBirdLarge(128, 75) <= 2; angryBirdLarge(128, 76) <= 2; angryBirdLarge(128, 77) <= 2; angryBirdLarge(128, 78) <= 2; angryBirdLarge(128, 79) <= 2; angryBirdLarge(128, 80) <= 2; angryBirdLarge(128, 81) <= 2; angryBirdLarge(128, 82) <= 2; angryBirdLarge(128, 83) <= 2; angryBirdLarge(128, 84) <= 2; angryBirdLarge(128, 85) <= 2; angryBirdLarge(128, 86) <= 2; angryBirdLarge(128, 87) <= 2; angryBirdLarge(128, 88) <= 2; angryBirdLarge(128, 89) <= 2; angryBirdLarge(128, 90) <= 2; angryBirdLarge(128, 91) <= 2; angryBirdLarge(128, 92) <= 2; angryBirdLarge(128, 93) <= 2; angryBirdLarge(128, 94) <= 2; angryBirdLarge(128, 95) <= 2; angryBirdLarge(128, 96) <= 2; angryBirdLarge(128, 97) <= 2; angryBirdLarge(128, 98) <= 2; angryBirdLarge(128, 99) <= 2; angryBirdLarge(128, 100) <= 2; angryBirdLarge(128, 101) <= 2; angryBirdLarge(128, 102) <= 2; angryBirdLarge(128, 103) <= 2; angryBirdLarge(128, 104) <= 2; angryBirdLarge(128, 105) <= 2; angryBirdLarge(128, 106) <= 2; angryBirdLarge(128, 107) <= 2; angryBirdLarge(128, 108) <= 2; angryBirdLarge(128, 109) <= 2; angryBirdLarge(128, 110) <= 2; angryBirdLarge(128, 111) <= 2; angryBirdLarge(128, 112) <= 2; angryBirdLarge(128, 113) <= 2; angryBirdLarge(128, 114) <= 2; angryBirdLarge(128, 115) <= 2; angryBirdLarge(128, 116) <= 2; angryBirdLarge(128, 117) <= 2; angryBirdLarge(128, 118) <= 2; angryBirdLarge(128, 119) <= 2; angryBirdLarge(128, 120) <= 2; angryBirdLarge(128, 121) <= 2; angryBirdLarge(128, 122) <= 2; angryBirdLarge(128, 123) <= 2; angryBirdLarge(128, 124) <= 2; angryBirdLarge(128, 125) <= 2; angryBirdLarge(128, 126) <= 5; angryBirdLarge(128, 127) <= 5; angryBirdLarge(128, 128) <= 5; angryBirdLarge(128, 129) <= 5; angryBirdLarge(128, 130) <= 5; angryBirdLarge(128, 131) <= 5; angryBirdLarge(128, 132) <= 0; angryBirdLarge(128, 133) <= 0; angryBirdLarge(128, 134) <= 0; angryBirdLarge(128, 135) <= 0; angryBirdLarge(128, 136) <= 0; angryBirdLarge(128, 137) <= 0; angryBirdLarge(128, 138) <= 0; angryBirdLarge(128, 139) <= 0; angryBirdLarge(128, 140) <= 0; angryBirdLarge(128, 141) <= 0; angryBirdLarge(128, 142) <= 0; angryBirdLarge(128, 143) <= 0; angryBirdLarge(128, 144) <= 0; angryBirdLarge(128, 145) <= 0; angryBirdLarge(128, 146) <= 0; angryBirdLarge(128, 147) <= 0; angryBirdLarge(128, 148) <= 0; angryBirdLarge(128, 149) <= 0; 
angryBirdLarge(129, 0) <= 0; angryBirdLarge(129, 1) <= 0; angryBirdLarge(129, 2) <= 0; angryBirdLarge(129, 3) <= 0; angryBirdLarge(129, 4) <= 0; angryBirdLarge(129, 5) <= 0; angryBirdLarge(129, 6) <= 0; angryBirdLarge(129, 7) <= 0; angryBirdLarge(129, 8) <= 0; angryBirdLarge(129, 9) <= 0; angryBirdLarge(129, 10) <= 0; angryBirdLarge(129, 11) <= 0; angryBirdLarge(129, 12) <= 0; angryBirdLarge(129, 13) <= 0; angryBirdLarge(129, 14) <= 0; angryBirdLarge(129, 15) <= 0; angryBirdLarge(129, 16) <= 0; angryBirdLarge(129, 17) <= 0; angryBirdLarge(129, 18) <= 0; angryBirdLarge(129, 19) <= 0; angryBirdLarge(129, 20) <= 0; angryBirdLarge(129, 21) <= 0; angryBirdLarge(129, 22) <= 0; angryBirdLarge(129, 23) <= 0; angryBirdLarge(129, 24) <= 0; angryBirdLarge(129, 25) <= 0; angryBirdLarge(129, 26) <= 0; angryBirdLarge(129, 27) <= 0; angryBirdLarge(129, 28) <= 0; angryBirdLarge(129, 29) <= 0; angryBirdLarge(129, 30) <= 0; angryBirdLarge(129, 31) <= 0; angryBirdLarge(129, 32) <= 0; angryBirdLarge(129, 33) <= 0; angryBirdLarge(129, 34) <= 0; angryBirdLarge(129, 35) <= 0; angryBirdLarge(129, 36) <= 0; angryBirdLarge(129, 37) <= 0; angryBirdLarge(129, 38) <= 0; angryBirdLarge(129, 39) <= 0; angryBirdLarge(129, 40) <= 0; angryBirdLarge(129, 41) <= 0; angryBirdLarge(129, 42) <= 0; angryBirdLarge(129, 43) <= 0; angryBirdLarge(129, 44) <= 0; angryBirdLarge(129, 45) <= 0; angryBirdLarge(129, 46) <= 0; angryBirdLarge(129, 47) <= 0; angryBirdLarge(129, 48) <= 5; angryBirdLarge(129, 49) <= 5; angryBirdLarge(129, 50) <= 5; angryBirdLarge(129, 51) <= 5; angryBirdLarge(129, 52) <= 5; angryBirdLarge(129, 53) <= 5; angryBirdLarge(129, 54) <= 5; angryBirdLarge(129, 55) <= 5; angryBirdLarge(129, 56) <= 5; angryBirdLarge(129, 57) <= 5; angryBirdLarge(129, 58) <= 5; angryBirdLarge(129, 59) <= 5; angryBirdLarge(129, 60) <= 2; angryBirdLarge(129, 61) <= 2; angryBirdLarge(129, 62) <= 2; angryBirdLarge(129, 63) <= 2; angryBirdLarge(129, 64) <= 2; angryBirdLarge(129, 65) <= 2; angryBirdLarge(129, 66) <= 2; angryBirdLarge(129, 67) <= 2; angryBirdLarge(129, 68) <= 2; angryBirdLarge(129, 69) <= 2; angryBirdLarge(129, 70) <= 2; angryBirdLarge(129, 71) <= 2; angryBirdLarge(129, 72) <= 2; angryBirdLarge(129, 73) <= 2; angryBirdLarge(129, 74) <= 2; angryBirdLarge(129, 75) <= 2; angryBirdLarge(129, 76) <= 2; angryBirdLarge(129, 77) <= 2; angryBirdLarge(129, 78) <= 2; angryBirdLarge(129, 79) <= 2; angryBirdLarge(129, 80) <= 2; angryBirdLarge(129, 81) <= 2; angryBirdLarge(129, 82) <= 2; angryBirdLarge(129, 83) <= 2; angryBirdLarge(129, 84) <= 2; angryBirdLarge(129, 85) <= 2; angryBirdLarge(129, 86) <= 2; angryBirdLarge(129, 87) <= 2; angryBirdLarge(129, 88) <= 2; angryBirdLarge(129, 89) <= 2; angryBirdLarge(129, 90) <= 2; angryBirdLarge(129, 91) <= 2; angryBirdLarge(129, 92) <= 2; angryBirdLarge(129, 93) <= 2; angryBirdLarge(129, 94) <= 2; angryBirdLarge(129, 95) <= 2; angryBirdLarge(129, 96) <= 2; angryBirdLarge(129, 97) <= 2; angryBirdLarge(129, 98) <= 2; angryBirdLarge(129, 99) <= 2; angryBirdLarge(129, 100) <= 2; angryBirdLarge(129, 101) <= 2; angryBirdLarge(129, 102) <= 2; angryBirdLarge(129, 103) <= 2; angryBirdLarge(129, 104) <= 2; angryBirdLarge(129, 105) <= 2; angryBirdLarge(129, 106) <= 2; angryBirdLarge(129, 107) <= 2; angryBirdLarge(129, 108) <= 2; angryBirdLarge(129, 109) <= 2; angryBirdLarge(129, 110) <= 2; angryBirdLarge(129, 111) <= 2; angryBirdLarge(129, 112) <= 2; angryBirdLarge(129, 113) <= 2; angryBirdLarge(129, 114) <= 2; angryBirdLarge(129, 115) <= 2; angryBirdLarge(129, 116) <= 2; angryBirdLarge(129, 117) <= 2; angryBirdLarge(129, 118) <= 2; angryBirdLarge(129, 119) <= 2; angryBirdLarge(129, 120) <= 2; angryBirdLarge(129, 121) <= 2; angryBirdLarge(129, 122) <= 2; angryBirdLarge(129, 123) <= 2; angryBirdLarge(129, 124) <= 2; angryBirdLarge(129, 125) <= 2; angryBirdLarge(129, 126) <= 5; angryBirdLarge(129, 127) <= 5; angryBirdLarge(129, 128) <= 5; angryBirdLarge(129, 129) <= 5; angryBirdLarge(129, 130) <= 5; angryBirdLarge(129, 131) <= 5; angryBirdLarge(129, 132) <= 0; angryBirdLarge(129, 133) <= 0; angryBirdLarge(129, 134) <= 0; angryBirdLarge(129, 135) <= 0; angryBirdLarge(129, 136) <= 0; angryBirdLarge(129, 137) <= 0; angryBirdLarge(129, 138) <= 0; angryBirdLarge(129, 139) <= 0; angryBirdLarge(129, 140) <= 0; angryBirdLarge(129, 141) <= 0; angryBirdLarge(129, 142) <= 0; angryBirdLarge(129, 143) <= 0; angryBirdLarge(129, 144) <= 0; angryBirdLarge(129, 145) <= 0; angryBirdLarge(129, 146) <= 0; angryBirdLarge(129, 147) <= 0; angryBirdLarge(129, 148) <= 0; angryBirdLarge(129, 149) <= 0; 
angryBirdLarge(130, 0) <= 0; angryBirdLarge(130, 1) <= 0; angryBirdLarge(130, 2) <= 0; angryBirdLarge(130, 3) <= 0; angryBirdLarge(130, 4) <= 0; angryBirdLarge(130, 5) <= 0; angryBirdLarge(130, 6) <= 0; angryBirdLarge(130, 7) <= 0; angryBirdLarge(130, 8) <= 0; angryBirdLarge(130, 9) <= 0; angryBirdLarge(130, 10) <= 0; angryBirdLarge(130, 11) <= 0; angryBirdLarge(130, 12) <= 0; angryBirdLarge(130, 13) <= 0; angryBirdLarge(130, 14) <= 0; angryBirdLarge(130, 15) <= 0; angryBirdLarge(130, 16) <= 0; angryBirdLarge(130, 17) <= 0; angryBirdLarge(130, 18) <= 0; angryBirdLarge(130, 19) <= 0; angryBirdLarge(130, 20) <= 0; angryBirdLarge(130, 21) <= 0; angryBirdLarge(130, 22) <= 0; angryBirdLarge(130, 23) <= 0; angryBirdLarge(130, 24) <= 0; angryBirdLarge(130, 25) <= 0; angryBirdLarge(130, 26) <= 0; angryBirdLarge(130, 27) <= 0; angryBirdLarge(130, 28) <= 0; angryBirdLarge(130, 29) <= 0; angryBirdLarge(130, 30) <= 0; angryBirdLarge(130, 31) <= 0; angryBirdLarge(130, 32) <= 0; angryBirdLarge(130, 33) <= 0; angryBirdLarge(130, 34) <= 0; angryBirdLarge(130, 35) <= 0; angryBirdLarge(130, 36) <= 0; angryBirdLarge(130, 37) <= 0; angryBirdLarge(130, 38) <= 0; angryBirdLarge(130, 39) <= 0; angryBirdLarge(130, 40) <= 0; angryBirdLarge(130, 41) <= 0; angryBirdLarge(130, 42) <= 0; angryBirdLarge(130, 43) <= 0; angryBirdLarge(130, 44) <= 0; angryBirdLarge(130, 45) <= 0; angryBirdLarge(130, 46) <= 0; angryBirdLarge(130, 47) <= 0; angryBirdLarge(130, 48) <= 5; angryBirdLarge(130, 49) <= 5; angryBirdLarge(130, 50) <= 5; angryBirdLarge(130, 51) <= 5; angryBirdLarge(130, 52) <= 5; angryBirdLarge(130, 53) <= 5; angryBirdLarge(130, 54) <= 5; angryBirdLarge(130, 55) <= 5; angryBirdLarge(130, 56) <= 5; angryBirdLarge(130, 57) <= 5; angryBirdLarge(130, 58) <= 5; angryBirdLarge(130, 59) <= 5; angryBirdLarge(130, 60) <= 2; angryBirdLarge(130, 61) <= 2; angryBirdLarge(130, 62) <= 2; angryBirdLarge(130, 63) <= 2; angryBirdLarge(130, 64) <= 2; angryBirdLarge(130, 65) <= 2; angryBirdLarge(130, 66) <= 2; angryBirdLarge(130, 67) <= 2; angryBirdLarge(130, 68) <= 2; angryBirdLarge(130, 69) <= 2; angryBirdLarge(130, 70) <= 2; angryBirdLarge(130, 71) <= 2; angryBirdLarge(130, 72) <= 2; angryBirdLarge(130, 73) <= 2; angryBirdLarge(130, 74) <= 2; angryBirdLarge(130, 75) <= 2; angryBirdLarge(130, 76) <= 2; angryBirdLarge(130, 77) <= 2; angryBirdLarge(130, 78) <= 2; angryBirdLarge(130, 79) <= 2; angryBirdLarge(130, 80) <= 2; angryBirdLarge(130, 81) <= 2; angryBirdLarge(130, 82) <= 2; angryBirdLarge(130, 83) <= 2; angryBirdLarge(130, 84) <= 2; angryBirdLarge(130, 85) <= 2; angryBirdLarge(130, 86) <= 2; angryBirdLarge(130, 87) <= 2; angryBirdLarge(130, 88) <= 2; angryBirdLarge(130, 89) <= 2; angryBirdLarge(130, 90) <= 2; angryBirdLarge(130, 91) <= 2; angryBirdLarge(130, 92) <= 2; angryBirdLarge(130, 93) <= 2; angryBirdLarge(130, 94) <= 2; angryBirdLarge(130, 95) <= 2; angryBirdLarge(130, 96) <= 2; angryBirdLarge(130, 97) <= 2; angryBirdLarge(130, 98) <= 2; angryBirdLarge(130, 99) <= 2; angryBirdLarge(130, 100) <= 2; angryBirdLarge(130, 101) <= 2; angryBirdLarge(130, 102) <= 2; angryBirdLarge(130, 103) <= 2; angryBirdLarge(130, 104) <= 2; angryBirdLarge(130, 105) <= 2; angryBirdLarge(130, 106) <= 2; angryBirdLarge(130, 107) <= 2; angryBirdLarge(130, 108) <= 2; angryBirdLarge(130, 109) <= 2; angryBirdLarge(130, 110) <= 2; angryBirdLarge(130, 111) <= 2; angryBirdLarge(130, 112) <= 2; angryBirdLarge(130, 113) <= 2; angryBirdLarge(130, 114) <= 2; angryBirdLarge(130, 115) <= 2; angryBirdLarge(130, 116) <= 2; angryBirdLarge(130, 117) <= 2; angryBirdLarge(130, 118) <= 2; angryBirdLarge(130, 119) <= 2; angryBirdLarge(130, 120) <= 2; angryBirdLarge(130, 121) <= 2; angryBirdLarge(130, 122) <= 2; angryBirdLarge(130, 123) <= 2; angryBirdLarge(130, 124) <= 2; angryBirdLarge(130, 125) <= 2; angryBirdLarge(130, 126) <= 5; angryBirdLarge(130, 127) <= 5; angryBirdLarge(130, 128) <= 5; angryBirdLarge(130, 129) <= 5; angryBirdLarge(130, 130) <= 5; angryBirdLarge(130, 131) <= 5; angryBirdLarge(130, 132) <= 0; angryBirdLarge(130, 133) <= 0; angryBirdLarge(130, 134) <= 0; angryBirdLarge(130, 135) <= 0; angryBirdLarge(130, 136) <= 0; angryBirdLarge(130, 137) <= 0; angryBirdLarge(130, 138) <= 0; angryBirdLarge(130, 139) <= 0; angryBirdLarge(130, 140) <= 0; angryBirdLarge(130, 141) <= 0; angryBirdLarge(130, 142) <= 0; angryBirdLarge(130, 143) <= 0; angryBirdLarge(130, 144) <= 0; angryBirdLarge(130, 145) <= 0; angryBirdLarge(130, 146) <= 0; angryBirdLarge(130, 147) <= 0; angryBirdLarge(130, 148) <= 0; angryBirdLarge(130, 149) <= 0; 
angryBirdLarge(131, 0) <= 0; angryBirdLarge(131, 1) <= 0; angryBirdLarge(131, 2) <= 0; angryBirdLarge(131, 3) <= 0; angryBirdLarge(131, 4) <= 0; angryBirdLarge(131, 5) <= 0; angryBirdLarge(131, 6) <= 0; angryBirdLarge(131, 7) <= 0; angryBirdLarge(131, 8) <= 0; angryBirdLarge(131, 9) <= 0; angryBirdLarge(131, 10) <= 0; angryBirdLarge(131, 11) <= 0; angryBirdLarge(131, 12) <= 0; angryBirdLarge(131, 13) <= 0; angryBirdLarge(131, 14) <= 0; angryBirdLarge(131, 15) <= 0; angryBirdLarge(131, 16) <= 0; angryBirdLarge(131, 17) <= 0; angryBirdLarge(131, 18) <= 0; angryBirdLarge(131, 19) <= 0; angryBirdLarge(131, 20) <= 0; angryBirdLarge(131, 21) <= 0; angryBirdLarge(131, 22) <= 0; angryBirdLarge(131, 23) <= 0; angryBirdLarge(131, 24) <= 0; angryBirdLarge(131, 25) <= 0; angryBirdLarge(131, 26) <= 0; angryBirdLarge(131, 27) <= 0; angryBirdLarge(131, 28) <= 0; angryBirdLarge(131, 29) <= 0; angryBirdLarge(131, 30) <= 0; angryBirdLarge(131, 31) <= 0; angryBirdLarge(131, 32) <= 0; angryBirdLarge(131, 33) <= 0; angryBirdLarge(131, 34) <= 0; angryBirdLarge(131, 35) <= 0; angryBirdLarge(131, 36) <= 0; angryBirdLarge(131, 37) <= 0; angryBirdLarge(131, 38) <= 0; angryBirdLarge(131, 39) <= 0; angryBirdLarge(131, 40) <= 0; angryBirdLarge(131, 41) <= 0; angryBirdLarge(131, 42) <= 0; angryBirdLarge(131, 43) <= 0; angryBirdLarge(131, 44) <= 0; angryBirdLarge(131, 45) <= 0; angryBirdLarge(131, 46) <= 0; angryBirdLarge(131, 47) <= 0; angryBirdLarge(131, 48) <= 5; angryBirdLarge(131, 49) <= 5; angryBirdLarge(131, 50) <= 5; angryBirdLarge(131, 51) <= 5; angryBirdLarge(131, 52) <= 5; angryBirdLarge(131, 53) <= 5; angryBirdLarge(131, 54) <= 5; angryBirdLarge(131, 55) <= 5; angryBirdLarge(131, 56) <= 5; angryBirdLarge(131, 57) <= 5; angryBirdLarge(131, 58) <= 5; angryBirdLarge(131, 59) <= 5; angryBirdLarge(131, 60) <= 2; angryBirdLarge(131, 61) <= 2; angryBirdLarge(131, 62) <= 2; angryBirdLarge(131, 63) <= 2; angryBirdLarge(131, 64) <= 2; angryBirdLarge(131, 65) <= 2; angryBirdLarge(131, 66) <= 2; angryBirdLarge(131, 67) <= 2; angryBirdLarge(131, 68) <= 2; angryBirdLarge(131, 69) <= 2; angryBirdLarge(131, 70) <= 2; angryBirdLarge(131, 71) <= 2; angryBirdLarge(131, 72) <= 2; angryBirdLarge(131, 73) <= 2; angryBirdLarge(131, 74) <= 2; angryBirdLarge(131, 75) <= 2; angryBirdLarge(131, 76) <= 2; angryBirdLarge(131, 77) <= 2; angryBirdLarge(131, 78) <= 2; angryBirdLarge(131, 79) <= 2; angryBirdLarge(131, 80) <= 2; angryBirdLarge(131, 81) <= 2; angryBirdLarge(131, 82) <= 2; angryBirdLarge(131, 83) <= 2; angryBirdLarge(131, 84) <= 2; angryBirdLarge(131, 85) <= 2; angryBirdLarge(131, 86) <= 2; angryBirdLarge(131, 87) <= 2; angryBirdLarge(131, 88) <= 2; angryBirdLarge(131, 89) <= 2; angryBirdLarge(131, 90) <= 2; angryBirdLarge(131, 91) <= 2; angryBirdLarge(131, 92) <= 2; angryBirdLarge(131, 93) <= 2; angryBirdLarge(131, 94) <= 2; angryBirdLarge(131, 95) <= 2; angryBirdLarge(131, 96) <= 2; angryBirdLarge(131, 97) <= 2; angryBirdLarge(131, 98) <= 2; angryBirdLarge(131, 99) <= 2; angryBirdLarge(131, 100) <= 2; angryBirdLarge(131, 101) <= 2; angryBirdLarge(131, 102) <= 2; angryBirdLarge(131, 103) <= 2; angryBirdLarge(131, 104) <= 2; angryBirdLarge(131, 105) <= 2; angryBirdLarge(131, 106) <= 2; angryBirdLarge(131, 107) <= 2; angryBirdLarge(131, 108) <= 2; angryBirdLarge(131, 109) <= 2; angryBirdLarge(131, 110) <= 2; angryBirdLarge(131, 111) <= 2; angryBirdLarge(131, 112) <= 2; angryBirdLarge(131, 113) <= 2; angryBirdLarge(131, 114) <= 2; angryBirdLarge(131, 115) <= 2; angryBirdLarge(131, 116) <= 2; angryBirdLarge(131, 117) <= 2; angryBirdLarge(131, 118) <= 2; angryBirdLarge(131, 119) <= 2; angryBirdLarge(131, 120) <= 2; angryBirdLarge(131, 121) <= 2; angryBirdLarge(131, 122) <= 2; angryBirdLarge(131, 123) <= 2; angryBirdLarge(131, 124) <= 2; angryBirdLarge(131, 125) <= 2; angryBirdLarge(131, 126) <= 5; angryBirdLarge(131, 127) <= 5; angryBirdLarge(131, 128) <= 5; angryBirdLarge(131, 129) <= 5; angryBirdLarge(131, 130) <= 5; angryBirdLarge(131, 131) <= 5; angryBirdLarge(131, 132) <= 0; angryBirdLarge(131, 133) <= 0; angryBirdLarge(131, 134) <= 0; angryBirdLarge(131, 135) <= 0; angryBirdLarge(131, 136) <= 0; angryBirdLarge(131, 137) <= 0; angryBirdLarge(131, 138) <= 0; angryBirdLarge(131, 139) <= 0; angryBirdLarge(131, 140) <= 0; angryBirdLarge(131, 141) <= 0; angryBirdLarge(131, 142) <= 0; angryBirdLarge(131, 143) <= 0; angryBirdLarge(131, 144) <= 0; angryBirdLarge(131, 145) <= 0; angryBirdLarge(131, 146) <= 0; angryBirdLarge(131, 147) <= 0; angryBirdLarge(131, 148) <= 0; angryBirdLarge(131, 149) <= 0; 
angryBirdLarge(132, 0) <= 0; angryBirdLarge(132, 1) <= 0; angryBirdLarge(132, 2) <= 0; angryBirdLarge(132, 3) <= 0; angryBirdLarge(132, 4) <= 0; angryBirdLarge(132, 5) <= 0; angryBirdLarge(132, 6) <= 0; angryBirdLarge(132, 7) <= 0; angryBirdLarge(132, 8) <= 0; angryBirdLarge(132, 9) <= 0; angryBirdLarge(132, 10) <= 0; angryBirdLarge(132, 11) <= 0; angryBirdLarge(132, 12) <= 0; angryBirdLarge(132, 13) <= 0; angryBirdLarge(132, 14) <= 0; angryBirdLarge(132, 15) <= 0; angryBirdLarge(132, 16) <= 0; angryBirdLarge(132, 17) <= 0; angryBirdLarge(132, 18) <= 0; angryBirdLarge(132, 19) <= 0; angryBirdLarge(132, 20) <= 0; angryBirdLarge(132, 21) <= 0; angryBirdLarge(132, 22) <= 0; angryBirdLarge(132, 23) <= 0; angryBirdLarge(132, 24) <= 0; angryBirdLarge(132, 25) <= 0; angryBirdLarge(132, 26) <= 0; angryBirdLarge(132, 27) <= 0; angryBirdLarge(132, 28) <= 0; angryBirdLarge(132, 29) <= 0; angryBirdLarge(132, 30) <= 0; angryBirdLarge(132, 31) <= 0; angryBirdLarge(132, 32) <= 0; angryBirdLarge(132, 33) <= 0; angryBirdLarge(132, 34) <= 0; angryBirdLarge(132, 35) <= 0; angryBirdLarge(132, 36) <= 0; angryBirdLarge(132, 37) <= 0; angryBirdLarge(132, 38) <= 0; angryBirdLarge(132, 39) <= 0; angryBirdLarge(132, 40) <= 0; angryBirdLarge(132, 41) <= 0; angryBirdLarge(132, 42) <= 0; angryBirdLarge(132, 43) <= 0; angryBirdLarge(132, 44) <= 0; angryBirdLarge(132, 45) <= 0; angryBirdLarge(132, 46) <= 0; angryBirdLarge(132, 47) <= 0; angryBirdLarge(132, 48) <= 0; angryBirdLarge(132, 49) <= 0; angryBirdLarge(132, 50) <= 0; angryBirdLarge(132, 51) <= 0; angryBirdLarge(132, 52) <= 0; angryBirdLarge(132, 53) <= 0; angryBirdLarge(132, 54) <= 0; angryBirdLarge(132, 55) <= 0; angryBirdLarge(132, 56) <= 0; angryBirdLarge(132, 57) <= 0; angryBirdLarge(132, 58) <= 0; angryBirdLarge(132, 59) <= 0; angryBirdLarge(132, 60) <= 5; angryBirdLarge(132, 61) <= 5; angryBirdLarge(132, 62) <= 5; angryBirdLarge(132, 63) <= 5; angryBirdLarge(132, 64) <= 5; angryBirdLarge(132, 65) <= 5; angryBirdLarge(132, 66) <= 5; angryBirdLarge(132, 67) <= 5; angryBirdLarge(132, 68) <= 5; angryBirdLarge(132, 69) <= 5; angryBirdLarge(132, 70) <= 5; angryBirdLarge(132, 71) <= 5; angryBirdLarge(132, 72) <= 5; angryBirdLarge(132, 73) <= 5; angryBirdLarge(132, 74) <= 5; angryBirdLarge(132, 75) <= 5; angryBirdLarge(132, 76) <= 5; angryBirdLarge(132, 77) <= 5; angryBirdLarge(132, 78) <= 5; angryBirdLarge(132, 79) <= 5; angryBirdLarge(132, 80) <= 5; angryBirdLarge(132, 81) <= 5; angryBirdLarge(132, 82) <= 5; angryBirdLarge(132, 83) <= 5; angryBirdLarge(132, 84) <= 5; angryBirdLarge(132, 85) <= 5; angryBirdLarge(132, 86) <= 5; angryBirdLarge(132, 87) <= 5; angryBirdLarge(132, 88) <= 5; angryBirdLarge(132, 89) <= 5; angryBirdLarge(132, 90) <= 5; angryBirdLarge(132, 91) <= 5; angryBirdLarge(132, 92) <= 5; angryBirdLarge(132, 93) <= 5; angryBirdLarge(132, 94) <= 5; angryBirdLarge(132, 95) <= 5; angryBirdLarge(132, 96) <= 5; angryBirdLarge(132, 97) <= 5; angryBirdLarge(132, 98) <= 5; angryBirdLarge(132, 99) <= 5; angryBirdLarge(132, 100) <= 5; angryBirdLarge(132, 101) <= 5; angryBirdLarge(132, 102) <= 5; angryBirdLarge(132, 103) <= 5; angryBirdLarge(132, 104) <= 5; angryBirdLarge(132, 105) <= 5; angryBirdLarge(132, 106) <= 5; angryBirdLarge(132, 107) <= 5; angryBirdLarge(132, 108) <= 5; angryBirdLarge(132, 109) <= 5; angryBirdLarge(132, 110) <= 5; angryBirdLarge(132, 111) <= 5; angryBirdLarge(132, 112) <= 5; angryBirdLarge(132, 113) <= 5; angryBirdLarge(132, 114) <= 5; angryBirdLarge(132, 115) <= 5; angryBirdLarge(132, 116) <= 5; angryBirdLarge(132, 117) <= 5; angryBirdLarge(132, 118) <= 5; angryBirdLarge(132, 119) <= 5; angryBirdLarge(132, 120) <= 5; angryBirdLarge(132, 121) <= 5; angryBirdLarge(132, 122) <= 5; angryBirdLarge(132, 123) <= 5; angryBirdLarge(132, 124) <= 5; angryBirdLarge(132, 125) <= 5; angryBirdLarge(132, 126) <= 0; angryBirdLarge(132, 127) <= 0; angryBirdLarge(132, 128) <= 0; angryBirdLarge(132, 129) <= 0; angryBirdLarge(132, 130) <= 0; angryBirdLarge(132, 131) <= 0; angryBirdLarge(132, 132) <= 0; angryBirdLarge(132, 133) <= 0; angryBirdLarge(132, 134) <= 0; angryBirdLarge(132, 135) <= 0; angryBirdLarge(132, 136) <= 0; angryBirdLarge(132, 137) <= 0; angryBirdLarge(132, 138) <= 0; angryBirdLarge(132, 139) <= 0; angryBirdLarge(132, 140) <= 0; angryBirdLarge(132, 141) <= 0; angryBirdLarge(132, 142) <= 0; angryBirdLarge(132, 143) <= 0; angryBirdLarge(132, 144) <= 0; angryBirdLarge(132, 145) <= 0; angryBirdLarge(132, 146) <= 0; angryBirdLarge(132, 147) <= 0; angryBirdLarge(132, 148) <= 0; angryBirdLarge(132, 149) <= 0; 
angryBirdLarge(133, 0) <= 0; angryBirdLarge(133, 1) <= 0; angryBirdLarge(133, 2) <= 0; angryBirdLarge(133, 3) <= 0; angryBirdLarge(133, 4) <= 0; angryBirdLarge(133, 5) <= 0; angryBirdLarge(133, 6) <= 0; angryBirdLarge(133, 7) <= 0; angryBirdLarge(133, 8) <= 0; angryBirdLarge(133, 9) <= 0; angryBirdLarge(133, 10) <= 0; angryBirdLarge(133, 11) <= 0; angryBirdLarge(133, 12) <= 0; angryBirdLarge(133, 13) <= 0; angryBirdLarge(133, 14) <= 0; angryBirdLarge(133, 15) <= 0; angryBirdLarge(133, 16) <= 0; angryBirdLarge(133, 17) <= 0; angryBirdLarge(133, 18) <= 0; angryBirdLarge(133, 19) <= 0; angryBirdLarge(133, 20) <= 0; angryBirdLarge(133, 21) <= 0; angryBirdLarge(133, 22) <= 0; angryBirdLarge(133, 23) <= 0; angryBirdLarge(133, 24) <= 0; angryBirdLarge(133, 25) <= 0; angryBirdLarge(133, 26) <= 0; angryBirdLarge(133, 27) <= 0; angryBirdLarge(133, 28) <= 0; angryBirdLarge(133, 29) <= 0; angryBirdLarge(133, 30) <= 0; angryBirdLarge(133, 31) <= 0; angryBirdLarge(133, 32) <= 0; angryBirdLarge(133, 33) <= 0; angryBirdLarge(133, 34) <= 0; angryBirdLarge(133, 35) <= 0; angryBirdLarge(133, 36) <= 0; angryBirdLarge(133, 37) <= 0; angryBirdLarge(133, 38) <= 0; angryBirdLarge(133, 39) <= 0; angryBirdLarge(133, 40) <= 0; angryBirdLarge(133, 41) <= 0; angryBirdLarge(133, 42) <= 0; angryBirdLarge(133, 43) <= 0; angryBirdLarge(133, 44) <= 0; angryBirdLarge(133, 45) <= 0; angryBirdLarge(133, 46) <= 0; angryBirdLarge(133, 47) <= 0; angryBirdLarge(133, 48) <= 0; angryBirdLarge(133, 49) <= 0; angryBirdLarge(133, 50) <= 0; angryBirdLarge(133, 51) <= 0; angryBirdLarge(133, 52) <= 0; angryBirdLarge(133, 53) <= 0; angryBirdLarge(133, 54) <= 0; angryBirdLarge(133, 55) <= 0; angryBirdLarge(133, 56) <= 0; angryBirdLarge(133, 57) <= 0; angryBirdLarge(133, 58) <= 0; angryBirdLarge(133, 59) <= 0; angryBirdLarge(133, 60) <= 5; angryBirdLarge(133, 61) <= 5; angryBirdLarge(133, 62) <= 5; angryBirdLarge(133, 63) <= 5; angryBirdLarge(133, 64) <= 5; angryBirdLarge(133, 65) <= 5; angryBirdLarge(133, 66) <= 5; angryBirdLarge(133, 67) <= 5; angryBirdLarge(133, 68) <= 5; angryBirdLarge(133, 69) <= 5; angryBirdLarge(133, 70) <= 5; angryBirdLarge(133, 71) <= 5; angryBirdLarge(133, 72) <= 5; angryBirdLarge(133, 73) <= 5; angryBirdLarge(133, 74) <= 5; angryBirdLarge(133, 75) <= 5; angryBirdLarge(133, 76) <= 5; angryBirdLarge(133, 77) <= 5; angryBirdLarge(133, 78) <= 5; angryBirdLarge(133, 79) <= 5; angryBirdLarge(133, 80) <= 5; angryBirdLarge(133, 81) <= 5; angryBirdLarge(133, 82) <= 5; angryBirdLarge(133, 83) <= 5; angryBirdLarge(133, 84) <= 5; angryBirdLarge(133, 85) <= 5; angryBirdLarge(133, 86) <= 5; angryBirdLarge(133, 87) <= 5; angryBirdLarge(133, 88) <= 5; angryBirdLarge(133, 89) <= 5; angryBirdLarge(133, 90) <= 5; angryBirdLarge(133, 91) <= 5; angryBirdLarge(133, 92) <= 5; angryBirdLarge(133, 93) <= 5; angryBirdLarge(133, 94) <= 5; angryBirdLarge(133, 95) <= 5; angryBirdLarge(133, 96) <= 5; angryBirdLarge(133, 97) <= 5; angryBirdLarge(133, 98) <= 5; angryBirdLarge(133, 99) <= 5; angryBirdLarge(133, 100) <= 5; angryBirdLarge(133, 101) <= 5; angryBirdLarge(133, 102) <= 5; angryBirdLarge(133, 103) <= 5; angryBirdLarge(133, 104) <= 5; angryBirdLarge(133, 105) <= 5; angryBirdLarge(133, 106) <= 5; angryBirdLarge(133, 107) <= 5; angryBirdLarge(133, 108) <= 5; angryBirdLarge(133, 109) <= 5; angryBirdLarge(133, 110) <= 5; angryBirdLarge(133, 111) <= 5; angryBirdLarge(133, 112) <= 5; angryBirdLarge(133, 113) <= 5; angryBirdLarge(133, 114) <= 5; angryBirdLarge(133, 115) <= 5; angryBirdLarge(133, 116) <= 5; angryBirdLarge(133, 117) <= 5; angryBirdLarge(133, 118) <= 5; angryBirdLarge(133, 119) <= 5; angryBirdLarge(133, 120) <= 5; angryBirdLarge(133, 121) <= 5; angryBirdLarge(133, 122) <= 5; angryBirdLarge(133, 123) <= 5; angryBirdLarge(133, 124) <= 5; angryBirdLarge(133, 125) <= 5; angryBirdLarge(133, 126) <= 0; angryBirdLarge(133, 127) <= 0; angryBirdLarge(133, 128) <= 0; angryBirdLarge(133, 129) <= 0; angryBirdLarge(133, 130) <= 0; angryBirdLarge(133, 131) <= 0; angryBirdLarge(133, 132) <= 0; angryBirdLarge(133, 133) <= 0; angryBirdLarge(133, 134) <= 0; angryBirdLarge(133, 135) <= 0; angryBirdLarge(133, 136) <= 0; angryBirdLarge(133, 137) <= 0; angryBirdLarge(133, 138) <= 0; angryBirdLarge(133, 139) <= 0; angryBirdLarge(133, 140) <= 0; angryBirdLarge(133, 141) <= 0; angryBirdLarge(133, 142) <= 0; angryBirdLarge(133, 143) <= 0; angryBirdLarge(133, 144) <= 0; angryBirdLarge(133, 145) <= 0; angryBirdLarge(133, 146) <= 0; angryBirdLarge(133, 147) <= 0; angryBirdLarge(133, 148) <= 0; angryBirdLarge(133, 149) <= 0; 
angryBirdLarge(134, 0) <= 0; angryBirdLarge(134, 1) <= 0; angryBirdLarge(134, 2) <= 0; angryBirdLarge(134, 3) <= 0; angryBirdLarge(134, 4) <= 0; angryBirdLarge(134, 5) <= 0; angryBirdLarge(134, 6) <= 0; angryBirdLarge(134, 7) <= 0; angryBirdLarge(134, 8) <= 0; angryBirdLarge(134, 9) <= 0; angryBirdLarge(134, 10) <= 0; angryBirdLarge(134, 11) <= 0; angryBirdLarge(134, 12) <= 0; angryBirdLarge(134, 13) <= 0; angryBirdLarge(134, 14) <= 0; angryBirdLarge(134, 15) <= 0; angryBirdLarge(134, 16) <= 0; angryBirdLarge(134, 17) <= 0; angryBirdLarge(134, 18) <= 0; angryBirdLarge(134, 19) <= 0; angryBirdLarge(134, 20) <= 0; angryBirdLarge(134, 21) <= 0; angryBirdLarge(134, 22) <= 0; angryBirdLarge(134, 23) <= 0; angryBirdLarge(134, 24) <= 0; angryBirdLarge(134, 25) <= 0; angryBirdLarge(134, 26) <= 0; angryBirdLarge(134, 27) <= 0; angryBirdLarge(134, 28) <= 0; angryBirdLarge(134, 29) <= 0; angryBirdLarge(134, 30) <= 0; angryBirdLarge(134, 31) <= 0; angryBirdLarge(134, 32) <= 0; angryBirdLarge(134, 33) <= 0; angryBirdLarge(134, 34) <= 0; angryBirdLarge(134, 35) <= 0; angryBirdLarge(134, 36) <= 0; angryBirdLarge(134, 37) <= 0; angryBirdLarge(134, 38) <= 0; angryBirdLarge(134, 39) <= 0; angryBirdLarge(134, 40) <= 0; angryBirdLarge(134, 41) <= 0; angryBirdLarge(134, 42) <= 0; angryBirdLarge(134, 43) <= 0; angryBirdLarge(134, 44) <= 0; angryBirdLarge(134, 45) <= 0; angryBirdLarge(134, 46) <= 0; angryBirdLarge(134, 47) <= 0; angryBirdLarge(134, 48) <= 0; angryBirdLarge(134, 49) <= 0; angryBirdLarge(134, 50) <= 0; angryBirdLarge(134, 51) <= 0; angryBirdLarge(134, 52) <= 0; angryBirdLarge(134, 53) <= 0; angryBirdLarge(134, 54) <= 0; angryBirdLarge(134, 55) <= 0; angryBirdLarge(134, 56) <= 0; angryBirdLarge(134, 57) <= 0; angryBirdLarge(134, 58) <= 0; angryBirdLarge(134, 59) <= 0; angryBirdLarge(134, 60) <= 5; angryBirdLarge(134, 61) <= 5; angryBirdLarge(134, 62) <= 5; angryBirdLarge(134, 63) <= 5; angryBirdLarge(134, 64) <= 5; angryBirdLarge(134, 65) <= 5; angryBirdLarge(134, 66) <= 5; angryBirdLarge(134, 67) <= 5; angryBirdLarge(134, 68) <= 5; angryBirdLarge(134, 69) <= 5; angryBirdLarge(134, 70) <= 5; angryBirdLarge(134, 71) <= 5; angryBirdLarge(134, 72) <= 5; angryBirdLarge(134, 73) <= 5; angryBirdLarge(134, 74) <= 5; angryBirdLarge(134, 75) <= 5; angryBirdLarge(134, 76) <= 5; angryBirdLarge(134, 77) <= 5; angryBirdLarge(134, 78) <= 5; angryBirdLarge(134, 79) <= 5; angryBirdLarge(134, 80) <= 5; angryBirdLarge(134, 81) <= 5; angryBirdLarge(134, 82) <= 5; angryBirdLarge(134, 83) <= 5; angryBirdLarge(134, 84) <= 5; angryBirdLarge(134, 85) <= 5; angryBirdLarge(134, 86) <= 5; angryBirdLarge(134, 87) <= 5; angryBirdLarge(134, 88) <= 5; angryBirdLarge(134, 89) <= 5; angryBirdLarge(134, 90) <= 5; angryBirdLarge(134, 91) <= 5; angryBirdLarge(134, 92) <= 5; angryBirdLarge(134, 93) <= 5; angryBirdLarge(134, 94) <= 5; angryBirdLarge(134, 95) <= 5; angryBirdLarge(134, 96) <= 5; angryBirdLarge(134, 97) <= 5; angryBirdLarge(134, 98) <= 5; angryBirdLarge(134, 99) <= 5; angryBirdLarge(134, 100) <= 5; angryBirdLarge(134, 101) <= 5; angryBirdLarge(134, 102) <= 5; angryBirdLarge(134, 103) <= 5; angryBirdLarge(134, 104) <= 5; angryBirdLarge(134, 105) <= 5; angryBirdLarge(134, 106) <= 5; angryBirdLarge(134, 107) <= 5; angryBirdLarge(134, 108) <= 5; angryBirdLarge(134, 109) <= 5; angryBirdLarge(134, 110) <= 5; angryBirdLarge(134, 111) <= 5; angryBirdLarge(134, 112) <= 5; angryBirdLarge(134, 113) <= 5; angryBirdLarge(134, 114) <= 5; angryBirdLarge(134, 115) <= 5; angryBirdLarge(134, 116) <= 5; angryBirdLarge(134, 117) <= 5; angryBirdLarge(134, 118) <= 5; angryBirdLarge(134, 119) <= 5; angryBirdLarge(134, 120) <= 5; angryBirdLarge(134, 121) <= 5; angryBirdLarge(134, 122) <= 5; angryBirdLarge(134, 123) <= 5; angryBirdLarge(134, 124) <= 5; angryBirdLarge(134, 125) <= 5; angryBirdLarge(134, 126) <= 0; angryBirdLarge(134, 127) <= 0; angryBirdLarge(134, 128) <= 0; angryBirdLarge(134, 129) <= 0; angryBirdLarge(134, 130) <= 0; angryBirdLarge(134, 131) <= 0; angryBirdLarge(134, 132) <= 0; angryBirdLarge(134, 133) <= 0; angryBirdLarge(134, 134) <= 0; angryBirdLarge(134, 135) <= 0; angryBirdLarge(134, 136) <= 0; angryBirdLarge(134, 137) <= 0; angryBirdLarge(134, 138) <= 0; angryBirdLarge(134, 139) <= 0; angryBirdLarge(134, 140) <= 0; angryBirdLarge(134, 141) <= 0; angryBirdLarge(134, 142) <= 0; angryBirdLarge(134, 143) <= 0; angryBirdLarge(134, 144) <= 0; angryBirdLarge(134, 145) <= 0; angryBirdLarge(134, 146) <= 0; angryBirdLarge(134, 147) <= 0; angryBirdLarge(134, 148) <= 0; angryBirdLarge(134, 149) <= 0; 
angryBirdLarge(135, 0) <= 0; angryBirdLarge(135, 1) <= 0; angryBirdLarge(135, 2) <= 0; angryBirdLarge(135, 3) <= 0; angryBirdLarge(135, 4) <= 0; angryBirdLarge(135, 5) <= 0; angryBirdLarge(135, 6) <= 0; angryBirdLarge(135, 7) <= 0; angryBirdLarge(135, 8) <= 0; angryBirdLarge(135, 9) <= 0; angryBirdLarge(135, 10) <= 0; angryBirdLarge(135, 11) <= 0; angryBirdLarge(135, 12) <= 0; angryBirdLarge(135, 13) <= 0; angryBirdLarge(135, 14) <= 0; angryBirdLarge(135, 15) <= 0; angryBirdLarge(135, 16) <= 0; angryBirdLarge(135, 17) <= 0; angryBirdLarge(135, 18) <= 0; angryBirdLarge(135, 19) <= 0; angryBirdLarge(135, 20) <= 0; angryBirdLarge(135, 21) <= 0; angryBirdLarge(135, 22) <= 0; angryBirdLarge(135, 23) <= 0; angryBirdLarge(135, 24) <= 0; angryBirdLarge(135, 25) <= 0; angryBirdLarge(135, 26) <= 0; angryBirdLarge(135, 27) <= 0; angryBirdLarge(135, 28) <= 0; angryBirdLarge(135, 29) <= 0; angryBirdLarge(135, 30) <= 0; angryBirdLarge(135, 31) <= 0; angryBirdLarge(135, 32) <= 0; angryBirdLarge(135, 33) <= 0; angryBirdLarge(135, 34) <= 0; angryBirdLarge(135, 35) <= 0; angryBirdLarge(135, 36) <= 0; angryBirdLarge(135, 37) <= 0; angryBirdLarge(135, 38) <= 0; angryBirdLarge(135, 39) <= 0; angryBirdLarge(135, 40) <= 0; angryBirdLarge(135, 41) <= 0; angryBirdLarge(135, 42) <= 0; angryBirdLarge(135, 43) <= 0; angryBirdLarge(135, 44) <= 0; angryBirdLarge(135, 45) <= 0; angryBirdLarge(135, 46) <= 0; angryBirdLarge(135, 47) <= 0; angryBirdLarge(135, 48) <= 0; angryBirdLarge(135, 49) <= 0; angryBirdLarge(135, 50) <= 0; angryBirdLarge(135, 51) <= 0; angryBirdLarge(135, 52) <= 0; angryBirdLarge(135, 53) <= 0; angryBirdLarge(135, 54) <= 0; angryBirdLarge(135, 55) <= 0; angryBirdLarge(135, 56) <= 0; angryBirdLarge(135, 57) <= 0; angryBirdLarge(135, 58) <= 0; angryBirdLarge(135, 59) <= 0; angryBirdLarge(135, 60) <= 5; angryBirdLarge(135, 61) <= 5; angryBirdLarge(135, 62) <= 5; angryBirdLarge(135, 63) <= 5; angryBirdLarge(135, 64) <= 5; angryBirdLarge(135, 65) <= 5; angryBirdLarge(135, 66) <= 5; angryBirdLarge(135, 67) <= 5; angryBirdLarge(135, 68) <= 5; angryBirdLarge(135, 69) <= 5; angryBirdLarge(135, 70) <= 5; angryBirdLarge(135, 71) <= 5; angryBirdLarge(135, 72) <= 5; angryBirdLarge(135, 73) <= 5; angryBirdLarge(135, 74) <= 5; angryBirdLarge(135, 75) <= 5; angryBirdLarge(135, 76) <= 5; angryBirdLarge(135, 77) <= 5; angryBirdLarge(135, 78) <= 5; angryBirdLarge(135, 79) <= 5; angryBirdLarge(135, 80) <= 5; angryBirdLarge(135, 81) <= 5; angryBirdLarge(135, 82) <= 5; angryBirdLarge(135, 83) <= 5; angryBirdLarge(135, 84) <= 5; angryBirdLarge(135, 85) <= 5; angryBirdLarge(135, 86) <= 5; angryBirdLarge(135, 87) <= 5; angryBirdLarge(135, 88) <= 5; angryBirdLarge(135, 89) <= 5; angryBirdLarge(135, 90) <= 5; angryBirdLarge(135, 91) <= 5; angryBirdLarge(135, 92) <= 5; angryBirdLarge(135, 93) <= 5; angryBirdLarge(135, 94) <= 5; angryBirdLarge(135, 95) <= 5; angryBirdLarge(135, 96) <= 5; angryBirdLarge(135, 97) <= 5; angryBirdLarge(135, 98) <= 5; angryBirdLarge(135, 99) <= 5; angryBirdLarge(135, 100) <= 5; angryBirdLarge(135, 101) <= 5; angryBirdLarge(135, 102) <= 5; angryBirdLarge(135, 103) <= 5; angryBirdLarge(135, 104) <= 5; angryBirdLarge(135, 105) <= 5; angryBirdLarge(135, 106) <= 5; angryBirdLarge(135, 107) <= 5; angryBirdLarge(135, 108) <= 5; angryBirdLarge(135, 109) <= 5; angryBirdLarge(135, 110) <= 5; angryBirdLarge(135, 111) <= 5; angryBirdLarge(135, 112) <= 5; angryBirdLarge(135, 113) <= 5; angryBirdLarge(135, 114) <= 5; angryBirdLarge(135, 115) <= 5; angryBirdLarge(135, 116) <= 5; angryBirdLarge(135, 117) <= 5; angryBirdLarge(135, 118) <= 5; angryBirdLarge(135, 119) <= 5; angryBirdLarge(135, 120) <= 5; angryBirdLarge(135, 121) <= 5; angryBirdLarge(135, 122) <= 5; angryBirdLarge(135, 123) <= 5; angryBirdLarge(135, 124) <= 5; angryBirdLarge(135, 125) <= 5; angryBirdLarge(135, 126) <= 0; angryBirdLarge(135, 127) <= 0; angryBirdLarge(135, 128) <= 0; angryBirdLarge(135, 129) <= 0; angryBirdLarge(135, 130) <= 0; angryBirdLarge(135, 131) <= 0; angryBirdLarge(135, 132) <= 0; angryBirdLarge(135, 133) <= 0; angryBirdLarge(135, 134) <= 0; angryBirdLarge(135, 135) <= 0; angryBirdLarge(135, 136) <= 0; angryBirdLarge(135, 137) <= 0; angryBirdLarge(135, 138) <= 0; angryBirdLarge(135, 139) <= 0; angryBirdLarge(135, 140) <= 0; angryBirdLarge(135, 141) <= 0; angryBirdLarge(135, 142) <= 0; angryBirdLarge(135, 143) <= 0; angryBirdLarge(135, 144) <= 0; angryBirdLarge(135, 145) <= 0; angryBirdLarge(135, 146) <= 0; angryBirdLarge(135, 147) <= 0; angryBirdLarge(135, 148) <= 0; angryBirdLarge(135, 149) <= 0; 
angryBirdLarge(136, 0) <= 0; angryBirdLarge(136, 1) <= 0; angryBirdLarge(136, 2) <= 0; angryBirdLarge(136, 3) <= 0; angryBirdLarge(136, 4) <= 0; angryBirdLarge(136, 5) <= 0; angryBirdLarge(136, 6) <= 0; angryBirdLarge(136, 7) <= 0; angryBirdLarge(136, 8) <= 0; angryBirdLarge(136, 9) <= 0; angryBirdLarge(136, 10) <= 0; angryBirdLarge(136, 11) <= 0; angryBirdLarge(136, 12) <= 0; angryBirdLarge(136, 13) <= 0; angryBirdLarge(136, 14) <= 0; angryBirdLarge(136, 15) <= 0; angryBirdLarge(136, 16) <= 0; angryBirdLarge(136, 17) <= 0; angryBirdLarge(136, 18) <= 0; angryBirdLarge(136, 19) <= 0; angryBirdLarge(136, 20) <= 0; angryBirdLarge(136, 21) <= 0; angryBirdLarge(136, 22) <= 0; angryBirdLarge(136, 23) <= 0; angryBirdLarge(136, 24) <= 0; angryBirdLarge(136, 25) <= 0; angryBirdLarge(136, 26) <= 0; angryBirdLarge(136, 27) <= 0; angryBirdLarge(136, 28) <= 0; angryBirdLarge(136, 29) <= 0; angryBirdLarge(136, 30) <= 0; angryBirdLarge(136, 31) <= 0; angryBirdLarge(136, 32) <= 0; angryBirdLarge(136, 33) <= 0; angryBirdLarge(136, 34) <= 0; angryBirdLarge(136, 35) <= 0; angryBirdLarge(136, 36) <= 0; angryBirdLarge(136, 37) <= 0; angryBirdLarge(136, 38) <= 0; angryBirdLarge(136, 39) <= 0; angryBirdLarge(136, 40) <= 0; angryBirdLarge(136, 41) <= 0; angryBirdLarge(136, 42) <= 0; angryBirdLarge(136, 43) <= 0; angryBirdLarge(136, 44) <= 0; angryBirdLarge(136, 45) <= 0; angryBirdLarge(136, 46) <= 0; angryBirdLarge(136, 47) <= 0; angryBirdLarge(136, 48) <= 0; angryBirdLarge(136, 49) <= 0; angryBirdLarge(136, 50) <= 0; angryBirdLarge(136, 51) <= 0; angryBirdLarge(136, 52) <= 0; angryBirdLarge(136, 53) <= 0; angryBirdLarge(136, 54) <= 0; angryBirdLarge(136, 55) <= 0; angryBirdLarge(136, 56) <= 0; angryBirdLarge(136, 57) <= 0; angryBirdLarge(136, 58) <= 0; angryBirdLarge(136, 59) <= 0; angryBirdLarge(136, 60) <= 5; angryBirdLarge(136, 61) <= 5; angryBirdLarge(136, 62) <= 5; angryBirdLarge(136, 63) <= 5; angryBirdLarge(136, 64) <= 5; angryBirdLarge(136, 65) <= 5; angryBirdLarge(136, 66) <= 5; angryBirdLarge(136, 67) <= 5; angryBirdLarge(136, 68) <= 5; angryBirdLarge(136, 69) <= 5; angryBirdLarge(136, 70) <= 5; angryBirdLarge(136, 71) <= 5; angryBirdLarge(136, 72) <= 5; angryBirdLarge(136, 73) <= 5; angryBirdLarge(136, 74) <= 5; angryBirdLarge(136, 75) <= 5; angryBirdLarge(136, 76) <= 5; angryBirdLarge(136, 77) <= 5; angryBirdLarge(136, 78) <= 5; angryBirdLarge(136, 79) <= 5; angryBirdLarge(136, 80) <= 5; angryBirdLarge(136, 81) <= 5; angryBirdLarge(136, 82) <= 5; angryBirdLarge(136, 83) <= 5; angryBirdLarge(136, 84) <= 5; angryBirdLarge(136, 85) <= 5; angryBirdLarge(136, 86) <= 5; angryBirdLarge(136, 87) <= 5; angryBirdLarge(136, 88) <= 5; angryBirdLarge(136, 89) <= 5; angryBirdLarge(136, 90) <= 5; angryBirdLarge(136, 91) <= 5; angryBirdLarge(136, 92) <= 5; angryBirdLarge(136, 93) <= 5; angryBirdLarge(136, 94) <= 5; angryBirdLarge(136, 95) <= 5; angryBirdLarge(136, 96) <= 5; angryBirdLarge(136, 97) <= 5; angryBirdLarge(136, 98) <= 5; angryBirdLarge(136, 99) <= 5; angryBirdLarge(136, 100) <= 5; angryBirdLarge(136, 101) <= 5; angryBirdLarge(136, 102) <= 5; angryBirdLarge(136, 103) <= 5; angryBirdLarge(136, 104) <= 5; angryBirdLarge(136, 105) <= 5; angryBirdLarge(136, 106) <= 5; angryBirdLarge(136, 107) <= 5; angryBirdLarge(136, 108) <= 5; angryBirdLarge(136, 109) <= 5; angryBirdLarge(136, 110) <= 5; angryBirdLarge(136, 111) <= 5; angryBirdLarge(136, 112) <= 5; angryBirdLarge(136, 113) <= 5; angryBirdLarge(136, 114) <= 5; angryBirdLarge(136, 115) <= 5; angryBirdLarge(136, 116) <= 5; angryBirdLarge(136, 117) <= 5; angryBirdLarge(136, 118) <= 5; angryBirdLarge(136, 119) <= 5; angryBirdLarge(136, 120) <= 5; angryBirdLarge(136, 121) <= 5; angryBirdLarge(136, 122) <= 5; angryBirdLarge(136, 123) <= 5; angryBirdLarge(136, 124) <= 5; angryBirdLarge(136, 125) <= 5; angryBirdLarge(136, 126) <= 0; angryBirdLarge(136, 127) <= 0; angryBirdLarge(136, 128) <= 0; angryBirdLarge(136, 129) <= 0; angryBirdLarge(136, 130) <= 0; angryBirdLarge(136, 131) <= 0; angryBirdLarge(136, 132) <= 0; angryBirdLarge(136, 133) <= 0; angryBirdLarge(136, 134) <= 0; angryBirdLarge(136, 135) <= 0; angryBirdLarge(136, 136) <= 0; angryBirdLarge(136, 137) <= 0; angryBirdLarge(136, 138) <= 0; angryBirdLarge(136, 139) <= 0; angryBirdLarge(136, 140) <= 0; angryBirdLarge(136, 141) <= 0; angryBirdLarge(136, 142) <= 0; angryBirdLarge(136, 143) <= 0; angryBirdLarge(136, 144) <= 0; angryBirdLarge(136, 145) <= 0; angryBirdLarge(136, 146) <= 0; angryBirdLarge(136, 147) <= 0; angryBirdLarge(136, 148) <= 0; angryBirdLarge(136, 149) <= 0; 
angryBirdLarge(137, 0) <= 0; angryBirdLarge(137, 1) <= 0; angryBirdLarge(137, 2) <= 0; angryBirdLarge(137, 3) <= 0; angryBirdLarge(137, 4) <= 0; angryBirdLarge(137, 5) <= 0; angryBirdLarge(137, 6) <= 0; angryBirdLarge(137, 7) <= 0; angryBirdLarge(137, 8) <= 0; angryBirdLarge(137, 9) <= 0; angryBirdLarge(137, 10) <= 0; angryBirdLarge(137, 11) <= 0; angryBirdLarge(137, 12) <= 0; angryBirdLarge(137, 13) <= 0; angryBirdLarge(137, 14) <= 0; angryBirdLarge(137, 15) <= 0; angryBirdLarge(137, 16) <= 0; angryBirdLarge(137, 17) <= 0; angryBirdLarge(137, 18) <= 0; angryBirdLarge(137, 19) <= 0; angryBirdLarge(137, 20) <= 0; angryBirdLarge(137, 21) <= 0; angryBirdLarge(137, 22) <= 0; angryBirdLarge(137, 23) <= 0; angryBirdLarge(137, 24) <= 0; angryBirdLarge(137, 25) <= 0; angryBirdLarge(137, 26) <= 0; angryBirdLarge(137, 27) <= 0; angryBirdLarge(137, 28) <= 0; angryBirdLarge(137, 29) <= 0; angryBirdLarge(137, 30) <= 0; angryBirdLarge(137, 31) <= 0; angryBirdLarge(137, 32) <= 0; angryBirdLarge(137, 33) <= 0; angryBirdLarge(137, 34) <= 0; angryBirdLarge(137, 35) <= 0; angryBirdLarge(137, 36) <= 0; angryBirdLarge(137, 37) <= 0; angryBirdLarge(137, 38) <= 0; angryBirdLarge(137, 39) <= 0; angryBirdLarge(137, 40) <= 0; angryBirdLarge(137, 41) <= 0; angryBirdLarge(137, 42) <= 0; angryBirdLarge(137, 43) <= 0; angryBirdLarge(137, 44) <= 0; angryBirdLarge(137, 45) <= 0; angryBirdLarge(137, 46) <= 0; angryBirdLarge(137, 47) <= 0; angryBirdLarge(137, 48) <= 0; angryBirdLarge(137, 49) <= 0; angryBirdLarge(137, 50) <= 0; angryBirdLarge(137, 51) <= 0; angryBirdLarge(137, 52) <= 0; angryBirdLarge(137, 53) <= 0; angryBirdLarge(137, 54) <= 0; angryBirdLarge(137, 55) <= 0; angryBirdLarge(137, 56) <= 0; angryBirdLarge(137, 57) <= 0; angryBirdLarge(137, 58) <= 0; angryBirdLarge(137, 59) <= 0; angryBirdLarge(137, 60) <= 5; angryBirdLarge(137, 61) <= 5; angryBirdLarge(137, 62) <= 5; angryBirdLarge(137, 63) <= 5; angryBirdLarge(137, 64) <= 5; angryBirdLarge(137, 65) <= 5; angryBirdLarge(137, 66) <= 5; angryBirdLarge(137, 67) <= 5; angryBirdLarge(137, 68) <= 5; angryBirdLarge(137, 69) <= 5; angryBirdLarge(137, 70) <= 5; angryBirdLarge(137, 71) <= 5; angryBirdLarge(137, 72) <= 5; angryBirdLarge(137, 73) <= 5; angryBirdLarge(137, 74) <= 5; angryBirdLarge(137, 75) <= 5; angryBirdLarge(137, 76) <= 5; angryBirdLarge(137, 77) <= 5; angryBirdLarge(137, 78) <= 5; angryBirdLarge(137, 79) <= 5; angryBirdLarge(137, 80) <= 5; angryBirdLarge(137, 81) <= 5; angryBirdLarge(137, 82) <= 5; angryBirdLarge(137, 83) <= 5; angryBirdLarge(137, 84) <= 5; angryBirdLarge(137, 85) <= 5; angryBirdLarge(137, 86) <= 5; angryBirdLarge(137, 87) <= 5; angryBirdLarge(137, 88) <= 5; angryBirdLarge(137, 89) <= 5; angryBirdLarge(137, 90) <= 5; angryBirdLarge(137, 91) <= 5; angryBirdLarge(137, 92) <= 5; angryBirdLarge(137, 93) <= 5; angryBirdLarge(137, 94) <= 5; angryBirdLarge(137, 95) <= 5; angryBirdLarge(137, 96) <= 5; angryBirdLarge(137, 97) <= 5; angryBirdLarge(137, 98) <= 5; angryBirdLarge(137, 99) <= 5; angryBirdLarge(137, 100) <= 5; angryBirdLarge(137, 101) <= 5; angryBirdLarge(137, 102) <= 5; angryBirdLarge(137, 103) <= 5; angryBirdLarge(137, 104) <= 5; angryBirdLarge(137, 105) <= 5; angryBirdLarge(137, 106) <= 5; angryBirdLarge(137, 107) <= 5; angryBirdLarge(137, 108) <= 5; angryBirdLarge(137, 109) <= 5; angryBirdLarge(137, 110) <= 5; angryBirdLarge(137, 111) <= 5; angryBirdLarge(137, 112) <= 5; angryBirdLarge(137, 113) <= 5; angryBirdLarge(137, 114) <= 5; angryBirdLarge(137, 115) <= 5; angryBirdLarge(137, 116) <= 5; angryBirdLarge(137, 117) <= 5; angryBirdLarge(137, 118) <= 5; angryBirdLarge(137, 119) <= 5; angryBirdLarge(137, 120) <= 5; angryBirdLarge(137, 121) <= 5; angryBirdLarge(137, 122) <= 5; angryBirdLarge(137, 123) <= 5; angryBirdLarge(137, 124) <= 5; angryBirdLarge(137, 125) <= 5; angryBirdLarge(137, 126) <= 0; angryBirdLarge(137, 127) <= 0; angryBirdLarge(137, 128) <= 0; angryBirdLarge(137, 129) <= 0; angryBirdLarge(137, 130) <= 0; angryBirdLarge(137, 131) <= 0; angryBirdLarge(137, 132) <= 0; angryBirdLarge(137, 133) <= 0; angryBirdLarge(137, 134) <= 0; angryBirdLarge(137, 135) <= 0; angryBirdLarge(137, 136) <= 0; angryBirdLarge(137, 137) <= 0; angryBirdLarge(137, 138) <= 0; angryBirdLarge(137, 139) <= 0; angryBirdLarge(137, 140) <= 0; angryBirdLarge(137, 141) <= 0; angryBirdLarge(137, 142) <= 0; angryBirdLarge(137, 143) <= 0; angryBirdLarge(137, 144) <= 0; angryBirdLarge(137, 145) <= 0; angryBirdLarge(137, 146) <= 0; angryBirdLarge(137, 147) <= 0; angryBirdLarge(137, 148) <= 0; angryBirdLarge(137, 149) <= 0; 
angryBirdLarge(138, 0) <= 0; angryBirdLarge(138, 1) <= 0; angryBirdLarge(138, 2) <= 0; angryBirdLarge(138, 3) <= 0; angryBirdLarge(138, 4) <= 0; angryBirdLarge(138, 5) <= 0; angryBirdLarge(138, 6) <= 0; angryBirdLarge(138, 7) <= 0; angryBirdLarge(138, 8) <= 0; angryBirdLarge(138, 9) <= 0; angryBirdLarge(138, 10) <= 0; angryBirdLarge(138, 11) <= 0; angryBirdLarge(138, 12) <= 0; angryBirdLarge(138, 13) <= 0; angryBirdLarge(138, 14) <= 0; angryBirdLarge(138, 15) <= 0; angryBirdLarge(138, 16) <= 0; angryBirdLarge(138, 17) <= 0; angryBirdLarge(138, 18) <= 0; angryBirdLarge(138, 19) <= 0; angryBirdLarge(138, 20) <= 0; angryBirdLarge(138, 21) <= 0; angryBirdLarge(138, 22) <= 0; angryBirdLarge(138, 23) <= 0; angryBirdLarge(138, 24) <= 0; angryBirdLarge(138, 25) <= 0; angryBirdLarge(138, 26) <= 0; angryBirdLarge(138, 27) <= 0; angryBirdLarge(138, 28) <= 0; angryBirdLarge(138, 29) <= 0; angryBirdLarge(138, 30) <= 0; angryBirdLarge(138, 31) <= 0; angryBirdLarge(138, 32) <= 0; angryBirdLarge(138, 33) <= 0; angryBirdLarge(138, 34) <= 0; angryBirdLarge(138, 35) <= 0; angryBirdLarge(138, 36) <= 0; angryBirdLarge(138, 37) <= 0; angryBirdLarge(138, 38) <= 0; angryBirdLarge(138, 39) <= 0; angryBirdLarge(138, 40) <= 0; angryBirdLarge(138, 41) <= 0; angryBirdLarge(138, 42) <= 0; angryBirdLarge(138, 43) <= 0; angryBirdLarge(138, 44) <= 0; angryBirdLarge(138, 45) <= 0; angryBirdLarge(138, 46) <= 0; angryBirdLarge(138, 47) <= 0; angryBirdLarge(138, 48) <= 0; angryBirdLarge(138, 49) <= 0; angryBirdLarge(138, 50) <= 0; angryBirdLarge(138, 51) <= 0; angryBirdLarge(138, 52) <= 0; angryBirdLarge(138, 53) <= 0; angryBirdLarge(138, 54) <= 0; angryBirdLarge(138, 55) <= 0; angryBirdLarge(138, 56) <= 0; angryBirdLarge(138, 57) <= 0; angryBirdLarge(138, 58) <= 0; angryBirdLarge(138, 59) <= 0; angryBirdLarge(138, 60) <= 0; angryBirdLarge(138, 61) <= 0; angryBirdLarge(138, 62) <= 0; angryBirdLarge(138, 63) <= 0; angryBirdLarge(138, 64) <= 0; angryBirdLarge(138, 65) <= 0; angryBirdLarge(138, 66) <= 0; angryBirdLarge(138, 67) <= 0; angryBirdLarge(138, 68) <= 0; angryBirdLarge(138, 69) <= 0; angryBirdLarge(138, 70) <= 0; angryBirdLarge(138, 71) <= 0; angryBirdLarge(138, 72) <= 0; angryBirdLarge(138, 73) <= 0; angryBirdLarge(138, 74) <= 0; angryBirdLarge(138, 75) <= 0; angryBirdLarge(138, 76) <= 0; angryBirdLarge(138, 77) <= 0; angryBirdLarge(138, 78) <= 0; angryBirdLarge(138, 79) <= 0; angryBirdLarge(138, 80) <= 0; angryBirdLarge(138, 81) <= 0; angryBirdLarge(138, 82) <= 0; angryBirdLarge(138, 83) <= 0; angryBirdLarge(138, 84) <= 0; angryBirdLarge(138, 85) <= 0; angryBirdLarge(138, 86) <= 0; angryBirdLarge(138, 87) <= 0; angryBirdLarge(138, 88) <= 0; angryBirdLarge(138, 89) <= 0; angryBirdLarge(138, 90) <= 0; angryBirdLarge(138, 91) <= 0; angryBirdLarge(138, 92) <= 0; angryBirdLarge(138, 93) <= 0; angryBirdLarge(138, 94) <= 0; angryBirdLarge(138, 95) <= 0; angryBirdLarge(138, 96) <= 0; angryBirdLarge(138, 97) <= 0; angryBirdLarge(138, 98) <= 0; angryBirdLarge(138, 99) <= 0; angryBirdLarge(138, 100) <= 0; angryBirdLarge(138, 101) <= 0; angryBirdLarge(138, 102) <= 0; angryBirdLarge(138, 103) <= 0; angryBirdLarge(138, 104) <= 0; angryBirdLarge(138, 105) <= 0; angryBirdLarge(138, 106) <= 0; angryBirdLarge(138, 107) <= 0; angryBirdLarge(138, 108) <= 0; angryBirdLarge(138, 109) <= 0; angryBirdLarge(138, 110) <= 0; angryBirdLarge(138, 111) <= 0; angryBirdLarge(138, 112) <= 0; angryBirdLarge(138, 113) <= 0; angryBirdLarge(138, 114) <= 0; angryBirdLarge(138, 115) <= 0; angryBirdLarge(138, 116) <= 0; angryBirdLarge(138, 117) <= 0; angryBirdLarge(138, 118) <= 0; angryBirdLarge(138, 119) <= 0; angryBirdLarge(138, 120) <= 0; angryBirdLarge(138, 121) <= 0; angryBirdLarge(138, 122) <= 0; angryBirdLarge(138, 123) <= 0; angryBirdLarge(138, 124) <= 0; angryBirdLarge(138, 125) <= 0; angryBirdLarge(138, 126) <= 0; angryBirdLarge(138, 127) <= 0; angryBirdLarge(138, 128) <= 0; angryBirdLarge(138, 129) <= 0; angryBirdLarge(138, 130) <= 0; angryBirdLarge(138, 131) <= 0; angryBirdLarge(138, 132) <= 0; angryBirdLarge(138, 133) <= 0; angryBirdLarge(138, 134) <= 0; angryBirdLarge(138, 135) <= 0; angryBirdLarge(138, 136) <= 0; angryBirdLarge(138, 137) <= 0; angryBirdLarge(138, 138) <= 0; angryBirdLarge(138, 139) <= 0; angryBirdLarge(138, 140) <= 0; angryBirdLarge(138, 141) <= 0; angryBirdLarge(138, 142) <= 0; angryBirdLarge(138, 143) <= 0; angryBirdLarge(138, 144) <= 0; angryBirdLarge(138, 145) <= 0; angryBirdLarge(138, 146) <= 0; angryBirdLarge(138, 147) <= 0; angryBirdLarge(138, 148) <= 0; angryBirdLarge(138, 149) <= 0; 
angryBirdLarge(139, 0) <= 0; angryBirdLarge(139, 1) <= 0; angryBirdLarge(139, 2) <= 0; angryBirdLarge(139, 3) <= 0; angryBirdLarge(139, 4) <= 0; angryBirdLarge(139, 5) <= 0; angryBirdLarge(139, 6) <= 0; angryBirdLarge(139, 7) <= 0; angryBirdLarge(139, 8) <= 0; angryBirdLarge(139, 9) <= 0; angryBirdLarge(139, 10) <= 0; angryBirdLarge(139, 11) <= 0; angryBirdLarge(139, 12) <= 0; angryBirdLarge(139, 13) <= 0; angryBirdLarge(139, 14) <= 0; angryBirdLarge(139, 15) <= 0; angryBirdLarge(139, 16) <= 0; angryBirdLarge(139, 17) <= 0; angryBirdLarge(139, 18) <= 0; angryBirdLarge(139, 19) <= 0; angryBirdLarge(139, 20) <= 0; angryBirdLarge(139, 21) <= 0; angryBirdLarge(139, 22) <= 0; angryBirdLarge(139, 23) <= 0; angryBirdLarge(139, 24) <= 0; angryBirdLarge(139, 25) <= 0; angryBirdLarge(139, 26) <= 0; angryBirdLarge(139, 27) <= 0; angryBirdLarge(139, 28) <= 0; angryBirdLarge(139, 29) <= 0; angryBirdLarge(139, 30) <= 0; angryBirdLarge(139, 31) <= 0; angryBirdLarge(139, 32) <= 0; angryBirdLarge(139, 33) <= 0; angryBirdLarge(139, 34) <= 0; angryBirdLarge(139, 35) <= 0; angryBirdLarge(139, 36) <= 0; angryBirdLarge(139, 37) <= 0; angryBirdLarge(139, 38) <= 0; angryBirdLarge(139, 39) <= 0; angryBirdLarge(139, 40) <= 0; angryBirdLarge(139, 41) <= 0; angryBirdLarge(139, 42) <= 0; angryBirdLarge(139, 43) <= 0; angryBirdLarge(139, 44) <= 0; angryBirdLarge(139, 45) <= 0; angryBirdLarge(139, 46) <= 0; angryBirdLarge(139, 47) <= 0; angryBirdLarge(139, 48) <= 0; angryBirdLarge(139, 49) <= 0; angryBirdLarge(139, 50) <= 0; angryBirdLarge(139, 51) <= 0; angryBirdLarge(139, 52) <= 0; angryBirdLarge(139, 53) <= 0; angryBirdLarge(139, 54) <= 0; angryBirdLarge(139, 55) <= 0; angryBirdLarge(139, 56) <= 0; angryBirdLarge(139, 57) <= 0; angryBirdLarge(139, 58) <= 0; angryBirdLarge(139, 59) <= 0; angryBirdLarge(139, 60) <= 0; angryBirdLarge(139, 61) <= 0; angryBirdLarge(139, 62) <= 0; angryBirdLarge(139, 63) <= 0; angryBirdLarge(139, 64) <= 0; angryBirdLarge(139, 65) <= 0; angryBirdLarge(139, 66) <= 0; angryBirdLarge(139, 67) <= 0; angryBirdLarge(139, 68) <= 0; angryBirdLarge(139, 69) <= 0; angryBirdLarge(139, 70) <= 0; angryBirdLarge(139, 71) <= 0; angryBirdLarge(139, 72) <= 0; angryBirdLarge(139, 73) <= 0; angryBirdLarge(139, 74) <= 0; angryBirdLarge(139, 75) <= 0; angryBirdLarge(139, 76) <= 0; angryBirdLarge(139, 77) <= 0; angryBirdLarge(139, 78) <= 0; angryBirdLarge(139, 79) <= 0; angryBirdLarge(139, 80) <= 0; angryBirdLarge(139, 81) <= 0; angryBirdLarge(139, 82) <= 0; angryBirdLarge(139, 83) <= 0; angryBirdLarge(139, 84) <= 0; angryBirdLarge(139, 85) <= 0; angryBirdLarge(139, 86) <= 0; angryBirdLarge(139, 87) <= 0; angryBirdLarge(139, 88) <= 0; angryBirdLarge(139, 89) <= 0; angryBirdLarge(139, 90) <= 0; angryBirdLarge(139, 91) <= 0; angryBirdLarge(139, 92) <= 0; angryBirdLarge(139, 93) <= 0; angryBirdLarge(139, 94) <= 0; angryBirdLarge(139, 95) <= 0; angryBirdLarge(139, 96) <= 0; angryBirdLarge(139, 97) <= 0; angryBirdLarge(139, 98) <= 0; angryBirdLarge(139, 99) <= 0; angryBirdLarge(139, 100) <= 0; angryBirdLarge(139, 101) <= 0; angryBirdLarge(139, 102) <= 0; angryBirdLarge(139, 103) <= 0; angryBirdLarge(139, 104) <= 0; angryBirdLarge(139, 105) <= 0; angryBirdLarge(139, 106) <= 0; angryBirdLarge(139, 107) <= 0; angryBirdLarge(139, 108) <= 0; angryBirdLarge(139, 109) <= 0; angryBirdLarge(139, 110) <= 0; angryBirdLarge(139, 111) <= 0; angryBirdLarge(139, 112) <= 0; angryBirdLarge(139, 113) <= 0; angryBirdLarge(139, 114) <= 0; angryBirdLarge(139, 115) <= 0; angryBirdLarge(139, 116) <= 0; angryBirdLarge(139, 117) <= 0; angryBirdLarge(139, 118) <= 0; angryBirdLarge(139, 119) <= 0; angryBirdLarge(139, 120) <= 0; angryBirdLarge(139, 121) <= 0; angryBirdLarge(139, 122) <= 0; angryBirdLarge(139, 123) <= 0; angryBirdLarge(139, 124) <= 0; angryBirdLarge(139, 125) <= 0; angryBirdLarge(139, 126) <= 0; angryBirdLarge(139, 127) <= 0; angryBirdLarge(139, 128) <= 0; angryBirdLarge(139, 129) <= 0; angryBirdLarge(139, 130) <= 0; angryBirdLarge(139, 131) <= 0; angryBirdLarge(139, 132) <= 0; angryBirdLarge(139, 133) <= 0; angryBirdLarge(139, 134) <= 0; angryBirdLarge(139, 135) <= 0; angryBirdLarge(139, 136) <= 0; angryBirdLarge(139, 137) <= 0; angryBirdLarge(139, 138) <= 0; angryBirdLarge(139, 139) <= 0; angryBirdLarge(139, 140) <= 0; angryBirdLarge(139, 141) <= 0; angryBirdLarge(139, 142) <= 0; angryBirdLarge(139, 143) <= 0; angryBirdLarge(139, 144) <= 0; angryBirdLarge(139, 145) <= 0; angryBirdLarge(139, 146) <= 0; angryBirdLarge(139, 147) <= 0; angryBirdLarge(139, 148) <= 0; angryBirdLarge(139, 149) <= 0; 
angryBirdLarge(140, 0) <= 0; angryBirdLarge(140, 1) <= 0; angryBirdLarge(140, 2) <= 0; angryBirdLarge(140, 3) <= 0; angryBirdLarge(140, 4) <= 0; angryBirdLarge(140, 5) <= 0; angryBirdLarge(140, 6) <= 0; angryBirdLarge(140, 7) <= 0; angryBirdLarge(140, 8) <= 0; angryBirdLarge(140, 9) <= 0; angryBirdLarge(140, 10) <= 0; angryBirdLarge(140, 11) <= 0; angryBirdLarge(140, 12) <= 0; angryBirdLarge(140, 13) <= 0; angryBirdLarge(140, 14) <= 0; angryBirdLarge(140, 15) <= 0; angryBirdLarge(140, 16) <= 0; angryBirdLarge(140, 17) <= 0; angryBirdLarge(140, 18) <= 0; angryBirdLarge(140, 19) <= 0; angryBirdLarge(140, 20) <= 0; angryBirdLarge(140, 21) <= 0; angryBirdLarge(140, 22) <= 0; angryBirdLarge(140, 23) <= 0; angryBirdLarge(140, 24) <= 0; angryBirdLarge(140, 25) <= 0; angryBirdLarge(140, 26) <= 0; angryBirdLarge(140, 27) <= 0; angryBirdLarge(140, 28) <= 0; angryBirdLarge(140, 29) <= 0; angryBirdLarge(140, 30) <= 0; angryBirdLarge(140, 31) <= 0; angryBirdLarge(140, 32) <= 0; angryBirdLarge(140, 33) <= 0; angryBirdLarge(140, 34) <= 0; angryBirdLarge(140, 35) <= 0; angryBirdLarge(140, 36) <= 0; angryBirdLarge(140, 37) <= 0; angryBirdLarge(140, 38) <= 0; angryBirdLarge(140, 39) <= 0; angryBirdLarge(140, 40) <= 0; angryBirdLarge(140, 41) <= 0; angryBirdLarge(140, 42) <= 0; angryBirdLarge(140, 43) <= 0; angryBirdLarge(140, 44) <= 0; angryBirdLarge(140, 45) <= 0; angryBirdLarge(140, 46) <= 0; angryBirdLarge(140, 47) <= 0; angryBirdLarge(140, 48) <= 0; angryBirdLarge(140, 49) <= 0; angryBirdLarge(140, 50) <= 0; angryBirdLarge(140, 51) <= 0; angryBirdLarge(140, 52) <= 0; angryBirdLarge(140, 53) <= 0; angryBirdLarge(140, 54) <= 0; angryBirdLarge(140, 55) <= 0; angryBirdLarge(140, 56) <= 0; angryBirdLarge(140, 57) <= 0; angryBirdLarge(140, 58) <= 0; angryBirdLarge(140, 59) <= 0; angryBirdLarge(140, 60) <= 0; angryBirdLarge(140, 61) <= 0; angryBirdLarge(140, 62) <= 0; angryBirdLarge(140, 63) <= 0; angryBirdLarge(140, 64) <= 0; angryBirdLarge(140, 65) <= 0; angryBirdLarge(140, 66) <= 0; angryBirdLarge(140, 67) <= 0; angryBirdLarge(140, 68) <= 0; angryBirdLarge(140, 69) <= 0; angryBirdLarge(140, 70) <= 0; angryBirdLarge(140, 71) <= 0; angryBirdLarge(140, 72) <= 0; angryBirdLarge(140, 73) <= 0; angryBirdLarge(140, 74) <= 0; angryBirdLarge(140, 75) <= 0; angryBirdLarge(140, 76) <= 0; angryBirdLarge(140, 77) <= 0; angryBirdLarge(140, 78) <= 0; angryBirdLarge(140, 79) <= 0; angryBirdLarge(140, 80) <= 0; angryBirdLarge(140, 81) <= 0; angryBirdLarge(140, 82) <= 0; angryBirdLarge(140, 83) <= 0; angryBirdLarge(140, 84) <= 0; angryBirdLarge(140, 85) <= 0; angryBirdLarge(140, 86) <= 0; angryBirdLarge(140, 87) <= 0; angryBirdLarge(140, 88) <= 0; angryBirdLarge(140, 89) <= 0; angryBirdLarge(140, 90) <= 0; angryBirdLarge(140, 91) <= 0; angryBirdLarge(140, 92) <= 0; angryBirdLarge(140, 93) <= 0; angryBirdLarge(140, 94) <= 0; angryBirdLarge(140, 95) <= 0; angryBirdLarge(140, 96) <= 0; angryBirdLarge(140, 97) <= 0; angryBirdLarge(140, 98) <= 0; angryBirdLarge(140, 99) <= 0; angryBirdLarge(140, 100) <= 0; angryBirdLarge(140, 101) <= 0; angryBirdLarge(140, 102) <= 0; angryBirdLarge(140, 103) <= 0; angryBirdLarge(140, 104) <= 0; angryBirdLarge(140, 105) <= 0; angryBirdLarge(140, 106) <= 0; angryBirdLarge(140, 107) <= 0; angryBirdLarge(140, 108) <= 0; angryBirdLarge(140, 109) <= 0; angryBirdLarge(140, 110) <= 0; angryBirdLarge(140, 111) <= 0; angryBirdLarge(140, 112) <= 0; angryBirdLarge(140, 113) <= 0; angryBirdLarge(140, 114) <= 0; angryBirdLarge(140, 115) <= 0; angryBirdLarge(140, 116) <= 0; angryBirdLarge(140, 117) <= 0; angryBirdLarge(140, 118) <= 0; angryBirdLarge(140, 119) <= 0; angryBirdLarge(140, 120) <= 0; angryBirdLarge(140, 121) <= 0; angryBirdLarge(140, 122) <= 0; angryBirdLarge(140, 123) <= 0; angryBirdLarge(140, 124) <= 0; angryBirdLarge(140, 125) <= 0; angryBirdLarge(140, 126) <= 0; angryBirdLarge(140, 127) <= 0; angryBirdLarge(140, 128) <= 0; angryBirdLarge(140, 129) <= 0; angryBirdLarge(140, 130) <= 0; angryBirdLarge(140, 131) <= 0; angryBirdLarge(140, 132) <= 0; angryBirdLarge(140, 133) <= 0; angryBirdLarge(140, 134) <= 0; angryBirdLarge(140, 135) <= 0; angryBirdLarge(140, 136) <= 0; angryBirdLarge(140, 137) <= 0; angryBirdLarge(140, 138) <= 0; angryBirdLarge(140, 139) <= 0; angryBirdLarge(140, 140) <= 0; angryBirdLarge(140, 141) <= 0; angryBirdLarge(140, 142) <= 0; angryBirdLarge(140, 143) <= 0; angryBirdLarge(140, 144) <= 0; angryBirdLarge(140, 145) <= 0; angryBirdLarge(140, 146) <= 0; angryBirdLarge(140, 147) <= 0; angryBirdLarge(140, 148) <= 0; angryBirdLarge(140, 149) <= 0; 
angryBirdLarge(141, 0) <= 0; angryBirdLarge(141, 1) <= 0; angryBirdLarge(141, 2) <= 0; angryBirdLarge(141, 3) <= 0; angryBirdLarge(141, 4) <= 0; angryBirdLarge(141, 5) <= 0; angryBirdLarge(141, 6) <= 0; angryBirdLarge(141, 7) <= 0; angryBirdLarge(141, 8) <= 0; angryBirdLarge(141, 9) <= 0; angryBirdLarge(141, 10) <= 0; angryBirdLarge(141, 11) <= 0; angryBirdLarge(141, 12) <= 0; angryBirdLarge(141, 13) <= 0; angryBirdLarge(141, 14) <= 0; angryBirdLarge(141, 15) <= 0; angryBirdLarge(141, 16) <= 0; angryBirdLarge(141, 17) <= 0; angryBirdLarge(141, 18) <= 0; angryBirdLarge(141, 19) <= 0; angryBirdLarge(141, 20) <= 0; angryBirdLarge(141, 21) <= 0; angryBirdLarge(141, 22) <= 0; angryBirdLarge(141, 23) <= 0; angryBirdLarge(141, 24) <= 0; angryBirdLarge(141, 25) <= 0; angryBirdLarge(141, 26) <= 0; angryBirdLarge(141, 27) <= 0; angryBirdLarge(141, 28) <= 0; angryBirdLarge(141, 29) <= 0; angryBirdLarge(141, 30) <= 0; angryBirdLarge(141, 31) <= 0; angryBirdLarge(141, 32) <= 0; angryBirdLarge(141, 33) <= 0; angryBirdLarge(141, 34) <= 0; angryBirdLarge(141, 35) <= 0; angryBirdLarge(141, 36) <= 0; angryBirdLarge(141, 37) <= 0; angryBirdLarge(141, 38) <= 0; angryBirdLarge(141, 39) <= 0; angryBirdLarge(141, 40) <= 0; angryBirdLarge(141, 41) <= 0; angryBirdLarge(141, 42) <= 0; angryBirdLarge(141, 43) <= 0; angryBirdLarge(141, 44) <= 0; angryBirdLarge(141, 45) <= 0; angryBirdLarge(141, 46) <= 0; angryBirdLarge(141, 47) <= 0; angryBirdLarge(141, 48) <= 0; angryBirdLarge(141, 49) <= 0; angryBirdLarge(141, 50) <= 0; angryBirdLarge(141, 51) <= 0; angryBirdLarge(141, 52) <= 0; angryBirdLarge(141, 53) <= 0; angryBirdLarge(141, 54) <= 0; angryBirdLarge(141, 55) <= 0; angryBirdLarge(141, 56) <= 0; angryBirdLarge(141, 57) <= 0; angryBirdLarge(141, 58) <= 0; angryBirdLarge(141, 59) <= 0; angryBirdLarge(141, 60) <= 0; angryBirdLarge(141, 61) <= 0; angryBirdLarge(141, 62) <= 0; angryBirdLarge(141, 63) <= 0; angryBirdLarge(141, 64) <= 0; angryBirdLarge(141, 65) <= 0; angryBirdLarge(141, 66) <= 0; angryBirdLarge(141, 67) <= 0; angryBirdLarge(141, 68) <= 0; angryBirdLarge(141, 69) <= 0; angryBirdLarge(141, 70) <= 0; angryBirdLarge(141, 71) <= 0; angryBirdLarge(141, 72) <= 0; angryBirdLarge(141, 73) <= 0; angryBirdLarge(141, 74) <= 0; angryBirdLarge(141, 75) <= 0; angryBirdLarge(141, 76) <= 0; angryBirdLarge(141, 77) <= 0; angryBirdLarge(141, 78) <= 0; angryBirdLarge(141, 79) <= 0; angryBirdLarge(141, 80) <= 0; angryBirdLarge(141, 81) <= 0; angryBirdLarge(141, 82) <= 0; angryBirdLarge(141, 83) <= 0; angryBirdLarge(141, 84) <= 0; angryBirdLarge(141, 85) <= 0; angryBirdLarge(141, 86) <= 0; angryBirdLarge(141, 87) <= 0; angryBirdLarge(141, 88) <= 0; angryBirdLarge(141, 89) <= 0; angryBirdLarge(141, 90) <= 0; angryBirdLarge(141, 91) <= 0; angryBirdLarge(141, 92) <= 0; angryBirdLarge(141, 93) <= 0; angryBirdLarge(141, 94) <= 0; angryBirdLarge(141, 95) <= 0; angryBirdLarge(141, 96) <= 0; angryBirdLarge(141, 97) <= 0; angryBirdLarge(141, 98) <= 0; angryBirdLarge(141, 99) <= 0; angryBirdLarge(141, 100) <= 0; angryBirdLarge(141, 101) <= 0; angryBirdLarge(141, 102) <= 0; angryBirdLarge(141, 103) <= 0; angryBirdLarge(141, 104) <= 0; angryBirdLarge(141, 105) <= 0; angryBirdLarge(141, 106) <= 0; angryBirdLarge(141, 107) <= 0; angryBirdLarge(141, 108) <= 0; angryBirdLarge(141, 109) <= 0; angryBirdLarge(141, 110) <= 0; angryBirdLarge(141, 111) <= 0; angryBirdLarge(141, 112) <= 0; angryBirdLarge(141, 113) <= 0; angryBirdLarge(141, 114) <= 0; angryBirdLarge(141, 115) <= 0; angryBirdLarge(141, 116) <= 0; angryBirdLarge(141, 117) <= 0; angryBirdLarge(141, 118) <= 0; angryBirdLarge(141, 119) <= 0; angryBirdLarge(141, 120) <= 0; angryBirdLarge(141, 121) <= 0; angryBirdLarge(141, 122) <= 0; angryBirdLarge(141, 123) <= 0; angryBirdLarge(141, 124) <= 0; angryBirdLarge(141, 125) <= 0; angryBirdLarge(141, 126) <= 0; angryBirdLarge(141, 127) <= 0; angryBirdLarge(141, 128) <= 0; angryBirdLarge(141, 129) <= 0; angryBirdLarge(141, 130) <= 0; angryBirdLarge(141, 131) <= 0; angryBirdLarge(141, 132) <= 0; angryBirdLarge(141, 133) <= 0; angryBirdLarge(141, 134) <= 0; angryBirdLarge(141, 135) <= 0; angryBirdLarge(141, 136) <= 0; angryBirdLarge(141, 137) <= 0; angryBirdLarge(141, 138) <= 0; angryBirdLarge(141, 139) <= 0; angryBirdLarge(141, 140) <= 0; angryBirdLarge(141, 141) <= 0; angryBirdLarge(141, 142) <= 0; angryBirdLarge(141, 143) <= 0; angryBirdLarge(141, 144) <= 0; angryBirdLarge(141, 145) <= 0; angryBirdLarge(141, 146) <= 0; angryBirdLarge(141, 147) <= 0; angryBirdLarge(141, 148) <= 0; angryBirdLarge(141, 149) <= 0; 
angryBirdLarge(142, 0) <= 0; angryBirdLarge(142, 1) <= 0; angryBirdLarge(142, 2) <= 0; angryBirdLarge(142, 3) <= 0; angryBirdLarge(142, 4) <= 0; angryBirdLarge(142, 5) <= 0; angryBirdLarge(142, 6) <= 0; angryBirdLarge(142, 7) <= 0; angryBirdLarge(142, 8) <= 0; angryBirdLarge(142, 9) <= 0; angryBirdLarge(142, 10) <= 0; angryBirdLarge(142, 11) <= 0; angryBirdLarge(142, 12) <= 0; angryBirdLarge(142, 13) <= 0; angryBirdLarge(142, 14) <= 0; angryBirdLarge(142, 15) <= 0; angryBirdLarge(142, 16) <= 0; angryBirdLarge(142, 17) <= 0; angryBirdLarge(142, 18) <= 0; angryBirdLarge(142, 19) <= 0; angryBirdLarge(142, 20) <= 0; angryBirdLarge(142, 21) <= 0; angryBirdLarge(142, 22) <= 0; angryBirdLarge(142, 23) <= 0; angryBirdLarge(142, 24) <= 0; angryBirdLarge(142, 25) <= 0; angryBirdLarge(142, 26) <= 0; angryBirdLarge(142, 27) <= 0; angryBirdLarge(142, 28) <= 0; angryBirdLarge(142, 29) <= 0; angryBirdLarge(142, 30) <= 0; angryBirdLarge(142, 31) <= 0; angryBirdLarge(142, 32) <= 0; angryBirdLarge(142, 33) <= 0; angryBirdLarge(142, 34) <= 0; angryBirdLarge(142, 35) <= 0; angryBirdLarge(142, 36) <= 0; angryBirdLarge(142, 37) <= 0; angryBirdLarge(142, 38) <= 0; angryBirdLarge(142, 39) <= 0; angryBirdLarge(142, 40) <= 0; angryBirdLarge(142, 41) <= 0; angryBirdLarge(142, 42) <= 0; angryBirdLarge(142, 43) <= 0; angryBirdLarge(142, 44) <= 0; angryBirdLarge(142, 45) <= 0; angryBirdLarge(142, 46) <= 0; angryBirdLarge(142, 47) <= 0; angryBirdLarge(142, 48) <= 0; angryBirdLarge(142, 49) <= 0; angryBirdLarge(142, 50) <= 0; angryBirdLarge(142, 51) <= 0; angryBirdLarge(142, 52) <= 0; angryBirdLarge(142, 53) <= 0; angryBirdLarge(142, 54) <= 0; angryBirdLarge(142, 55) <= 0; angryBirdLarge(142, 56) <= 0; angryBirdLarge(142, 57) <= 0; angryBirdLarge(142, 58) <= 0; angryBirdLarge(142, 59) <= 0; angryBirdLarge(142, 60) <= 0; angryBirdLarge(142, 61) <= 0; angryBirdLarge(142, 62) <= 0; angryBirdLarge(142, 63) <= 0; angryBirdLarge(142, 64) <= 0; angryBirdLarge(142, 65) <= 0; angryBirdLarge(142, 66) <= 0; angryBirdLarge(142, 67) <= 0; angryBirdLarge(142, 68) <= 0; angryBirdLarge(142, 69) <= 0; angryBirdLarge(142, 70) <= 0; angryBirdLarge(142, 71) <= 0; angryBirdLarge(142, 72) <= 0; angryBirdLarge(142, 73) <= 0; angryBirdLarge(142, 74) <= 0; angryBirdLarge(142, 75) <= 0; angryBirdLarge(142, 76) <= 0; angryBirdLarge(142, 77) <= 0; angryBirdLarge(142, 78) <= 0; angryBirdLarge(142, 79) <= 0; angryBirdLarge(142, 80) <= 0; angryBirdLarge(142, 81) <= 0; angryBirdLarge(142, 82) <= 0; angryBirdLarge(142, 83) <= 0; angryBirdLarge(142, 84) <= 0; angryBirdLarge(142, 85) <= 0; angryBirdLarge(142, 86) <= 0; angryBirdLarge(142, 87) <= 0; angryBirdLarge(142, 88) <= 0; angryBirdLarge(142, 89) <= 0; angryBirdLarge(142, 90) <= 0; angryBirdLarge(142, 91) <= 0; angryBirdLarge(142, 92) <= 0; angryBirdLarge(142, 93) <= 0; angryBirdLarge(142, 94) <= 0; angryBirdLarge(142, 95) <= 0; angryBirdLarge(142, 96) <= 0; angryBirdLarge(142, 97) <= 0; angryBirdLarge(142, 98) <= 0; angryBirdLarge(142, 99) <= 0; angryBirdLarge(142, 100) <= 0; angryBirdLarge(142, 101) <= 0; angryBirdLarge(142, 102) <= 0; angryBirdLarge(142, 103) <= 0; angryBirdLarge(142, 104) <= 0; angryBirdLarge(142, 105) <= 0; angryBirdLarge(142, 106) <= 0; angryBirdLarge(142, 107) <= 0; angryBirdLarge(142, 108) <= 0; angryBirdLarge(142, 109) <= 0; angryBirdLarge(142, 110) <= 0; angryBirdLarge(142, 111) <= 0; angryBirdLarge(142, 112) <= 0; angryBirdLarge(142, 113) <= 0; angryBirdLarge(142, 114) <= 0; angryBirdLarge(142, 115) <= 0; angryBirdLarge(142, 116) <= 0; angryBirdLarge(142, 117) <= 0; angryBirdLarge(142, 118) <= 0; angryBirdLarge(142, 119) <= 0; angryBirdLarge(142, 120) <= 0; angryBirdLarge(142, 121) <= 0; angryBirdLarge(142, 122) <= 0; angryBirdLarge(142, 123) <= 0; angryBirdLarge(142, 124) <= 0; angryBirdLarge(142, 125) <= 0; angryBirdLarge(142, 126) <= 0; angryBirdLarge(142, 127) <= 0; angryBirdLarge(142, 128) <= 0; angryBirdLarge(142, 129) <= 0; angryBirdLarge(142, 130) <= 0; angryBirdLarge(142, 131) <= 0; angryBirdLarge(142, 132) <= 0; angryBirdLarge(142, 133) <= 0; angryBirdLarge(142, 134) <= 0; angryBirdLarge(142, 135) <= 0; angryBirdLarge(142, 136) <= 0; angryBirdLarge(142, 137) <= 0; angryBirdLarge(142, 138) <= 0; angryBirdLarge(142, 139) <= 0; angryBirdLarge(142, 140) <= 0; angryBirdLarge(142, 141) <= 0; angryBirdLarge(142, 142) <= 0; angryBirdLarge(142, 143) <= 0; angryBirdLarge(142, 144) <= 0; angryBirdLarge(142, 145) <= 0; angryBirdLarge(142, 146) <= 0; angryBirdLarge(142, 147) <= 0; angryBirdLarge(142, 148) <= 0; angryBirdLarge(142, 149) <= 0; 
angryBirdLarge(143, 0) <= 0; angryBirdLarge(143, 1) <= 0; angryBirdLarge(143, 2) <= 0; angryBirdLarge(143, 3) <= 0; angryBirdLarge(143, 4) <= 0; angryBirdLarge(143, 5) <= 0; angryBirdLarge(143, 6) <= 0; angryBirdLarge(143, 7) <= 0; angryBirdLarge(143, 8) <= 0; angryBirdLarge(143, 9) <= 0; angryBirdLarge(143, 10) <= 0; angryBirdLarge(143, 11) <= 0; angryBirdLarge(143, 12) <= 0; angryBirdLarge(143, 13) <= 0; angryBirdLarge(143, 14) <= 0; angryBirdLarge(143, 15) <= 0; angryBirdLarge(143, 16) <= 0; angryBirdLarge(143, 17) <= 0; angryBirdLarge(143, 18) <= 0; angryBirdLarge(143, 19) <= 0; angryBirdLarge(143, 20) <= 0; angryBirdLarge(143, 21) <= 0; angryBirdLarge(143, 22) <= 0; angryBirdLarge(143, 23) <= 0; angryBirdLarge(143, 24) <= 0; angryBirdLarge(143, 25) <= 0; angryBirdLarge(143, 26) <= 0; angryBirdLarge(143, 27) <= 0; angryBirdLarge(143, 28) <= 0; angryBirdLarge(143, 29) <= 0; angryBirdLarge(143, 30) <= 0; angryBirdLarge(143, 31) <= 0; angryBirdLarge(143, 32) <= 0; angryBirdLarge(143, 33) <= 0; angryBirdLarge(143, 34) <= 0; angryBirdLarge(143, 35) <= 0; angryBirdLarge(143, 36) <= 0; angryBirdLarge(143, 37) <= 0; angryBirdLarge(143, 38) <= 0; angryBirdLarge(143, 39) <= 0; angryBirdLarge(143, 40) <= 0; angryBirdLarge(143, 41) <= 0; angryBirdLarge(143, 42) <= 0; angryBirdLarge(143, 43) <= 0; angryBirdLarge(143, 44) <= 0; angryBirdLarge(143, 45) <= 0; angryBirdLarge(143, 46) <= 0; angryBirdLarge(143, 47) <= 0; angryBirdLarge(143, 48) <= 0; angryBirdLarge(143, 49) <= 0; angryBirdLarge(143, 50) <= 0; angryBirdLarge(143, 51) <= 0; angryBirdLarge(143, 52) <= 0; angryBirdLarge(143, 53) <= 0; angryBirdLarge(143, 54) <= 0; angryBirdLarge(143, 55) <= 0; angryBirdLarge(143, 56) <= 0; angryBirdLarge(143, 57) <= 0; angryBirdLarge(143, 58) <= 0; angryBirdLarge(143, 59) <= 0; angryBirdLarge(143, 60) <= 0; angryBirdLarge(143, 61) <= 0; angryBirdLarge(143, 62) <= 0; angryBirdLarge(143, 63) <= 0; angryBirdLarge(143, 64) <= 0; angryBirdLarge(143, 65) <= 0; angryBirdLarge(143, 66) <= 0; angryBirdLarge(143, 67) <= 0; angryBirdLarge(143, 68) <= 0; angryBirdLarge(143, 69) <= 0; angryBirdLarge(143, 70) <= 0; angryBirdLarge(143, 71) <= 0; angryBirdLarge(143, 72) <= 0; angryBirdLarge(143, 73) <= 0; angryBirdLarge(143, 74) <= 0; angryBirdLarge(143, 75) <= 0; angryBirdLarge(143, 76) <= 0; angryBirdLarge(143, 77) <= 0; angryBirdLarge(143, 78) <= 0; angryBirdLarge(143, 79) <= 0; angryBirdLarge(143, 80) <= 0; angryBirdLarge(143, 81) <= 0; angryBirdLarge(143, 82) <= 0; angryBirdLarge(143, 83) <= 0; angryBirdLarge(143, 84) <= 0; angryBirdLarge(143, 85) <= 0; angryBirdLarge(143, 86) <= 0; angryBirdLarge(143, 87) <= 0; angryBirdLarge(143, 88) <= 0; angryBirdLarge(143, 89) <= 0; angryBirdLarge(143, 90) <= 0; angryBirdLarge(143, 91) <= 0; angryBirdLarge(143, 92) <= 0; angryBirdLarge(143, 93) <= 0; angryBirdLarge(143, 94) <= 0; angryBirdLarge(143, 95) <= 0; angryBirdLarge(143, 96) <= 0; angryBirdLarge(143, 97) <= 0; angryBirdLarge(143, 98) <= 0; angryBirdLarge(143, 99) <= 0; angryBirdLarge(143, 100) <= 0; angryBirdLarge(143, 101) <= 0; angryBirdLarge(143, 102) <= 0; angryBirdLarge(143, 103) <= 0; angryBirdLarge(143, 104) <= 0; angryBirdLarge(143, 105) <= 0; angryBirdLarge(143, 106) <= 0; angryBirdLarge(143, 107) <= 0; angryBirdLarge(143, 108) <= 0; angryBirdLarge(143, 109) <= 0; angryBirdLarge(143, 110) <= 0; angryBirdLarge(143, 111) <= 0; angryBirdLarge(143, 112) <= 0; angryBirdLarge(143, 113) <= 0; angryBirdLarge(143, 114) <= 0; angryBirdLarge(143, 115) <= 0; angryBirdLarge(143, 116) <= 0; angryBirdLarge(143, 117) <= 0; angryBirdLarge(143, 118) <= 0; angryBirdLarge(143, 119) <= 0; angryBirdLarge(143, 120) <= 0; angryBirdLarge(143, 121) <= 0; angryBirdLarge(143, 122) <= 0; angryBirdLarge(143, 123) <= 0; angryBirdLarge(143, 124) <= 0; angryBirdLarge(143, 125) <= 0; angryBirdLarge(143, 126) <= 0; angryBirdLarge(143, 127) <= 0; angryBirdLarge(143, 128) <= 0; angryBirdLarge(143, 129) <= 0; angryBirdLarge(143, 130) <= 0; angryBirdLarge(143, 131) <= 0; angryBirdLarge(143, 132) <= 0; angryBirdLarge(143, 133) <= 0; angryBirdLarge(143, 134) <= 0; angryBirdLarge(143, 135) <= 0; angryBirdLarge(143, 136) <= 0; angryBirdLarge(143, 137) <= 0; angryBirdLarge(143, 138) <= 0; angryBirdLarge(143, 139) <= 0; angryBirdLarge(143, 140) <= 0; angryBirdLarge(143, 141) <= 0; angryBirdLarge(143, 142) <= 0; angryBirdLarge(143, 143) <= 0; angryBirdLarge(143, 144) <= 0; angryBirdLarge(143, 145) <= 0; angryBirdLarge(143, 146) <= 0; angryBirdLarge(143, 147) <= 0; angryBirdLarge(143, 148) <= 0; angryBirdLarge(143, 149) <= 0; 




end Behavioral;
