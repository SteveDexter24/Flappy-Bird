library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package playpkg is
    type play2D is array(0 to 29, 0 to 269) of integer;
end package;

use work.playpkg.all;

entity play is
    Port (play_W: out play2D);
end play;

architecture Behavioral of play is

begin

play_W(0, 0) <= 1; play_W(0, 1) <= 1; play_W(0, 2) <= 1; play_W(0, 3) <= 1; play_W(0, 4) <= 1; play_W(0, 5) <= 1; play_W(0, 6) <= 1; play_W(0, 7) <= 1; play_W(0, 8) <= 1; play_W(0, 9) <= 1; play_W(0, 10) <= 1; play_W(0, 11) <= 1; play_W(0, 12) <= 1; play_W(0, 13) <= 1; play_W(0, 14) <= 1; play_W(0, 15) <= 1; play_W(0, 16) <= 1; play_W(0, 17) <= 1; play_W(0, 18) <= 0; play_W(0, 19) <= 0; play_W(0, 20) <= 0; play_W(0, 21) <= 0; play_W(0, 22) <= 0; play_W(0, 23) <= 0; play_W(0, 24) <= 0; play_W(0, 25) <= 0; play_W(0, 26) <= 0; play_W(0, 27) <= 1; play_W(0, 28) <= 1; play_W(0, 29) <= 1; play_W(0, 30) <= 1; play_W(0, 31) <= 1; play_W(0, 32) <= 1; play_W(0, 33) <= 1; play_W(0, 34) <= 1; play_W(0, 35) <= 1; play_W(0, 36) <= 1; play_W(0, 37) <= 1; play_W(0, 38) <= 1; play_W(0, 39) <= 0; play_W(0, 40) <= 0; play_W(0, 41) <= 0; play_W(0, 42) <= 0; play_W(0, 43) <= 0; play_W(0, 44) <= 0; play_W(0, 45) <= 0; play_W(0, 46) <= 0; play_W(0, 47) <= 0; play_W(0, 48) <= 0; play_W(0, 49) <= 0; play_W(0, 50) <= 0; play_W(0, 51) <= 0; play_W(0, 52) <= 0; play_W(0, 53) <= 0; play_W(0, 54) <= 0; play_W(0, 55) <= 0; play_W(0, 56) <= 0; play_W(0, 57) <= 0; play_W(0, 58) <= 0; play_W(0, 59) <= 0; play_W(0, 60) <= 0; play_W(0, 61) <= 0; play_W(0, 62) <= 0; play_W(0, 63) <= 1; play_W(0, 64) <= 1; play_W(0, 65) <= 1; play_W(0, 66) <= 0; play_W(0, 67) <= 0; play_W(0, 68) <= 0; play_W(0, 69) <= 0; play_W(0, 70) <= 0; play_W(0, 71) <= 0; play_W(0, 72) <= 0; play_W(0, 73) <= 0; play_W(0, 74) <= 0; play_W(0, 75) <= 0; play_W(0, 76) <= 0; play_W(0, 77) <= 0; play_W(0, 78) <= 0; play_W(0, 79) <= 0; play_W(0, 80) <= 0; play_W(0, 81) <= 1; play_W(0, 82) <= 1; play_W(0, 83) <= 1; play_W(0, 84) <= 1; play_W(0, 85) <= 1; play_W(0, 86) <= 1; play_W(0, 87) <= 0; play_W(0, 88) <= 0; play_W(0, 89) <= 0; play_W(0, 90) <= 0; play_W(0, 91) <= 0; play_W(0, 92) <= 0; play_W(0, 93) <= 0; play_W(0, 94) <= 0; play_W(0, 95) <= 0; play_W(0, 96) <= 0; play_W(0, 97) <= 0; play_W(0, 98) <= 0; play_W(0, 99) <= 1; play_W(0, 100) <= 1; play_W(0, 101) <= 1; play_W(0, 102) <= 1; play_W(0, 103) <= 1; play_W(0, 104) <= 1; play_W(0, 105) <= 0; play_W(0, 106) <= 0; play_W(0, 107) <= 0; play_W(0, 108) <= 0; play_W(0, 109) <= 0; play_W(0, 110) <= 0; play_W(0, 111) <= 0; play_W(0, 112) <= 0; play_W(0, 113) <= 0; play_W(0, 114) <= 0; play_W(0, 115) <= 0; play_W(0, 116) <= 0; play_W(0, 117) <= 0; play_W(0, 118) <= 0; play_W(0, 119) <= 0; play_W(0, 120) <= 0; play_W(0, 121) <= 0; play_W(0, 122) <= 0; play_W(0, 123) <= 0; play_W(0, 124) <= 0; play_W(0, 125) <= 0; play_W(0, 126) <= 0; play_W(0, 127) <= 0; play_W(0, 128) <= 0; play_W(0, 129) <= 0; play_W(0, 130) <= 0; play_W(0, 131) <= 0; play_W(0, 132) <= 0; play_W(0, 133) <= 0; play_W(0, 134) <= 0; play_W(0, 135) <= 0; play_W(0, 136) <= 0; play_W(0, 137) <= 0; play_W(0, 138) <= 0; play_W(0, 139) <= 0; play_W(0, 140) <= 0; play_W(0, 141) <= 0; play_W(0, 142) <= 0; play_W(0, 143) <= 0; play_W(0, 144) <= 0; play_W(0, 145) <= 0; play_W(0, 146) <= 0; play_W(0, 147) <= 0; play_W(0, 148) <= 0; play_W(0, 149) <= 0; play_W(0, 150) <= 0; play_W(0, 151) <= 0; play_W(0, 152) <= 0; play_W(0, 153) <= 0; play_W(0, 154) <= 0; play_W(0, 155) <= 0; play_W(0, 156) <= 0; play_W(0, 157) <= 0; play_W(0, 158) <= 0; play_W(0, 159) <= 0; play_W(0, 160) <= 0; play_W(0, 161) <= 0; play_W(0, 162) <= 1; play_W(0, 163) <= 1; play_W(0, 164) <= 1; play_W(0, 165) <= 1; play_W(0, 166) <= 1; play_W(0, 167) <= 1; play_W(0, 168) <= 1; play_W(0, 169) <= 1; play_W(0, 170) <= 1; play_W(0, 171) <= 1; play_W(0, 172) <= 1; play_W(0, 173) <= 1; play_W(0, 174) <= 1; play_W(0, 175) <= 1; play_W(0, 176) <= 1; play_W(0, 177) <= 1; play_W(0, 178) <= 1; play_W(0, 179) <= 1; play_W(0, 180) <= 0; play_W(0, 181) <= 0; play_W(0, 182) <= 0; play_W(0, 183) <= 0; play_W(0, 184) <= 0; play_W(0, 185) <= 0; play_W(0, 186) <= 0; play_W(0, 187) <= 0; play_W(0, 188) <= 0; play_W(0, 189) <= 1; play_W(0, 190) <= 1; play_W(0, 191) <= 1; play_W(0, 192) <= 1; play_W(0, 193) <= 1; play_W(0, 194) <= 1; play_W(0, 195) <= 1; play_W(0, 196) <= 1; play_W(0, 197) <= 1; play_W(0, 198) <= 1; play_W(0, 199) <= 1; play_W(0, 200) <= 1; play_W(0, 201) <= 1; play_W(0, 202) <= 1; play_W(0, 203) <= 1; play_W(0, 204) <= 1; play_W(0, 205) <= 1; play_W(0, 206) <= 1; play_W(0, 207) <= 1; play_W(0, 208) <= 1; play_W(0, 209) <= 1; play_W(0, 210) <= 1; play_W(0, 211) <= 1; play_W(0, 212) <= 1; play_W(0, 213) <= 0; play_W(0, 214) <= 0; play_W(0, 215) <= 0; play_W(0, 216) <= 1; play_W(0, 217) <= 1; play_W(0, 218) <= 1; play_W(0, 219) <= 1; play_W(0, 220) <= 1; play_W(0, 221) <= 1; play_W(0, 222) <= 0; play_W(0, 223) <= 0; play_W(0, 224) <= 0; play_W(0, 225) <= 0; play_W(0, 226) <= 0; play_W(0, 227) <= 0; play_W(0, 228) <= 0; play_W(0, 229) <= 0; play_W(0, 230) <= 0; play_W(0, 231) <= 1; play_W(0, 232) <= 1; play_W(0, 233) <= 1; play_W(0, 234) <= 1; play_W(0, 235) <= 1; play_W(0, 236) <= 1; play_W(0, 237) <= 0; play_W(0, 238) <= 0; play_W(0, 239) <= 0; play_W(0, 240) <= 0; play_W(0, 241) <= 0; play_W(0, 242) <= 0; play_W(0, 243) <= 1; play_W(0, 244) <= 1; play_W(0, 245) <= 1; play_W(0, 246) <= 1; play_W(0, 247) <= 1; play_W(0, 248) <= 1; play_W(0, 249) <= 1; play_W(0, 250) <= 1; play_W(0, 251) <= 1; play_W(0, 252) <= 1; play_W(0, 253) <= 1; play_W(0, 254) <= 1; play_W(0, 255) <= 1; play_W(0, 256) <= 1; play_W(0, 257) <= 1; play_W(0, 258) <= 1; play_W(0, 259) <= 1; play_W(0, 260) <= 1; play_W(0, 261) <= 0; play_W(0, 262) <= 0; play_W(0, 263) <= 0; play_W(0, 264) <= 0; play_W(0, 265) <= 0; play_W(0, 266) <= 0; play_W(0, 267) <= 0; play_W(0, 268) <= 0; play_W(0, 269) <= 0; 
play_W(1, 0) <= 1; play_W(1, 1) <= 1; play_W(1, 2) <= 1; play_W(1, 3) <= 1; play_W(1, 4) <= 1; play_W(1, 5) <= 1; play_W(1, 6) <= 1; play_W(1, 7) <= 1; play_W(1, 8) <= 1; play_W(1, 9) <= 1; play_W(1, 10) <= 1; play_W(1, 11) <= 1; play_W(1, 12) <= 1; play_W(1, 13) <= 1; play_W(1, 14) <= 1; play_W(1, 15) <= 1; play_W(1, 16) <= 1; play_W(1, 17) <= 1; play_W(1, 18) <= 0; play_W(1, 19) <= 0; play_W(1, 20) <= 0; play_W(1, 21) <= 0; play_W(1, 22) <= 0; play_W(1, 23) <= 0; play_W(1, 24) <= 0; play_W(1, 25) <= 0; play_W(1, 26) <= 0; play_W(1, 27) <= 1; play_W(1, 28) <= 1; play_W(1, 29) <= 1; play_W(1, 30) <= 1; play_W(1, 31) <= 1; play_W(1, 32) <= 1; play_W(1, 33) <= 1; play_W(1, 34) <= 1; play_W(1, 35) <= 1; play_W(1, 36) <= 1; play_W(1, 37) <= 1; play_W(1, 38) <= 1; play_W(1, 39) <= 0; play_W(1, 40) <= 0; play_W(1, 41) <= 0; play_W(1, 42) <= 0; play_W(1, 43) <= 0; play_W(1, 44) <= 0; play_W(1, 45) <= 0; play_W(1, 46) <= 0; play_W(1, 47) <= 0; play_W(1, 48) <= 0; play_W(1, 49) <= 0; play_W(1, 50) <= 0; play_W(1, 51) <= 0; play_W(1, 52) <= 0; play_W(1, 53) <= 0; play_W(1, 54) <= 0; play_W(1, 55) <= 0; play_W(1, 56) <= 0; play_W(1, 57) <= 0; play_W(1, 58) <= 0; play_W(1, 59) <= 0; play_W(1, 60) <= 0; play_W(1, 61) <= 0; play_W(1, 62) <= 0; play_W(1, 63) <= 1; play_W(1, 64) <= 1; play_W(1, 65) <= 1; play_W(1, 66) <= 0; play_W(1, 67) <= 0; play_W(1, 68) <= 0; play_W(1, 69) <= 0; play_W(1, 70) <= 0; play_W(1, 71) <= 0; play_W(1, 72) <= 0; play_W(1, 73) <= 0; play_W(1, 74) <= 0; play_W(1, 75) <= 0; play_W(1, 76) <= 0; play_W(1, 77) <= 0; play_W(1, 78) <= 0; play_W(1, 79) <= 0; play_W(1, 80) <= 0; play_W(1, 81) <= 1; play_W(1, 82) <= 1; play_W(1, 83) <= 1; play_W(1, 84) <= 1; play_W(1, 85) <= 1; play_W(1, 86) <= 1; play_W(1, 87) <= 0; play_W(1, 88) <= 0; play_W(1, 89) <= 0; play_W(1, 90) <= 0; play_W(1, 91) <= 0; play_W(1, 92) <= 0; play_W(1, 93) <= 0; play_W(1, 94) <= 0; play_W(1, 95) <= 0; play_W(1, 96) <= 0; play_W(1, 97) <= 0; play_W(1, 98) <= 0; play_W(1, 99) <= 1; play_W(1, 100) <= 1; play_W(1, 101) <= 1; play_W(1, 102) <= 1; play_W(1, 103) <= 1; play_W(1, 104) <= 1; play_W(1, 105) <= 0; play_W(1, 106) <= 0; play_W(1, 107) <= 0; play_W(1, 108) <= 0; play_W(1, 109) <= 0; play_W(1, 110) <= 0; play_W(1, 111) <= 0; play_W(1, 112) <= 0; play_W(1, 113) <= 0; play_W(1, 114) <= 0; play_W(1, 115) <= 0; play_W(1, 116) <= 0; play_W(1, 117) <= 0; play_W(1, 118) <= 0; play_W(1, 119) <= 0; play_W(1, 120) <= 0; play_W(1, 121) <= 0; play_W(1, 122) <= 0; play_W(1, 123) <= 0; play_W(1, 124) <= 0; play_W(1, 125) <= 0; play_W(1, 126) <= 0; play_W(1, 127) <= 0; play_W(1, 128) <= 0; play_W(1, 129) <= 0; play_W(1, 130) <= 0; play_W(1, 131) <= 0; play_W(1, 132) <= 0; play_W(1, 133) <= 0; play_W(1, 134) <= 0; play_W(1, 135) <= 0; play_W(1, 136) <= 0; play_W(1, 137) <= 0; play_W(1, 138) <= 0; play_W(1, 139) <= 0; play_W(1, 140) <= 0; play_W(1, 141) <= 0; play_W(1, 142) <= 0; play_W(1, 143) <= 0; play_W(1, 144) <= 0; play_W(1, 145) <= 0; play_W(1, 146) <= 0; play_W(1, 147) <= 0; play_W(1, 148) <= 0; play_W(1, 149) <= 0; play_W(1, 150) <= 0; play_W(1, 151) <= 0; play_W(1, 152) <= 0; play_W(1, 153) <= 0; play_W(1, 154) <= 0; play_W(1, 155) <= 0; play_W(1, 156) <= 0; play_W(1, 157) <= 0; play_W(1, 158) <= 0; play_W(1, 159) <= 0; play_W(1, 160) <= 0; play_W(1, 161) <= 0; play_W(1, 162) <= 1; play_W(1, 163) <= 1; play_W(1, 164) <= 1; play_W(1, 165) <= 1; play_W(1, 166) <= 1; play_W(1, 167) <= 1; play_W(1, 168) <= 1; play_W(1, 169) <= 1; play_W(1, 170) <= 1; play_W(1, 171) <= 1; play_W(1, 172) <= 1; play_W(1, 173) <= 1; play_W(1, 174) <= 1; play_W(1, 175) <= 1; play_W(1, 176) <= 1; play_W(1, 177) <= 1; play_W(1, 178) <= 1; play_W(1, 179) <= 1; play_W(1, 180) <= 0; play_W(1, 181) <= 0; play_W(1, 182) <= 0; play_W(1, 183) <= 0; play_W(1, 184) <= 0; play_W(1, 185) <= 0; play_W(1, 186) <= 0; play_W(1, 187) <= 0; play_W(1, 188) <= 0; play_W(1, 189) <= 1; play_W(1, 190) <= 1; play_W(1, 191) <= 1; play_W(1, 192) <= 1; play_W(1, 193) <= 1; play_W(1, 194) <= 1; play_W(1, 195) <= 1; play_W(1, 196) <= 1; play_W(1, 197) <= 1; play_W(1, 198) <= 1; play_W(1, 199) <= 1; play_W(1, 200) <= 1; play_W(1, 201) <= 1; play_W(1, 202) <= 1; play_W(1, 203) <= 1; play_W(1, 204) <= 1; play_W(1, 205) <= 1; play_W(1, 206) <= 1; play_W(1, 207) <= 1; play_W(1, 208) <= 1; play_W(1, 209) <= 1; play_W(1, 210) <= 1; play_W(1, 211) <= 1; play_W(1, 212) <= 1; play_W(1, 213) <= 0; play_W(1, 214) <= 0; play_W(1, 215) <= 0; play_W(1, 216) <= 1; play_W(1, 217) <= 1; play_W(1, 218) <= 1; play_W(1, 219) <= 1; play_W(1, 220) <= 1; play_W(1, 221) <= 1; play_W(1, 222) <= 0; play_W(1, 223) <= 0; play_W(1, 224) <= 0; play_W(1, 225) <= 0; play_W(1, 226) <= 0; play_W(1, 227) <= 0; play_W(1, 228) <= 0; play_W(1, 229) <= 0; play_W(1, 230) <= 0; play_W(1, 231) <= 1; play_W(1, 232) <= 1; play_W(1, 233) <= 1; play_W(1, 234) <= 1; play_W(1, 235) <= 1; play_W(1, 236) <= 1; play_W(1, 237) <= 0; play_W(1, 238) <= 0; play_W(1, 239) <= 0; play_W(1, 240) <= 0; play_W(1, 241) <= 0; play_W(1, 242) <= 0; play_W(1, 243) <= 1; play_W(1, 244) <= 1; play_W(1, 245) <= 1; play_W(1, 246) <= 1; play_W(1, 247) <= 1; play_W(1, 248) <= 1; play_W(1, 249) <= 1; play_W(1, 250) <= 1; play_W(1, 251) <= 1; play_W(1, 252) <= 1; play_W(1, 253) <= 1; play_W(1, 254) <= 1; play_W(1, 255) <= 1; play_W(1, 256) <= 1; play_W(1, 257) <= 1; play_W(1, 258) <= 1; play_W(1, 259) <= 1; play_W(1, 260) <= 1; play_W(1, 261) <= 0; play_W(1, 262) <= 0; play_W(1, 263) <= 0; play_W(1, 264) <= 0; play_W(1, 265) <= 0; play_W(1, 266) <= 0; play_W(1, 267) <= 0; play_W(1, 268) <= 0; play_W(1, 269) <= 0; 
play_W(2, 0) <= 1; play_W(2, 1) <= 1; play_W(2, 2) <= 1; play_W(2, 3) <= 1; play_W(2, 4) <= 1; play_W(2, 5) <= 1; play_W(2, 6) <= 1; play_W(2, 7) <= 1; play_W(2, 8) <= 1; play_W(2, 9) <= 1; play_W(2, 10) <= 1; play_W(2, 11) <= 1; play_W(2, 12) <= 1; play_W(2, 13) <= 1; play_W(2, 14) <= 1; play_W(2, 15) <= 1; play_W(2, 16) <= 1; play_W(2, 17) <= 1; play_W(2, 18) <= 0; play_W(2, 19) <= 0; play_W(2, 20) <= 0; play_W(2, 21) <= 0; play_W(2, 22) <= 0; play_W(2, 23) <= 0; play_W(2, 24) <= 0; play_W(2, 25) <= 0; play_W(2, 26) <= 0; play_W(2, 27) <= 1; play_W(2, 28) <= 1; play_W(2, 29) <= 1; play_W(2, 30) <= 1; play_W(2, 31) <= 1; play_W(2, 32) <= 1; play_W(2, 33) <= 1; play_W(2, 34) <= 1; play_W(2, 35) <= 1; play_W(2, 36) <= 1; play_W(2, 37) <= 1; play_W(2, 38) <= 1; play_W(2, 39) <= 0; play_W(2, 40) <= 0; play_W(2, 41) <= 0; play_W(2, 42) <= 0; play_W(2, 43) <= 0; play_W(2, 44) <= 0; play_W(2, 45) <= 0; play_W(2, 46) <= 0; play_W(2, 47) <= 0; play_W(2, 48) <= 0; play_W(2, 49) <= 0; play_W(2, 50) <= 0; play_W(2, 51) <= 0; play_W(2, 52) <= 0; play_W(2, 53) <= 0; play_W(2, 54) <= 0; play_W(2, 55) <= 0; play_W(2, 56) <= 0; play_W(2, 57) <= 0; play_W(2, 58) <= 0; play_W(2, 59) <= 0; play_W(2, 60) <= 0; play_W(2, 61) <= 0; play_W(2, 62) <= 0; play_W(2, 63) <= 1; play_W(2, 64) <= 1; play_W(2, 65) <= 1; play_W(2, 66) <= 0; play_W(2, 67) <= 0; play_W(2, 68) <= 0; play_W(2, 69) <= 0; play_W(2, 70) <= 0; play_W(2, 71) <= 0; play_W(2, 72) <= 0; play_W(2, 73) <= 0; play_W(2, 74) <= 0; play_W(2, 75) <= 0; play_W(2, 76) <= 0; play_W(2, 77) <= 0; play_W(2, 78) <= 0; play_W(2, 79) <= 0; play_W(2, 80) <= 0; play_W(2, 81) <= 1; play_W(2, 82) <= 1; play_W(2, 83) <= 1; play_W(2, 84) <= 1; play_W(2, 85) <= 1; play_W(2, 86) <= 1; play_W(2, 87) <= 0; play_W(2, 88) <= 0; play_W(2, 89) <= 0; play_W(2, 90) <= 0; play_W(2, 91) <= 0; play_W(2, 92) <= 0; play_W(2, 93) <= 0; play_W(2, 94) <= 0; play_W(2, 95) <= 0; play_W(2, 96) <= 0; play_W(2, 97) <= 0; play_W(2, 98) <= 0; play_W(2, 99) <= 1; play_W(2, 100) <= 1; play_W(2, 101) <= 1; play_W(2, 102) <= 1; play_W(2, 103) <= 1; play_W(2, 104) <= 1; play_W(2, 105) <= 0; play_W(2, 106) <= 0; play_W(2, 107) <= 0; play_W(2, 108) <= 0; play_W(2, 109) <= 0; play_W(2, 110) <= 0; play_W(2, 111) <= 0; play_W(2, 112) <= 0; play_W(2, 113) <= 0; play_W(2, 114) <= 0; play_W(2, 115) <= 0; play_W(2, 116) <= 0; play_W(2, 117) <= 0; play_W(2, 118) <= 0; play_W(2, 119) <= 0; play_W(2, 120) <= 0; play_W(2, 121) <= 0; play_W(2, 122) <= 0; play_W(2, 123) <= 0; play_W(2, 124) <= 0; play_W(2, 125) <= 0; play_W(2, 126) <= 0; play_W(2, 127) <= 0; play_W(2, 128) <= 0; play_W(2, 129) <= 0; play_W(2, 130) <= 0; play_W(2, 131) <= 0; play_W(2, 132) <= 0; play_W(2, 133) <= 0; play_W(2, 134) <= 0; play_W(2, 135) <= 0; play_W(2, 136) <= 0; play_W(2, 137) <= 0; play_W(2, 138) <= 0; play_W(2, 139) <= 0; play_W(2, 140) <= 0; play_W(2, 141) <= 0; play_W(2, 142) <= 0; play_W(2, 143) <= 0; play_W(2, 144) <= 0; play_W(2, 145) <= 0; play_W(2, 146) <= 0; play_W(2, 147) <= 0; play_W(2, 148) <= 0; play_W(2, 149) <= 0; play_W(2, 150) <= 0; play_W(2, 151) <= 0; play_W(2, 152) <= 0; play_W(2, 153) <= 0; play_W(2, 154) <= 0; play_W(2, 155) <= 0; play_W(2, 156) <= 0; play_W(2, 157) <= 0; play_W(2, 158) <= 0; play_W(2, 159) <= 0; play_W(2, 160) <= 0; play_W(2, 161) <= 0; play_W(2, 162) <= 1; play_W(2, 163) <= 1; play_W(2, 164) <= 1; play_W(2, 165) <= 1; play_W(2, 166) <= 1; play_W(2, 167) <= 1; play_W(2, 168) <= 1; play_W(2, 169) <= 1; play_W(2, 170) <= 1; play_W(2, 171) <= 1; play_W(2, 172) <= 1; play_W(2, 173) <= 1; play_W(2, 174) <= 1; play_W(2, 175) <= 1; play_W(2, 176) <= 1; play_W(2, 177) <= 1; play_W(2, 178) <= 1; play_W(2, 179) <= 1; play_W(2, 180) <= 0; play_W(2, 181) <= 0; play_W(2, 182) <= 0; play_W(2, 183) <= 0; play_W(2, 184) <= 0; play_W(2, 185) <= 0; play_W(2, 186) <= 0; play_W(2, 187) <= 0; play_W(2, 188) <= 0; play_W(2, 189) <= 1; play_W(2, 190) <= 1; play_W(2, 191) <= 1; play_W(2, 192) <= 1; play_W(2, 193) <= 1; play_W(2, 194) <= 1; play_W(2, 195) <= 1; play_W(2, 196) <= 1; play_W(2, 197) <= 1; play_W(2, 198) <= 1; play_W(2, 199) <= 1; play_W(2, 200) <= 1; play_W(2, 201) <= 1; play_W(2, 202) <= 1; play_W(2, 203) <= 1; play_W(2, 204) <= 1; play_W(2, 205) <= 1; play_W(2, 206) <= 1; play_W(2, 207) <= 1; play_W(2, 208) <= 1; play_W(2, 209) <= 1; play_W(2, 210) <= 1; play_W(2, 211) <= 1; play_W(2, 212) <= 1; play_W(2, 213) <= 0; play_W(2, 214) <= 0; play_W(2, 215) <= 0; play_W(2, 216) <= 1; play_W(2, 217) <= 1; play_W(2, 218) <= 1; play_W(2, 219) <= 1; play_W(2, 220) <= 1; play_W(2, 221) <= 1; play_W(2, 222) <= 0; play_W(2, 223) <= 0; play_W(2, 224) <= 0; play_W(2, 225) <= 0; play_W(2, 226) <= 0; play_W(2, 227) <= 0; play_W(2, 228) <= 0; play_W(2, 229) <= 0; play_W(2, 230) <= 0; play_W(2, 231) <= 1; play_W(2, 232) <= 1; play_W(2, 233) <= 1; play_W(2, 234) <= 1; play_W(2, 235) <= 1; play_W(2, 236) <= 1; play_W(2, 237) <= 0; play_W(2, 238) <= 0; play_W(2, 239) <= 0; play_W(2, 240) <= 0; play_W(2, 241) <= 0; play_W(2, 242) <= 0; play_W(2, 243) <= 1; play_W(2, 244) <= 1; play_W(2, 245) <= 1; play_W(2, 246) <= 1; play_W(2, 247) <= 1; play_W(2, 248) <= 1; play_W(2, 249) <= 1; play_W(2, 250) <= 1; play_W(2, 251) <= 1; play_W(2, 252) <= 1; play_W(2, 253) <= 1; play_W(2, 254) <= 1; play_W(2, 255) <= 1; play_W(2, 256) <= 1; play_W(2, 257) <= 1; play_W(2, 258) <= 1; play_W(2, 259) <= 1; play_W(2, 260) <= 1; play_W(2, 261) <= 0; play_W(2, 262) <= 0; play_W(2, 263) <= 0; play_W(2, 264) <= 0; play_W(2, 265) <= 0; play_W(2, 266) <= 0; play_W(2, 267) <= 0; play_W(2, 268) <= 0; play_W(2, 269) <= 0; 
play_W(3, 0) <= 0; play_W(3, 1) <= 0; play_W(3, 2) <= 0; play_W(3, 3) <= 1; play_W(3, 4) <= 1; play_W(3, 5) <= 1; play_W(3, 6) <= 1; play_W(3, 7) <= 1; play_W(3, 8) <= 1; play_W(3, 9) <= 0; play_W(3, 10) <= 0; play_W(3, 11) <= 0; play_W(3, 12) <= 0; play_W(3, 13) <= 0; play_W(3, 14) <= 0; play_W(3, 15) <= 1; play_W(3, 16) <= 1; play_W(3, 17) <= 1; play_W(3, 18) <= 1; play_W(3, 19) <= 1; play_W(3, 20) <= 1; play_W(3, 21) <= 0; play_W(3, 22) <= 0; play_W(3, 23) <= 0; play_W(3, 24) <= 0; play_W(3, 25) <= 0; play_W(3, 26) <= 0; play_W(3, 27) <= 0; play_W(3, 28) <= 0; play_W(3, 29) <= 0; play_W(3, 30) <= 1; play_W(3, 31) <= 1; play_W(3, 32) <= 1; play_W(3, 33) <= 1; play_W(3, 34) <= 1; play_W(3, 35) <= 1; play_W(3, 36) <= 0; play_W(3, 37) <= 0; play_W(3, 38) <= 0; play_W(3, 39) <= 0; play_W(3, 40) <= 0; play_W(3, 41) <= 0; play_W(3, 42) <= 0; play_W(3, 43) <= 0; play_W(3, 44) <= 0; play_W(3, 45) <= 0; play_W(3, 46) <= 0; play_W(3, 47) <= 0; play_W(3, 48) <= 0; play_W(3, 49) <= 0; play_W(3, 50) <= 0; play_W(3, 51) <= 0; play_W(3, 52) <= 0; play_W(3, 53) <= 0; play_W(3, 54) <= 0; play_W(3, 55) <= 0; play_W(3, 56) <= 0; play_W(3, 57) <= 0; play_W(3, 58) <= 0; play_W(3, 59) <= 0; play_W(3, 60) <= 1; play_W(3, 61) <= 1; play_W(3, 62) <= 1; play_W(3, 63) <= 1; play_W(3, 64) <= 1; play_W(3, 65) <= 1; play_W(3, 66) <= 1; play_W(3, 67) <= 1; play_W(3, 68) <= 1; play_W(3, 69) <= 0; play_W(3, 70) <= 0; play_W(3, 71) <= 0; play_W(3, 72) <= 0; play_W(3, 73) <= 0; play_W(3, 74) <= 0; play_W(3, 75) <= 0; play_W(3, 76) <= 0; play_W(3, 77) <= 0; play_W(3, 78) <= 0; play_W(3, 79) <= 0; play_W(3, 80) <= 0; play_W(3, 81) <= 1; play_W(3, 82) <= 1; play_W(3, 83) <= 1; play_W(3, 84) <= 1; play_W(3, 85) <= 1; play_W(3, 86) <= 1; play_W(3, 87) <= 0; play_W(3, 88) <= 0; play_W(3, 89) <= 0; play_W(3, 90) <= 0; play_W(3, 91) <= 0; play_W(3, 92) <= 0; play_W(3, 93) <= 0; play_W(3, 94) <= 0; play_W(3, 95) <= 0; play_W(3, 96) <= 0; play_W(3, 97) <= 0; play_W(3, 98) <= 0; play_W(3, 99) <= 1; play_W(3, 100) <= 1; play_W(3, 101) <= 1; play_W(3, 102) <= 1; play_W(3, 103) <= 1; play_W(3, 104) <= 1; play_W(3, 105) <= 0; play_W(3, 106) <= 0; play_W(3, 107) <= 0; play_W(3, 108) <= 0; play_W(3, 109) <= 0; play_W(3, 110) <= 0; play_W(3, 111) <= 0; play_W(3, 112) <= 0; play_W(3, 113) <= 0; play_W(3, 114) <= 0; play_W(3, 115) <= 0; play_W(3, 116) <= 0; play_W(3, 117) <= 0; play_W(3, 118) <= 0; play_W(3, 119) <= 0; play_W(3, 120) <= 0; play_W(3, 121) <= 0; play_W(3, 122) <= 0; play_W(3, 123) <= 0; play_W(3, 124) <= 0; play_W(3, 125) <= 0; play_W(3, 126) <= 0; play_W(3, 127) <= 0; play_W(3, 128) <= 0; play_W(3, 129) <= 0; play_W(3, 130) <= 0; play_W(3, 131) <= 0; play_W(3, 132) <= 0; play_W(3, 133) <= 0; play_W(3, 134) <= 0; play_W(3, 135) <= 0; play_W(3, 136) <= 0; play_W(3, 137) <= 0; play_W(3, 138) <= 0; play_W(3, 139) <= 0; play_W(3, 140) <= 0; play_W(3, 141) <= 0; play_W(3, 142) <= 0; play_W(3, 143) <= 0; play_W(3, 144) <= 0; play_W(3, 145) <= 0; play_W(3, 146) <= 0; play_W(3, 147) <= 0; play_W(3, 148) <= 0; play_W(3, 149) <= 0; play_W(3, 150) <= 0; play_W(3, 151) <= 0; play_W(3, 152) <= 0; play_W(3, 153) <= 0; play_W(3, 154) <= 0; play_W(3, 155) <= 0; play_W(3, 156) <= 0; play_W(3, 157) <= 0; play_W(3, 158) <= 0; play_W(3, 159) <= 0; play_W(3, 160) <= 0; play_W(3, 161) <= 0; play_W(3, 162) <= 0; play_W(3, 163) <= 0; play_W(3, 164) <= 0; play_W(3, 165) <= 1; play_W(3, 166) <= 1; play_W(3, 167) <= 1; play_W(3, 168) <= 1; play_W(3, 169) <= 1; play_W(3, 170) <= 1; play_W(3, 171) <= 0; play_W(3, 172) <= 0; play_W(3, 173) <= 0; play_W(3, 174) <= 0; play_W(3, 175) <= 0; play_W(3, 176) <= 0; play_W(3, 177) <= 1; play_W(3, 178) <= 1; play_W(3, 179) <= 1; play_W(3, 180) <= 1; play_W(3, 181) <= 1; play_W(3, 182) <= 1; play_W(3, 183) <= 0; play_W(3, 184) <= 0; play_W(3, 185) <= 0; play_W(3, 186) <= 0; play_W(3, 187) <= 0; play_W(3, 188) <= 0; play_W(3, 189) <= 1; play_W(3, 190) <= 1; play_W(3, 191) <= 1; play_W(3, 192) <= 1; play_W(3, 193) <= 1; play_W(3, 194) <= 1; play_W(3, 195) <= 0; play_W(3, 196) <= 0; play_W(3, 197) <= 0; play_W(3, 198) <= 1; play_W(3, 199) <= 1; play_W(3, 200) <= 1; play_W(3, 201) <= 1; play_W(3, 202) <= 1; play_W(3, 203) <= 1; play_W(3, 204) <= 0; play_W(3, 205) <= 0; play_W(3, 206) <= 0; play_W(3, 207) <= 1; play_W(3, 208) <= 1; play_W(3, 209) <= 1; play_W(3, 210) <= 1; play_W(3, 211) <= 1; play_W(3, 212) <= 1; play_W(3, 213) <= 0; play_W(3, 214) <= 0; play_W(3, 215) <= 0; play_W(3, 216) <= 1; play_W(3, 217) <= 1; play_W(3, 218) <= 1; play_W(3, 219) <= 1; play_W(3, 220) <= 1; play_W(3, 221) <= 1; play_W(3, 222) <= 1; play_W(3, 223) <= 1; play_W(3, 224) <= 1; play_W(3, 225) <= 0; play_W(3, 226) <= 0; play_W(3, 227) <= 0; play_W(3, 228) <= 0; play_W(3, 229) <= 0; play_W(3, 230) <= 0; play_W(3, 231) <= 1; play_W(3, 232) <= 1; play_W(3, 233) <= 1; play_W(3, 234) <= 1; play_W(3, 235) <= 1; play_W(3, 236) <= 1; play_W(3, 237) <= 0; play_W(3, 238) <= 0; play_W(3, 239) <= 0; play_W(3, 240) <= 0; play_W(3, 241) <= 0; play_W(3, 242) <= 0; play_W(3, 243) <= 0; play_W(3, 244) <= 0; play_W(3, 245) <= 0; play_W(3, 246) <= 1; play_W(3, 247) <= 1; play_W(3, 248) <= 1; play_W(3, 249) <= 1; play_W(3, 250) <= 1; play_W(3, 251) <= 1; play_W(3, 252) <= 0; play_W(3, 253) <= 0; play_W(3, 254) <= 0; play_W(3, 255) <= 0; play_W(3, 256) <= 0; play_W(3, 257) <= 0; play_W(3, 258) <= 1; play_W(3, 259) <= 1; play_W(3, 260) <= 1; play_W(3, 261) <= 1; play_W(3, 262) <= 1; play_W(3, 263) <= 1; play_W(3, 264) <= 0; play_W(3, 265) <= 0; play_W(3, 266) <= 0; play_W(3, 267) <= 0; play_W(3, 268) <= 0; play_W(3, 269) <= 0; 
play_W(4, 0) <= 0; play_W(4, 1) <= 0; play_W(4, 2) <= 0; play_W(4, 3) <= 1; play_W(4, 4) <= 1; play_W(4, 5) <= 1; play_W(4, 6) <= 1; play_W(4, 7) <= 1; play_W(4, 8) <= 1; play_W(4, 9) <= 0; play_W(4, 10) <= 0; play_W(4, 11) <= 0; play_W(4, 12) <= 0; play_W(4, 13) <= 0; play_W(4, 14) <= 0; play_W(4, 15) <= 1; play_W(4, 16) <= 1; play_W(4, 17) <= 1; play_W(4, 18) <= 1; play_W(4, 19) <= 1; play_W(4, 20) <= 1; play_W(4, 21) <= 0; play_W(4, 22) <= 0; play_W(4, 23) <= 0; play_W(4, 24) <= 0; play_W(4, 25) <= 0; play_W(4, 26) <= 0; play_W(4, 27) <= 0; play_W(4, 28) <= 0; play_W(4, 29) <= 0; play_W(4, 30) <= 1; play_W(4, 31) <= 1; play_W(4, 32) <= 1; play_W(4, 33) <= 1; play_W(4, 34) <= 1; play_W(4, 35) <= 1; play_W(4, 36) <= 0; play_W(4, 37) <= 0; play_W(4, 38) <= 0; play_W(4, 39) <= 0; play_W(4, 40) <= 0; play_W(4, 41) <= 0; play_W(4, 42) <= 0; play_W(4, 43) <= 0; play_W(4, 44) <= 0; play_W(4, 45) <= 0; play_W(4, 46) <= 0; play_W(4, 47) <= 0; play_W(4, 48) <= 0; play_W(4, 49) <= 0; play_W(4, 50) <= 0; play_W(4, 51) <= 0; play_W(4, 52) <= 0; play_W(4, 53) <= 0; play_W(4, 54) <= 0; play_W(4, 55) <= 0; play_W(4, 56) <= 0; play_W(4, 57) <= 0; play_W(4, 58) <= 0; play_W(4, 59) <= 0; play_W(4, 60) <= 1; play_W(4, 61) <= 1; play_W(4, 62) <= 1; play_W(4, 63) <= 1; play_W(4, 64) <= 1; play_W(4, 65) <= 1; play_W(4, 66) <= 1; play_W(4, 67) <= 1; play_W(4, 68) <= 1; play_W(4, 69) <= 0; play_W(4, 70) <= 0; play_W(4, 71) <= 0; play_W(4, 72) <= 0; play_W(4, 73) <= 0; play_W(4, 74) <= 0; play_W(4, 75) <= 0; play_W(4, 76) <= 0; play_W(4, 77) <= 0; play_W(4, 78) <= 0; play_W(4, 79) <= 0; play_W(4, 80) <= 0; play_W(4, 81) <= 1; play_W(4, 82) <= 1; play_W(4, 83) <= 1; play_W(4, 84) <= 1; play_W(4, 85) <= 1; play_W(4, 86) <= 1; play_W(4, 87) <= 0; play_W(4, 88) <= 0; play_W(4, 89) <= 0; play_W(4, 90) <= 0; play_W(4, 91) <= 0; play_W(4, 92) <= 0; play_W(4, 93) <= 0; play_W(4, 94) <= 0; play_W(4, 95) <= 0; play_W(4, 96) <= 0; play_W(4, 97) <= 0; play_W(4, 98) <= 0; play_W(4, 99) <= 1; play_W(4, 100) <= 1; play_W(4, 101) <= 1; play_W(4, 102) <= 1; play_W(4, 103) <= 1; play_W(4, 104) <= 1; play_W(4, 105) <= 0; play_W(4, 106) <= 0; play_W(4, 107) <= 0; play_W(4, 108) <= 0; play_W(4, 109) <= 0; play_W(4, 110) <= 0; play_W(4, 111) <= 0; play_W(4, 112) <= 0; play_W(4, 113) <= 0; play_W(4, 114) <= 0; play_W(4, 115) <= 0; play_W(4, 116) <= 0; play_W(4, 117) <= 0; play_W(4, 118) <= 0; play_W(4, 119) <= 0; play_W(4, 120) <= 0; play_W(4, 121) <= 0; play_W(4, 122) <= 0; play_W(4, 123) <= 0; play_W(4, 124) <= 0; play_W(4, 125) <= 0; play_W(4, 126) <= 0; play_W(4, 127) <= 0; play_W(4, 128) <= 0; play_W(4, 129) <= 0; play_W(4, 130) <= 0; play_W(4, 131) <= 0; play_W(4, 132) <= 0; play_W(4, 133) <= 0; play_W(4, 134) <= 0; play_W(4, 135) <= 0; play_W(4, 136) <= 0; play_W(4, 137) <= 0; play_W(4, 138) <= 0; play_W(4, 139) <= 0; play_W(4, 140) <= 0; play_W(4, 141) <= 0; play_W(4, 142) <= 0; play_W(4, 143) <= 0; play_W(4, 144) <= 0; play_W(4, 145) <= 0; play_W(4, 146) <= 0; play_W(4, 147) <= 0; play_W(4, 148) <= 0; play_W(4, 149) <= 0; play_W(4, 150) <= 0; play_W(4, 151) <= 0; play_W(4, 152) <= 0; play_W(4, 153) <= 0; play_W(4, 154) <= 0; play_W(4, 155) <= 0; play_W(4, 156) <= 0; play_W(4, 157) <= 0; play_W(4, 158) <= 0; play_W(4, 159) <= 0; play_W(4, 160) <= 0; play_W(4, 161) <= 0; play_W(4, 162) <= 0; play_W(4, 163) <= 0; play_W(4, 164) <= 0; play_W(4, 165) <= 1; play_W(4, 166) <= 1; play_W(4, 167) <= 1; play_W(4, 168) <= 1; play_W(4, 169) <= 1; play_W(4, 170) <= 1; play_W(4, 171) <= 0; play_W(4, 172) <= 0; play_W(4, 173) <= 0; play_W(4, 174) <= 0; play_W(4, 175) <= 0; play_W(4, 176) <= 0; play_W(4, 177) <= 1; play_W(4, 178) <= 1; play_W(4, 179) <= 1; play_W(4, 180) <= 1; play_W(4, 181) <= 1; play_W(4, 182) <= 1; play_W(4, 183) <= 0; play_W(4, 184) <= 0; play_W(4, 185) <= 0; play_W(4, 186) <= 0; play_W(4, 187) <= 0; play_W(4, 188) <= 0; play_W(4, 189) <= 1; play_W(4, 190) <= 1; play_W(4, 191) <= 1; play_W(4, 192) <= 1; play_W(4, 193) <= 1; play_W(4, 194) <= 1; play_W(4, 195) <= 0; play_W(4, 196) <= 0; play_W(4, 197) <= 0; play_W(4, 198) <= 1; play_W(4, 199) <= 1; play_W(4, 200) <= 1; play_W(4, 201) <= 1; play_W(4, 202) <= 1; play_W(4, 203) <= 1; play_W(4, 204) <= 0; play_W(4, 205) <= 0; play_W(4, 206) <= 0; play_W(4, 207) <= 1; play_W(4, 208) <= 1; play_W(4, 209) <= 1; play_W(4, 210) <= 1; play_W(4, 211) <= 1; play_W(4, 212) <= 1; play_W(4, 213) <= 0; play_W(4, 214) <= 0; play_W(4, 215) <= 0; play_W(4, 216) <= 1; play_W(4, 217) <= 1; play_W(4, 218) <= 1; play_W(4, 219) <= 1; play_W(4, 220) <= 1; play_W(4, 221) <= 1; play_W(4, 222) <= 1; play_W(4, 223) <= 1; play_W(4, 224) <= 1; play_W(4, 225) <= 0; play_W(4, 226) <= 0; play_W(4, 227) <= 0; play_W(4, 228) <= 0; play_W(4, 229) <= 0; play_W(4, 230) <= 0; play_W(4, 231) <= 1; play_W(4, 232) <= 1; play_W(4, 233) <= 1; play_W(4, 234) <= 1; play_W(4, 235) <= 1; play_W(4, 236) <= 1; play_W(4, 237) <= 0; play_W(4, 238) <= 0; play_W(4, 239) <= 0; play_W(4, 240) <= 0; play_W(4, 241) <= 0; play_W(4, 242) <= 0; play_W(4, 243) <= 0; play_W(4, 244) <= 0; play_W(4, 245) <= 0; play_W(4, 246) <= 1; play_W(4, 247) <= 1; play_W(4, 248) <= 1; play_W(4, 249) <= 1; play_W(4, 250) <= 1; play_W(4, 251) <= 1; play_W(4, 252) <= 0; play_W(4, 253) <= 0; play_W(4, 254) <= 0; play_W(4, 255) <= 0; play_W(4, 256) <= 0; play_W(4, 257) <= 0; play_W(4, 258) <= 1; play_W(4, 259) <= 1; play_W(4, 260) <= 1; play_W(4, 261) <= 1; play_W(4, 262) <= 1; play_W(4, 263) <= 1; play_W(4, 264) <= 0; play_W(4, 265) <= 0; play_W(4, 266) <= 0; play_W(4, 267) <= 0; play_W(4, 268) <= 0; play_W(4, 269) <= 0; 
play_W(5, 0) <= 0; play_W(5, 1) <= 0; play_W(5, 2) <= 0; play_W(5, 3) <= 1; play_W(5, 4) <= 1; play_W(5, 5) <= 1; play_W(5, 6) <= 1; play_W(5, 7) <= 1; play_W(5, 8) <= 1; play_W(5, 9) <= 0; play_W(5, 10) <= 0; play_W(5, 11) <= 0; play_W(5, 12) <= 0; play_W(5, 13) <= 0; play_W(5, 14) <= 0; play_W(5, 15) <= 1; play_W(5, 16) <= 1; play_W(5, 17) <= 1; play_W(5, 18) <= 1; play_W(5, 19) <= 1; play_W(5, 20) <= 1; play_W(5, 21) <= 0; play_W(5, 22) <= 0; play_W(5, 23) <= 0; play_W(5, 24) <= 0; play_W(5, 25) <= 0; play_W(5, 26) <= 0; play_W(5, 27) <= 0; play_W(5, 28) <= 0; play_W(5, 29) <= 0; play_W(5, 30) <= 1; play_W(5, 31) <= 1; play_W(5, 32) <= 1; play_W(5, 33) <= 1; play_W(5, 34) <= 1; play_W(5, 35) <= 1; play_W(5, 36) <= 0; play_W(5, 37) <= 0; play_W(5, 38) <= 0; play_W(5, 39) <= 0; play_W(5, 40) <= 0; play_W(5, 41) <= 0; play_W(5, 42) <= 0; play_W(5, 43) <= 0; play_W(5, 44) <= 0; play_W(5, 45) <= 0; play_W(5, 46) <= 0; play_W(5, 47) <= 0; play_W(5, 48) <= 0; play_W(5, 49) <= 0; play_W(5, 50) <= 0; play_W(5, 51) <= 0; play_W(5, 52) <= 0; play_W(5, 53) <= 0; play_W(5, 54) <= 0; play_W(5, 55) <= 0; play_W(5, 56) <= 0; play_W(5, 57) <= 0; play_W(5, 58) <= 0; play_W(5, 59) <= 0; play_W(5, 60) <= 1; play_W(5, 61) <= 1; play_W(5, 62) <= 1; play_W(5, 63) <= 1; play_W(5, 64) <= 1; play_W(5, 65) <= 1; play_W(5, 66) <= 1; play_W(5, 67) <= 1; play_W(5, 68) <= 1; play_W(5, 69) <= 0; play_W(5, 70) <= 0; play_W(5, 71) <= 0; play_W(5, 72) <= 0; play_W(5, 73) <= 0; play_W(5, 74) <= 0; play_W(5, 75) <= 0; play_W(5, 76) <= 0; play_W(5, 77) <= 0; play_W(5, 78) <= 0; play_W(5, 79) <= 0; play_W(5, 80) <= 0; play_W(5, 81) <= 1; play_W(5, 82) <= 1; play_W(5, 83) <= 1; play_W(5, 84) <= 1; play_W(5, 85) <= 1; play_W(5, 86) <= 1; play_W(5, 87) <= 0; play_W(5, 88) <= 0; play_W(5, 89) <= 0; play_W(5, 90) <= 0; play_W(5, 91) <= 0; play_W(5, 92) <= 0; play_W(5, 93) <= 0; play_W(5, 94) <= 0; play_W(5, 95) <= 0; play_W(5, 96) <= 0; play_W(5, 97) <= 0; play_W(5, 98) <= 0; play_W(5, 99) <= 1; play_W(5, 100) <= 1; play_W(5, 101) <= 1; play_W(5, 102) <= 1; play_W(5, 103) <= 1; play_W(5, 104) <= 1; play_W(5, 105) <= 0; play_W(5, 106) <= 0; play_W(5, 107) <= 0; play_W(5, 108) <= 0; play_W(5, 109) <= 0; play_W(5, 110) <= 0; play_W(5, 111) <= 0; play_W(5, 112) <= 0; play_W(5, 113) <= 0; play_W(5, 114) <= 0; play_W(5, 115) <= 0; play_W(5, 116) <= 0; play_W(5, 117) <= 0; play_W(5, 118) <= 0; play_W(5, 119) <= 0; play_W(5, 120) <= 0; play_W(5, 121) <= 0; play_W(5, 122) <= 0; play_W(5, 123) <= 0; play_W(5, 124) <= 0; play_W(5, 125) <= 0; play_W(5, 126) <= 0; play_W(5, 127) <= 0; play_W(5, 128) <= 0; play_W(5, 129) <= 0; play_W(5, 130) <= 0; play_W(5, 131) <= 0; play_W(5, 132) <= 0; play_W(5, 133) <= 0; play_W(5, 134) <= 0; play_W(5, 135) <= 0; play_W(5, 136) <= 0; play_W(5, 137) <= 0; play_W(5, 138) <= 0; play_W(5, 139) <= 0; play_W(5, 140) <= 0; play_W(5, 141) <= 0; play_W(5, 142) <= 0; play_W(5, 143) <= 0; play_W(5, 144) <= 0; play_W(5, 145) <= 0; play_W(5, 146) <= 0; play_W(5, 147) <= 0; play_W(5, 148) <= 0; play_W(5, 149) <= 0; play_W(5, 150) <= 0; play_W(5, 151) <= 0; play_W(5, 152) <= 0; play_W(5, 153) <= 0; play_W(5, 154) <= 0; play_W(5, 155) <= 0; play_W(5, 156) <= 0; play_W(5, 157) <= 0; play_W(5, 158) <= 0; play_W(5, 159) <= 0; play_W(5, 160) <= 0; play_W(5, 161) <= 0; play_W(5, 162) <= 0; play_W(5, 163) <= 0; play_W(5, 164) <= 0; play_W(5, 165) <= 1; play_W(5, 166) <= 1; play_W(5, 167) <= 1; play_W(5, 168) <= 1; play_W(5, 169) <= 1; play_W(5, 170) <= 1; play_W(5, 171) <= 0; play_W(5, 172) <= 0; play_W(5, 173) <= 0; play_W(5, 174) <= 0; play_W(5, 175) <= 0; play_W(5, 176) <= 0; play_W(5, 177) <= 1; play_W(5, 178) <= 1; play_W(5, 179) <= 1; play_W(5, 180) <= 1; play_W(5, 181) <= 1; play_W(5, 182) <= 1; play_W(5, 183) <= 0; play_W(5, 184) <= 0; play_W(5, 185) <= 0; play_W(5, 186) <= 0; play_W(5, 187) <= 0; play_W(5, 188) <= 0; play_W(5, 189) <= 1; play_W(5, 190) <= 1; play_W(5, 191) <= 1; play_W(5, 192) <= 1; play_W(5, 193) <= 1; play_W(5, 194) <= 1; play_W(5, 195) <= 0; play_W(5, 196) <= 0; play_W(5, 197) <= 0; play_W(5, 198) <= 1; play_W(5, 199) <= 1; play_W(5, 200) <= 1; play_W(5, 201) <= 1; play_W(5, 202) <= 1; play_W(5, 203) <= 1; play_W(5, 204) <= 0; play_W(5, 205) <= 0; play_W(5, 206) <= 0; play_W(5, 207) <= 1; play_W(5, 208) <= 1; play_W(5, 209) <= 1; play_W(5, 210) <= 1; play_W(5, 211) <= 1; play_W(5, 212) <= 1; play_W(5, 213) <= 0; play_W(5, 214) <= 0; play_W(5, 215) <= 0; play_W(5, 216) <= 1; play_W(5, 217) <= 1; play_W(5, 218) <= 1; play_W(5, 219) <= 1; play_W(5, 220) <= 1; play_W(5, 221) <= 1; play_W(5, 222) <= 1; play_W(5, 223) <= 1; play_W(5, 224) <= 1; play_W(5, 225) <= 0; play_W(5, 226) <= 0; play_W(5, 227) <= 0; play_W(5, 228) <= 0; play_W(5, 229) <= 0; play_W(5, 230) <= 0; play_W(5, 231) <= 1; play_W(5, 232) <= 1; play_W(5, 233) <= 1; play_W(5, 234) <= 1; play_W(5, 235) <= 1; play_W(5, 236) <= 1; play_W(5, 237) <= 0; play_W(5, 238) <= 0; play_W(5, 239) <= 0; play_W(5, 240) <= 0; play_W(5, 241) <= 0; play_W(5, 242) <= 0; play_W(5, 243) <= 0; play_W(5, 244) <= 0; play_W(5, 245) <= 0; play_W(5, 246) <= 1; play_W(5, 247) <= 1; play_W(5, 248) <= 1; play_W(5, 249) <= 1; play_W(5, 250) <= 1; play_W(5, 251) <= 1; play_W(5, 252) <= 0; play_W(5, 253) <= 0; play_W(5, 254) <= 0; play_W(5, 255) <= 0; play_W(5, 256) <= 0; play_W(5, 257) <= 0; play_W(5, 258) <= 1; play_W(5, 259) <= 1; play_W(5, 260) <= 1; play_W(5, 261) <= 1; play_W(5, 262) <= 1; play_W(5, 263) <= 1; play_W(5, 264) <= 0; play_W(5, 265) <= 0; play_W(5, 266) <= 0; play_W(5, 267) <= 0; play_W(5, 268) <= 0; play_W(5, 269) <= 0; 
play_W(6, 0) <= 0; play_W(6, 1) <= 0; play_W(6, 2) <= 0; play_W(6, 3) <= 1; play_W(6, 4) <= 1; play_W(6, 5) <= 1; play_W(6, 6) <= 1; play_W(6, 7) <= 1; play_W(6, 8) <= 1; play_W(6, 9) <= 0; play_W(6, 10) <= 0; play_W(6, 11) <= 0; play_W(6, 12) <= 0; play_W(6, 13) <= 0; play_W(6, 14) <= 0; play_W(6, 15) <= 1; play_W(6, 16) <= 1; play_W(6, 17) <= 1; play_W(6, 18) <= 1; play_W(6, 19) <= 1; play_W(6, 20) <= 1; play_W(6, 21) <= 0; play_W(6, 22) <= 0; play_W(6, 23) <= 0; play_W(6, 24) <= 0; play_W(6, 25) <= 0; play_W(6, 26) <= 0; play_W(6, 27) <= 0; play_W(6, 28) <= 0; play_W(6, 29) <= 0; play_W(6, 30) <= 1; play_W(6, 31) <= 1; play_W(6, 32) <= 1; play_W(6, 33) <= 1; play_W(6, 34) <= 1; play_W(6, 35) <= 1; play_W(6, 36) <= 0; play_W(6, 37) <= 0; play_W(6, 38) <= 0; play_W(6, 39) <= 0; play_W(6, 40) <= 0; play_W(6, 41) <= 0; play_W(6, 42) <= 0; play_W(6, 43) <= 0; play_W(6, 44) <= 0; play_W(6, 45) <= 0; play_W(6, 46) <= 0; play_W(6, 47) <= 0; play_W(6, 48) <= 0; play_W(6, 49) <= 0; play_W(6, 50) <= 0; play_W(6, 51) <= 0; play_W(6, 52) <= 0; play_W(6, 53) <= 0; play_W(6, 54) <= 0; play_W(6, 55) <= 0; play_W(6, 56) <= 0; play_W(6, 57) <= 1; play_W(6, 58) <= 1; play_W(6, 59) <= 1; play_W(6, 60) <= 1; play_W(6, 61) <= 1; play_W(6, 62) <= 1; play_W(6, 63) <= 0; play_W(6, 64) <= 0; play_W(6, 65) <= 0; play_W(6, 66) <= 1; play_W(6, 67) <= 1; play_W(6, 68) <= 1; play_W(6, 69) <= 1; play_W(6, 70) <= 1; play_W(6, 71) <= 1; play_W(6, 72) <= 0; play_W(6, 73) <= 0; play_W(6, 74) <= 0; play_W(6, 75) <= 0; play_W(6, 76) <= 0; play_W(6, 77) <= 0; play_W(6, 78) <= 0; play_W(6, 79) <= 0; play_W(6, 80) <= 0; play_W(6, 81) <= 1; play_W(6, 82) <= 1; play_W(6, 83) <= 1; play_W(6, 84) <= 1; play_W(6, 85) <= 1; play_W(6, 86) <= 1; play_W(6, 87) <= 0; play_W(6, 88) <= 0; play_W(6, 89) <= 0; play_W(6, 90) <= 0; play_W(6, 91) <= 0; play_W(6, 92) <= 0; play_W(6, 93) <= 0; play_W(6, 94) <= 0; play_W(6, 95) <= 0; play_W(6, 96) <= 0; play_W(6, 97) <= 0; play_W(6, 98) <= 0; play_W(6, 99) <= 1; play_W(6, 100) <= 1; play_W(6, 101) <= 1; play_W(6, 102) <= 1; play_W(6, 103) <= 1; play_W(6, 104) <= 1; play_W(6, 105) <= 0; play_W(6, 106) <= 0; play_W(6, 107) <= 0; play_W(6, 108) <= 0; play_W(6, 109) <= 0; play_W(6, 110) <= 0; play_W(6, 111) <= 0; play_W(6, 112) <= 0; play_W(6, 113) <= 0; play_W(6, 114) <= 0; play_W(6, 115) <= 0; play_W(6, 116) <= 0; play_W(6, 117) <= 1; play_W(6, 118) <= 1; play_W(6, 119) <= 1; play_W(6, 120) <= 1; play_W(6, 121) <= 1; play_W(6, 122) <= 1; play_W(6, 123) <= 0; play_W(6, 124) <= 0; play_W(6, 125) <= 0; play_W(6, 126) <= 0; play_W(6, 127) <= 0; play_W(6, 128) <= 0; play_W(6, 129) <= 0; play_W(6, 130) <= 0; play_W(6, 131) <= 0; play_W(6, 132) <= 0; play_W(6, 133) <= 0; play_W(6, 134) <= 0; play_W(6, 135) <= 0; play_W(6, 136) <= 0; play_W(6, 137) <= 0; play_W(6, 138) <= 0; play_W(6, 139) <= 0; play_W(6, 140) <= 0; play_W(6, 141) <= 0; play_W(6, 142) <= 0; play_W(6, 143) <= 0; play_W(6, 144) <= 0; play_W(6, 145) <= 0; play_W(6, 146) <= 0; play_W(6, 147) <= 0; play_W(6, 148) <= 0; play_W(6, 149) <= 0; play_W(6, 150) <= 0; play_W(6, 151) <= 0; play_W(6, 152) <= 0; play_W(6, 153) <= 0; play_W(6, 154) <= 0; play_W(6, 155) <= 0; play_W(6, 156) <= 0; play_W(6, 157) <= 0; play_W(6, 158) <= 0; play_W(6, 159) <= 0; play_W(6, 160) <= 0; play_W(6, 161) <= 0; play_W(6, 162) <= 0; play_W(6, 163) <= 0; play_W(6, 164) <= 0; play_W(6, 165) <= 1; play_W(6, 166) <= 1; play_W(6, 167) <= 1; play_W(6, 168) <= 1; play_W(6, 169) <= 1; play_W(6, 170) <= 1; play_W(6, 171) <= 0; play_W(6, 172) <= 0; play_W(6, 173) <= 0; play_W(6, 174) <= 0; play_W(6, 175) <= 0; play_W(6, 176) <= 0; play_W(6, 177) <= 1; play_W(6, 178) <= 1; play_W(6, 179) <= 1; play_W(6, 180) <= 1; play_W(6, 181) <= 1; play_W(6, 182) <= 1; play_W(6, 183) <= 0; play_W(6, 184) <= 0; play_W(6, 185) <= 0; play_W(6, 186) <= 0; play_W(6, 187) <= 0; play_W(6, 188) <= 0; play_W(6, 189) <= 1; play_W(6, 190) <= 1; play_W(6, 191) <= 1; play_W(6, 192) <= 0; play_W(6, 193) <= 0; play_W(6, 194) <= 0; play_W(6, 195) <= 0; play_W(6, 196) <= 0; play_W(6, 197) <= 0; play_W(6, 198) <= 1; play_W(6, 199) <= 1; play_W(6, 200) <= 1; play_W(6, 201) <= 1; play_W(6, 202) <= 1; play_W(6, 203) <= 1; play_W(6, 204) <= 0; play_W(6, 205) <= 0; play_W(6, 206) <= 0; play_W(6, 207) <= 0; play_W(6, 208) <= 0; play_W(6, 209) <= 0; play_W(6, 210) <= 1; play_W(6, 211) <= 1; play_W(6, 212) <= 1; play_W(6, 213) <= 0; play_W(6, 214) <= 0; play_W(6, 215) <= 0; play_W(6, 216) <= 1; play_W(6, 217) <= 1; play_W(6, 218) <= 1; play_W(6, 219) <= 1; play_W(6, 220) <= 1; play_W(6, 221) <= 1; play_W(6, 222) <= 1; play_W(6, 223) <= 1; play_W(6, 224) <= 1; play_W(6, 225) <= 1; play_W(6, 226) <= 1; play_W(6, 227) <= 1; play_W(6, 228) <= 0; play_W(6, 229) <= 0; play_W(6, 230) <= 0; play_W(6, 231) <= 1; play_W(6, 232) <= 1; play_W(6, 233) <= 1; play_W(6, 234) <= 1; play_W(6, 235) <= 1; play_W(6, 236) <= 1; play_W(6, 237) <= 0; play_W(6, 238) <= 0; play_W(6, 239) <= 0; play_W(6, 240) <= 0; play_W(6, 241) <= 0; play_W(6, 242) <= 0; play_W(6, 243) <= 0; play_W(6, 244) <= 0; play_W(6, 245) <= 0; play_W(6, 246) <= 1; play_W(6, 247) <= 1; play_W(6, 248) <= 1; play_W(6, 249) <= 1; play_W(6, 250) <= 1; play_W(6, 251) <= 1; play_W(6, 252) <= 0; play_W(6, 253) <= 0; play_W(6, 254) <= 0; play_W(6, 255) <= 0; play_W(6, 256) <= 0; play_W(6, 257) <= 0; play_W(6, 258) <= 1; play_W(6, 259) <= 1; play_W(6, 260) <= 1; play_W(6, 261) <= 1; play_W(6, 262) <= 1; play_W(6, 263) <= 1; play_W(6, 264) <= 0; play_W(6, 265) <= 0; play_W(6, 266) <= 0; play_W(6, 267) <= 0; play_W(6, 268) <= 0; play_W(6, 269) <= 0; 
play_W(7, 0) <= 0; play_W(7, 1) <= 0; play_W(7, 2) <= 0; play_W(7, 3) <= 1; play_W(7, 4) <= 1; play_W(7, 5) <= 1; play_W(7, 6) <= 1; play_W(7, 7) <= 1; play_W(7, 8) <= 1; play_W(7, 9) <= 0; play_W(7, 10) <= 0; play_W(7, 11) <= 0; play_W(7, 12) <= 0; play_W(7, 13) <= 0; play_W(7, 14) <= 0; play_W(7, 15) <= 1; play_W(7, 16) <= 1; play_W(7, 17) <= 1; play_W(7, 18) <= 1; play_W(7, 19) <= 1; play_W(7, 20) <= 1; play_W(7, 21) <= 0; play_W(7, 22) <= 0; play_W(7, 23) <= 0; play_W(7, 24) <= 0; play_W(7, 25) <= 0; play_W(7, 26) <= 0; play_W(7, 27) <= 0; play_W(7, 28) <= 0; play_W(7, 29) <= 0; play_W(7, 30) <= 1; play_W(7, 31) <= 1; play_W(7, 32) <= 1; play_W(7, 33) <= 1; play_W(7, 34) <= 1; play_W(7, 35) <= 1; play_W(7, 36) <= 0; play_W(7, 37) <= 0; play_W(7, 38) <= 0; play_W(7, 39) <= 0; play_W(7, 40) <= 0; play_W(7, 41) <= 0; play_W(7, 42) <= 0; play_W(7, 43) <= 0; play_W(7, 44) <= 0; play_W(7, 45) <= 0; play_W(7, 46) <= 0; play_W(7, 47) <= 0; play_W(7, 48) <= 0; play_W(7, 49) <= 0; play_W(7, 50) <= 0; play_W(7, 51) <= 0; play_W(7, 52) <= 0; play_W(7, 53) <= 0; play_W(7, 54) <= 0; play_W(7, 55) <= 0; play_W(7, 56) <= 0; play_W(7, 57) <= 1; play_W(7, 58) <= 1; play_W(7, 59) <= 1; play_W(7, 60) <= 1; play_W(7, 61) <= 1; play_W(7, 62) <= 1; play_W(7, 63) <= 0; play_W(7, 64) <= 0; play_W(7, 65) <= 0; play_W(7, 66) <= 1; play_W(7, 67) <= 1; play_W(7, 68) <= 1; play_W(7, 69) <= 1; play_W(7, 70) <= 1; play_W(7, 71) <= 1; play_W(7, 72) <= 0; play_W(7, 73) <= 0; play_W(7, 74) <= 0; play_W(7, 75) <= 0; play_W(7, 76) <= 0; play_W(7, 77) <= 0; play_W(7, 78) <= 0; play_W(7, 79) <= 0; play_W(7, 80) <= 0; play_W(7, 81) <= 1; play_W(7, 82) <= 1; play_W(7, 83) <= 1; play_W(7, 84) <= 1; play_W(7, 85) <= 1; play_W(7, 86) <= 1; play_W(7, 87) <= 0; play_W(7, 88) <= 0; play_W(7, 89) <= 0; play_W(7, 90) <= 0; play_W(7, 91) <= 0; play_W(7, 92) <= 0; play_W(7, 93) <= 0; play_W(7, 94) <= 0; play_W(7, 95) <= 0; play_W(7, 96) <= 0; play_W(7, 97) <= 0; play_W(7, 98) <= 0; play_W(7, 99) <= 1; play_W(7, 100) <= 1; play_W(7, 101) <= 1; play_W(7, 102) <= 1; play_W(7, 103) <= 1; play_W(7, 104) <= 1; play_W(7, 105) <= 0; play_W(7, 106) <= 0; play_W(7, 107) <= 0; play_W(7, 108) <= 0; play_W(7, 109) <= 0; play_W(7, 110) <= 0; play_W(7, 111) <= 0; play_W(7, 112) <= 0; play_W(7, 113) <= 0; play_W(7, 114) <= 0; play_W(7, 115) <= 0; play_W(7, 116) <= 0; play_W(7, 117) <= 1; play_W(7, 118) <= 1; play_W(7, 119) <= 1; play_W(7, 120) <= 1; play_W(7, 121) <= 1; play_W(7, 122) <= 1; play_W(7, 123) <= 0; play_W(7, 124) <= 0; play_W(7, 125) <= 0; play_W(7, 126) <= 0; play_W(7, 127) <= 0; play_W(7, 128) <= 0; play_W(7, 129) <= 0; play_W(7, 130) <= 0; play_W(7, 131) <= 0; play_W(7, 132) <= 0; play_W(7, 133) <= 0; play_W(7, 134) <= 0; play_W(7, 135) <= 0; play_W(7, 136) <= 0; play_W(7, 137) <= 0; play_W(7, 138) <= 0; play_W(7, 139) <= 0; play_W(7, 140) <= 0; play_W(7, 141) <= 0; play_W(7, 142) <= 0; play_W(7, 143) <= 0; play_W(7, 144) <= 0; play_W(7, 145) <= 0; play_W(7, 146) <= 0; play_W(7, 147) <= 0; play_W(7, 148) <= 0; play_W(7, 149) <= 0; play_W(7, 150) <= 0; play_W(7, 151) <= 0; play_W(7, 152) <= 0; play_W(7, 153) <= 0; play_W(7, 154) <= 0; play_W(7, 155) <= 0; play_W(7, 156) <= 0; play_W(7, 157) <= 0; play_W(7, 158) <= 0; play_W(7, 159) <= 0; play_W(7, 160) <= 0; play_W(7, 161) <= 0; play_W(7, 162) <= 0; play_W(7, 163) <= 0; play_W(7, 164) <= 0; play_W(7, 165) <= 1; play_W(7, 166) <= 1; play_W(7, 167) <= 1; play_W(7, 168) <= 1; play_W(7, 169) <= 1; play_W(7, 170) <= 1; play_W(7, 171) <= 0; play_W(7, 172) <= 0; play_W(7, 173) <= 0; play_W(7, 174) <= 0; play_W(7, 175) <= 0; play_W(7, 176) <= 0; play_W(7, 177) <= 1; play_W(7, 178) <= 1; play_W(7, 179) <= 1; play_W(7, 180) <= 1; play_W(7, 181) <= 1; play_W(7, 182) <= 1; play_W(7, 183) <= 0; play_W(7, 184) <= 0; play_W(7, 185) <= 0; play_W(7, 186) <= 0; play_W(7, 187) <= 0; play_W(7, 188) <= 0; play_W(7, 189) <= 1; play_W(7, 190) <= 1; play_W(7, 191) <= 1; play_W(7, 192) <= 0; play_W(7, 193) <= 0; play_W(7, 194) <= 0; play_W(7, 195) <= 0; play_W(7, 196) <= 0; play_W(7, 197) <= 0; play_W(7, 198) <= 1; play_W(7, 199) <= 1; play_W(7, 200) <= 1; play_W(7, 201) <= 1; play_W(7, 202) <= 1; play_W(7, 203) <= 1; play_W(7, 204) <= 0; play_W(7, 205) <= 0; play_W(7, 206) <= 0; play_W(7, 207) <= 0; play_W(7, 208) <= 0; play_W(7, 209) <= 0; play_W(7, 210) <= 1; play_W(7, 211) <= 1; play_W(7, 212) <= 1; play_W(7, 213) <= 0; play_W(7, 214) <= 0; play_W(7, 215) <= 0; play_W(7, 216) <= 1; play_W(7, 217) <= 1; play_W(7, 218) <= 1; play_W(7, 219) <= 1; play_W(7, 220) <= 1; play_W(7, 221) <= 1; play_W(7, 222) <= 1; play_W(7, 223) <= 1; play_W(7, 224) <= 1; play_W(7, 225) <= 1; play_W(7, 226) <= 1; play_W(7, 227) <= 1; play_W(7, 228) <= 0; play_W(7, 229) <= 0; play_W(7, 230) <= 0; play_W(7, 231) <= 1; play_W(7, 232) <= 1; play_W(7, 233) <= 1; play_W(7, 234) <= 1; play_W(7, 235) <= 1; play_W(7, 236) <= 1; play_W(7, 237) <= 0; play_W(7, 238) <= 0; play_W(7, 239) <= 0; play_W(7, 240) <= 0; play_W(7, 241) <= 0; play_W(7, 242) <= 0; play_W(7, 243) <= 0; play_W(7, 244) <= 0; play_W(7, 245) <= 0; play_W(7, 246) <= 1; play_W(7, 247) <= 1; play_W(7, 248) <= 1; play_W(7, 249) <= 1; play_W(7, 250) <= 1; play_W(7, 251) <= 1; play_W(7, 252) <= 0; play_W(7, 253) <= 0; play_W(7, 254) <= 0; play_W(7, 255) <= 0; play_W(7, 256) <= 0; play_W(7, 257) <= 0; play_W(7, 258) <= 1; play_W(7, 259) <= 1; play_W(7, 260) <= 1; play_W(7, 261) <= 1; play_W(7, 262) <= 1; play_W(7, 263) <= 1; play_W(7, 264) <= 0; play_W(7, 265) <= 0; play_W(7, 266) <= 0; play_W(7, 267) <= 0; play_W(7, 268) <= 0; play_W(7, 269) <= 0; 
play_W(8, 0) <= 0; play_W(8, 1) <= 0; play_W(8, 2) <= 0; play_W(8, 3) <= 1; play_W(8, 4) <= 1; play_W(8, 5) <= 1; play_W(8, 6) <= 1; play_W(8, 7) <= 1; play_W(8, 8) <= 1; play_W(8, 9) <= 0; play_W(8, 10) <= 0; play_W(8, 11) <= 0; play_W(8, 12) <= 0; play_W(8, 13) <= 0; play_W(8, 14) <= 0; play_W(8, 15) <= 1; play_W(8, 16) <= 1; play_W(8, 17) <= 1; play_W(8, 18) <= 1; play_W(8, 19) <= 1; play_W(8, 20) <= 1; play_W(8, 21) <= 0; play_W(8, 22) <= 0; play_W(8, 23) <= 0; play_W(8, 24) <= 0; play_W(8, 25) <= 0; play_W(8, 26) <= 0; play_W(8, 27) <= 0; play_W(8, 28) <= 0; play_W(8, 29) <= 0; play_W(8, 30) <= 1; play_W(8, 31) <= 1; play_W(8, 32) <= 1; play_W(8, 33) <= 1; play_W(8, 34) <= 1; play_W(8, 35) <= 1; play_W(8, 36) <= 0; play_W(8, 37) <= 0; play_W(8, 38) <= 0; play_W(8, 39) <= 0; play_W(8, 40) <= 0; play_W(8, 41) <= 0; play_W(8, 42) <= 0; play_W(8, 43) <= 0; play_W(8, 44) <= 0; play_W(8, 45) <= 0; play_W(8, 46) <= 0; play_W(8, 47) <= 0; play_W(8, 48) <= 0; play_W(8, 49) <= 0; play_W(8, 50) <= 0; play_W(8, 51) <= 0; play_W(8, 52) <= 0; play_W(8, 53) <= 0; play_W(8, 54) <= 0; play_W(8, 55) <= 0; play_W(8, 56) <= 0; play_W(8, 57) <= 1; play_W(8, 58) <= 1; play_W(8, 59) <= 1; play_W(8, 60) <= 1; play_W(8, 61) <= 1; play_W(8, 62) <= 1; play_W(8, 63) <= 0; play_W(8, 64) <= 0; play_W(8, 65) <= 0; play_W(8, 66) <= 1; play_W(8, 67) <= 1; play_W(8, 68) <= 1; play_W(8, 69) <= 1; play_W(8, 70) <= 1; play_W(8, 71) <= 1; play_W(8, 72) <= 0; play_W(8, 73) <= 0; play_W(8, 74) <= 0; play_W(8, 75) <= 0; play_W(8, 76) <= 0; play_W(8, 77) <= 0; play_W(8, 78) <= 0; play_W(8, 79) <= 0; play_W(8, 80) <= 0; play_W(8, 81) <= 1; play_W(8, 82) <= 1; play_W(8, 83) <= 1; play_W(8, 84) <= 1; play_W(8, 85) <= 1; play_W(8, 86) <= 1; play_W(8, 87) <= 0; play_W(8, 88) <= 0; play_W(8, 89) <= 0; play_W(8, 90) <= 0; play_W(8, 91) <= 0; play_W(8, 92) <= 0; play_W(8, 93) <= 0; play_W(8, 94) <= 0; play_W(8, 95) <= 0; play_W(8, 96) <= 0; play_W(8, 97) <= 0; play_W(8, 98) <= 0; play_W(8, 99) <= 1; play_W(8, 100) <= 1; play_W(8, 101) <= 1; play_W(8, 102) <= 1; play_W(8, 103) <= 1; play_W(8, 104) <= 1; play_W(8, 105) <= 0; play_W(8, 106) <= 0; play_W(8, 107) <= 0; play_W(8, 108) <= 0; play_W(8, 109) <= 0; play_W(8, 110) <= 0; play_W(8, 111) <= 0; play_W(8, 112) <= 0; play_W(8, 113) <= 0; play_W(8, 114) <= 0; play_W(8, 115) <= 0; play_W(8, 116) <= 0; play_W(8, 117) <= 1; play_W(8, 118) <= 1; play_W(8, 119) <= 1; play_W(8, 120) <= 1; play_W(8, 121) <= 1; play_W(8, 122) <= 1; play_W(8, 123) <= 0; play_W(8, 124) <= 0; play_W(8, 125) <= 0; play_W(8, 126) <= 0; play_W(8, 127) <= 0; play_W(8, 128) <= 0; play_W(8, 129) <= 0; play_W(8, 130) <= 0; play_W(8, 131) <= 0; play_W(8, 132) <= 0; play_W(8, 133) <= 0; play_W(8, 134) <= 0; play_W(8, 135) <= 0; play_W(8, 136) <= 0; play_W(8, 137) <= 0; play_W(8, 138) <= 0; play_W(8, 139) <= 0; play_W(8, 140) <= 0; play_W(8, 141) <= 0; play_W(8, 142) <= 0; play_W(8, 143) <= 0; play_W(8, 144) <= 0; play_W(8, 145) <= 0; play_W(8, 146) <= 0; play_W(8, 147) <= 0; play_W(8, 148) <= 0; play_W(8, 149) <= 0; play_W(8, 150) <= 0; play_W(8, 151) <= 0; play_W(8, 152) <= 0; play_W(8, 153) <= 0; play_W(8, 154) <= 0; play_W(8, 155) <= 0; play_W(8, 156) <= 0; play_W(8, 157) <= 0; play_W(8, 158) <= 0; play_W(8, 159) <= 0; play_W(8, 160) <= 0; play_W(8, 161) <= 0; play_W(8, 162) <= 0; play_W(8, 163) <= 0; play_W(8, 164) <= 0; play_W(8, 165) <= 1; play_W(8, 166) <= 1; play_W(8, 167) <= 1; play_W(8, 168) <= 1; play_W(8, 169) <= 1; play_W(8, 170) <= 1; play_W(8, 171) <= 0; play_W(8, 172) <= 0; play_W(8, 173) <= 0; play_W(8, 174) <= 0; play_W(8, 175) <= 0; play_W(8, 176) <= 0; play_W(8, 177) <= 1; play_W(8, 178) <= 1; play_W(8, 179) <= 1; play_W(8, 180) <= 1; play_W(8, 181) <= 1; play_W(8, 182) <= 1; play_W(8, 183) <= 0; play_W(8, 184) <= 0; play_W(8, 185) <= 0; play_W(8, 186) <= 0; play_W(8, 187) <= 0; play_W(8, 188) <= 0; play_W(8, 189) <= 1; play_W(8, 190) <= 1; play_W(8, 191) <= 1; play_W(8, 192) <= 0; play_W(8, 193) <= 0; play_W(8, 194) <= 0; play_W(8, 195) <= 0; play_W(8, 196) <= 0; play_W(8, 197) <= 0; play_W(8, 198) <= 1; play_W(8, 199) <= 1; play_W(8, 200) <= 1; play_W(8, 201) <= 1; play_W(8, 202) <= 1; play_W(8, 203) <= 1; play_W(8, 204) <= 0; play_W(8, 205) <= 0; play_W(8, 206) <= 0; play_W(8, 207) <= 0; play_W(8, 208) <= 0; play_W(8, 209) <= 0; play_W(8, 210) <= 1; play_W(8, 211) <= 1; play_W(8, 212) <= 1; play_W(8, 213) <= 0; play_W(8, 214) <= 0; play_W(8, 215) <= 0; play_W(8, 216) <= 1; play_W(8, 217) <= 1; play_W(8, 218) <= 1; play_W(8, 219) <= 1; play_W(8, 220) <= 1; play_W(8, 221) <= 1; play_W(8, 222) <= 1; play_W(8, 223) <= 1; play_W(8, 224) <= 1; play_W(8, 225) <= 1; play_W(8, 226) <= 1; play_W(8, 227) <= 1; play_W(8, 228) <= 0; play_W(8, 229) <= 0; play_W(8, 230) <= 0; play_W(8, 231) <= 1; play_W(8, 232) <= 1; play_W(8, 233) <= 1; play_W(8, 234) <= 1; play_W(8, 235) <= 1; play_W(8, 236) <= 1; play_W(8, 237) <= 0; play_W(8, 238) <= 0; play_W(8, 239) <= 0; play_W(8, 240) <= 0; play_W(8, 241) <= 0; play_W(8, 242) <= 0; play_W(8, 243) <= 0; play_W(8, 244) <= 0; play_W(8, 245) <= 0; play_W(8, 246) <= 1; play_W(8, 247) <= 1; play_W(8, 248) <= 1; play_W(8, 249) <= 1; play_W(8, 250) <= 1; play_W(8, 251) <= 1; play_W(8, 252) <= 0; play_W(8, 253) <= 0; play_W(8, 254) <= 0; play_W(8, 255) <= 0; play_W(8, 256) <= 0; play_W(8, 257) <= 0; play_W(8, 258) <= 1; play_W(8, 259) <= 1; play_W(8, 260) <= 1; play_W(8, 261) <= 1; play_W(8, 262) <= 1; play_W(8, 263) <= 1; play_W(8, 264) <= 0; play_W(8, 265) <= 0; play_W(8, 266) <= 0; play_W(8, 267) <= 0; play_W(8, 268) <= 0; play_W(8, 269) <= 0; 
play_W(9, 0) <= 0; play_W(9, 1) <= 0; play_W(9, 2) <= 0; play_W(9, 3) <= 1; play_W(9, 4) <= 1; play_W(9, 5) <= 1; play_W(9, 6) <= 1; play_W(9, 7) <= 1; play_W(9, 8) <= 1; play_W(9, 9) <= 0; play_W(9, 10) <= 0; play_W(9, 11) <= 0; play_W(9, 12) <= 0; play_W(9, 13) <= 0; play_W(9, 14) <= 0; play_W(9, 15) <= 1; play_W(9, 16) <= 1; play_W(9, 17) <= 1; play_W(9, 18) <= 1; play_W(9, 19) <= 1; play_W(9, 20) <= 1; play_W(9, 21) <= 0; play_W(9, 22) <= 0; play_W(9, 23) <= 0; play_W(9, 24) <= 0; play_W(9, 25) <= 0; play_W(9, 26) <= 0; play_W(9, 27) <= 0; play_W(9, 28) <= 0; play_W(9, 29) <= 0; play_W(9, 30) <= 1; play_W(9, 31) <= 1; play_W(9, 32) <= 1; play_W(9, 33) <= 1; play_W(9, 34) <= 1; play_W(9, 35) <= 1; play_W(9, 36) <= 0; play_W(9, 37) <= 0; play_W(9, 38) <= 0; play_W(9, 39) <= 0; play_W(9, 40) <= 0; play_W(9, 41) <= 0; play_W(9, 42) <= 0; play_W(9, 43) <= 0; play_W(9, 44) <= 0; play_W(9, 45) <= 0; play_W(9, 46) <= 0; play_W(9, 47) <= 0; play_W(9, 48) <= 0; play_W(9, 49) <= 0; play_W(9, 50) <= 0; play_W(9, 51) <= 0; play_W(9, 52) <= 0; play_W(9, 53) <= 0; play_W(9, 54) <= 1; play_W(9, 55) <= 1; play_W(9, 56) <= 1; play_W(9, 57) <= 1; play_W(9, 58) <= 1; play_W(9, 59) <= 1; play_W(9, 60) <= 0; play_W(9, 61) <= 0; play_W(9, 62) <= 0; play_W(9, 63) <= 0; play_W(9, 64) <= 0; play_W(9, 65) <= 0; play_W(9, 66) <= 0; play_W(9, 67) <= 0; play_W(9, 68) <= 0; play_W(9, 69) <= 1; play_W(9, 70) <= 1; play_W(9, 71) <= 1; play_W(9, 72) <= 1; play_W(9, 73) <= 1; play_W(9, 74) <= 1; play_W(9, 75) <= 0; play_W(9, 76) <= 0; play_W(9, 77) <= 0; play_W(9, 78) <= 0; play_W(9, 79) <= 0; play_W(9, 80) <= 0; play_W(9, 81) <= 0; play_W(9, 82) <= 0; play_W(9, 83) <= 0; play_W(9, 84) <= 1; play_W(9, 85) <= 1; play_W(9, 86) <= 1; play_W(9, 87) <= 1; play_W(9, 88) <= 1; play_W(9, 89) <= 1; play_W(9, 90) <= 0; play_W(9, 91) <= 0; play_W(9, 92) <= 0; play_W(9, 93) <= 0; play_W(9, 94) <= 0; play_W(9, 95) <= 0; play_W(9, 96) <= 1; play_W(9, 97) <= 1; play_W(9, 98) <= 1; play_W(9, 99) <= 1; play_W(9, 100) <= 1; play_W(9, 101) <= 1; play_W(9, 102) <= 0; play_W(9, 103) <= 0; play_W(9, 104) <= 0; play_W(9, 105) <= 0; play_W(9, 106) <= 0; play_W(9, 107) <= 0; play_W(9, 108) <= 0; play_W(9, 109) <= 0; play_W(9, 110) <= 0; play_W(9, 111) <= 0; play_W(9, 112) <= 0; play_W(9, 113) <= 0; play_W(9, 114) <= 0; play_W(9, 115) <= 0; play_W(9, 116) <= 0; play_W(9, 117) <= 1; play_W(9, 118) <= 1; play_W(9, 119) <= 1; play_W(9, 120) <= 1; play_W(9, 121) <= 1; play_W(9, 122) <= 1; play_W(9, 123) <= 0; play_W(9, 124) <= 0; play_W(9, 125) <= 0; play_W(9, 126) <= 0; play_W(9, 127) <= 0; play_W(9, 128) <= 0; play_W(9, 129) <= 0; play_W(9, 130) <= 0; play_W(9, 131) <= 0; play_W(9, 132) <= 0; play_W(9, 133) <= 0; play_W(9, 134) <= 0; play_W(9, 135) <= 0; play_W(9, 136) <= 0; play_W(9, 137) <= 0; play_W(9, 138) <= 0; play_W(9, 139) <= 0; play_W(9, 140) <= 0; play_W(9, 141) <= 0; play_W(9, 142) <= 0; play_W(9, 143) <= 0; play_W(9, 144) <= 0; play_W(9, 145) <= 0; play_W(9, 146) <= 0; play_W(9, 147) <= 0; play_W(9, 148) <= 0; play_W(9, 149) <= 0; play_W(9, 150) <= 0; play_W(9, 151) <= 0; play_W(9, 152) <= 0; play_W(9, 153) <= 0; play_W(9, 154) <= 0; play_W(9, 155) <= 0; play_W(9, 156) <= 0; play_W(9, 157) <= 0; play_W(9, 158) <= 0; play_W(9, 159) <= 0; play_W(9, 160) <= 0; play_W(9, 161) <= 0; play_W(9, 162) <= 0; play_W(9, 163) <= 0; play_W(9, 164) <= 0; play_W(9, 165) <= 1; play_W(9, 166) <= 1; play_W(9, 167) <= 1; play_W(9, 168) <= 1; play_W(9, 169) <= 1; play_W(9, 170) <= 1; play_W(9, 171) <= 0; play_W(9, 172) <= 0; play_W(9, 173) <= 0; play_W(9, 174) <= 0; play_W(9, 175) <= 0; play_W(9, 176) <= 0; play_W(9, 177) <= 1; play_W(9, 178) <= 1; play_W(9, 179) <= 1; play_W(9, 180) <= 1; play_W(9, 181) <= 1; play_W(9, 182) <= 1; play_W(9, 183) <= 0; play_W(9, 184) <= 0; play_W(9, 185) <= 0; play_W(9, 186) <= 0; play_W(9, 187) <= 0; play_W(9, 188) <= 0; play_W(9, 189) <= 0; play_W(9, 190) <= 0; play_W(9, 191) <= 0; play_W(9, 192) <= 0; play_W(9, 193) <= 0; play_W(9, 194) <= 0; play_W(9, 195) <= 0; play_W(9, 196) <= 0; play_W(9, 197) <= 0; play_W(9, 198) <= 1; play_W(9, 199) <= 1; play_W(9, 200) <= 1; play_W(9, 201) <= 1; play_W(9, 202) <= 1; play_W(9, 203) <= 1; play_W(9, 204) <= 0; play_W(9, 205) <= 0; play_W(9, 206) <= 0; play_W(9, 207) <= 0; play_W(9, 208) <= 0; play_W(9, 209) <= 0; play_W(9, 210) <= 0; play_W(9, 211) <= 0; play_W(9, 212) <= 0; play_W(9, 213) <= 0; play_W(9, 214) <= 0; play_W(9, 215) <= 0; play_W(9, 216) <= 1; play_W(9, 217) <= 1; play_W(9, 218) <= 1; play_W(9, 219) <= 1; play_W(9, 220) <= 1; play_W(9, 221) <= 1; play_W(9, 222) <= 1; play_W(9, 223) <= 1; play_W(9, 224) <= 1; play_W(9, 225) <= 1; play_W(9, 226) <= 1; play_W(9, 227) <= 1; play_W(9, 228) <= 1; play_W(9, 229) <= 1; play_W(9, 230) <= 1; play_W(9, 231) <= 1; play_W(9, 232) <= 1; play_W(9, 233) <= 1; play_W(9, 234) <= 1; play_W(9, 235) <= 1; play_W(9, 236) <= 1; play_W(9, 237) <= 0; play_W(9, 238) <= 0; play_W(9, 239) <= 0; play_W(9, 240) <= 0; play_W(9, 241) <= 0; play_W(9, 242) <= 0; play_W(9, 243) <= 0; play_W(9, 244) <= 0; play_W(9, 245) <= 0; play_W(9, 246) <= 1; play_W(9, 247) <= 1; play_W(9, 248) <= 1; play_W(9, 249) <= 1; play_W(9, 250) <= 1; play_W(9, 251) <= 1; play_W(9, 252) <= 0; play_W(9, 253) <= 0; play_W(9, 254) <= 0; play_W(9, 255) <= 0; play_W(9, 256) <= 0; play_W(9, 257) <= 0; play_W(9, 258) <= 1; play_W(9, 259) <= 1; play_W(9, 260) <= 1; play_W(9, 261) <= 1; play_W(9, 262) <= 1; play_W(9, 263) <= 1; play_W(9, 264) <= 0; play_W(9, 265) <= 0; play_W(9, 266) <= 0; play_W(9, 267) <= 0; play_W(9, 268) <= 0; play_W(9, 269) <= 0; 
play_W(10, 0) <= 0; play_W(10, 1) <= 0; play_W(10, 2) <= 0; play_W(10, 3) <= 1; play_W(10, 4) <= 1; play_W(10, 5) <= 1; play_W(10, 6) <= 1; play_W(10, 7) <= 1; play_W(10, 8) <= 1; play_W(10, 9) <= 0; play_W(10, 10) <= 0; play_W(10, 11) <= 0; play_W(10, 12) <= 0; play_W(10, 13) <= 0; play_W(10, 14) <= 0; play_W(10, 15) <= 1; play_W(10, 16) <= 1; play_W(10, 17) <= 1; play_W(10, 18) <= 1; play_W(10, 19) <= 1; play_W(10, 20) <= 1; play_W(10, 21) <= 0; play_W(10, 22) <= 0; play_W(10, 23) <= 0; play_W(10, 24) <= 0; play_W(10, 25) <= 0; play_W(10, 26) <= 0; play_W(10, 27) <= 0; play_W(10, 28) <= 0; play_W(10, 29) <= 0; play_W(10, 30) <= 1; play_W(10, 31) <= 1; play_W(10, 32) <= 1; play_W(10, 33) <= 1; play_W(10, 34) <= 1; play_W(10, 35) <= 1; play_W(10, 36) <= 0; play_W(10, 37) <= 0; play_W(10, 38) <= 0; play_W(10, 39) <= 0; play_W(10, 40) <= 0; play_W(10, 41) <= 0; play_W(10, 42) <= 0; play_W(10, 43) <= 0; play_W(10, 44) <= 0; play_W(10, 45) <= 0; play_W(10, 46) <= 0; play_W(10, 47) <= 0; play_W(10, 48) <= 0; play_W(10, 49) <= 0; play_W(10, 50) <= 0; play_W(10, 51) <= 0; play_W(10, 52) <= 0; play_W(10, 53) <= 0; play_W(10, 54) <= 1; play_W(10, 55) <= 1; play_W(10, 56) <= 1; play_W(10, 57) <= 1; play_W(10, 58) <= 1; play_W(10, 59) <= 1; play_W(10, 60) <= 0; play_W(10, 61) <= 0; play_W(10, 62) <= 0; play_W(10, 63) <= 0; play_W(10, 64) <= 0; play_W(10, 65) <= 0; play_W(10, 66) <= 0; play_W(10, 67) <= 0; play_W(10, 68) <= 0; play_W(10, 69) <= 1; play_W(10, 70) <= 1; play_W(10, 71) <= 1; play_W(10, 72) <= 1; play_W(10, 73) <= 1; play_W(10, 74) <= 1; play_W(10, 75) <= 0; play_W(10, 76) <= 0; play_W(10, 77) <= 0; play_W(10, 78) <= 0; play_W(10, 79) <= 0; play_W(10, 80) <= 0; play_W(10, 81) <= 0; play_W(10, 82) <= 0; play_W(10, 83) <= 0; play_W(10, 84) <= 1; play_W(10, 85) <= 1; play_W(10, 86) <= 1; play_W(10, 87) <= 1; play_W(10, 88) <= 1; play_W(10, 89) <= 1; play_W(10, 90) <= 0; play_W(10, 91) <= 0; play_W(10, 92) <= 0; play_W(10, 93) <= 0; play_W(10, 94) <= 0; play_W(10, 95) <= 0; play_W(10, 96) <= 1; play_W(10, 97) <= 1; play_W(10, 98) <= 1; play_W(10, 99) <= 1; play_W(10, 100) <= 1; play_W(10, 101) <= 1; play_W(10, 102) <= 0; play_W(10, 103) <= 0; play_W(10, 104) <= 0; play_W(10, 105) <= 0; play_W(10, 106) <= 0; play_W(10, 107) <= 0; play_W(10, 108) <= 0; play_W(10, 109) <= 0; play_W(10, 110) <= 0; play_W(10, 111) <= 0; play_W(10, 112) <= 0; play_W(10, 113) <= 0; play_W(10, 114) <= 0; play_W(10, 115) <= 0; play_W(10, 116) <= 0; play_W(10, 117) <= 1; play_W(10, 118) <= 1; play_W(10, 119) <= 1; play_W(10, 120) <= 1; play_W(10, 121) <= 1; play_W(10, 122) <= 1; play_W(10, 123) <= 0; play_W(10, 124) <= 0; play_W(10, 125) <= 0; play_W(10, 126) <= 0; play_W(10, 127) <= 0; play_W(10, 128) <= 0; play_W(10, 129) <= 0; play_W(10, 130) <= 0; play_W(10, 131) <= 0; play_W(10, 132) <= 0; play_W(10, 133) <= 0; play_W(10, 134) <= 0; play_W(10, 135) <= 0; play_W(10, 136) <= 0; play_W(10, 137) <= 0; play_W(10, 138) <= 0; play_W(10, 139) <= 0; play_W(10, 140) <= 0; play_W(10, 141) <= 0; play_W(10, 142) <= 0; play_W(10, 143) <= 0; play_W(10, 144) <= 0; play_W(10, 145) <= 0; play_W(10, 146) <= 0; play_W(10, 147) <= 0; play_W(10, 148) <= 0; play_W(10, 149) <= 0; play_W(10, 150) <= 0; play_W(10, 151) <= 0; play_W(10, 152) <= 0; play_W(10, 153) <= 0; play_W(10, 154) <= 0; play_W(10, 155) <= 0; play_W(10, 156) <= 0; play_W(10, 157) <= 0; play_W(10, 158) <= 0; play_W(10, 159) <= 0; play_W(10, 160) <= 0; play_W(10, 161) <= 0; play_W(10, 162) <= 0; play_W(10, 163) <= 0; play_W(10, 164) <= 0; play_W(10, 165) <= 1; play_W(10, 166) <= 1; play_W(10, 167) <= 1; play_W(10, 168) <= 1; play_W(10, 169) <= 1; play_W(10, 170) <= 1; play_W(10, 171) <= 0; play_W(10, 172) <= 0; play_W(10, 173) <= 0; play_W(10, 174) <= 0; play_W(10, 175) <= 0; play_W(10, 176) <= 0; play_W(10, 177) <= 1; play_W(10, 178) <= 1; play_W(10, 179) <= 1; play_W(10, 180) <= 1; play_W(10, 181) <= 1; play_W(10, 182) <= 1; play_W(10, 183) <= 0; play_W(10, 184) <= 0; play_W(10, 185) <= 0; play_W(10, 186) <= 0; play_W(10, 187) <= 0; play_W(10, 188) <= 0; play_W(10, 189) <= 0; play_W(10, 190) <= 0; play_W(10, 191) <= 0; play_W(10, 192) <= 0; play_W(10, 193) <= 0; play_W(10, 194) <= 0; play_W(10, 195) <= 0; play_W(10, 196) <= 0; play_W(10, 197) <= 0; play_W(10, 198) <= 1; play_W(10, 199) <= 1; play_W(10, 200) <= 1; play_W(10, 201) <= 1; play_W(10, 202) <= 1; play_W(10, 203) <= 1; play_W(10, 204) <= 0; play_W(10, 205) <= 0; play_W(10, 206) <= 0; play_W(10, 207) <= 0; play_W(10, 208) <= 0; play_W(10, 209) <= 0; play_W(10, 210) <= 0; play_W(10, 211) <= 0; play_W(10, 212) <= 0; play_W(10, 213) <= 0; play_W(10, 214) <= 0; play_W(10, 215) <= 0; play_W(10, 216) <= 1; play_W(10, 217) <= 1; play_W(10, 218) <= 1; play_W(10, 219) <= 1; play_W(10, 220) <= 1; play_W(10, 221) <= 1; play_W(10, 222) <= 1; play_W(10, 223) <= 1; play_W(10, 224) <= 1; play_W(10, 225) <= 1; play_W(10, 226) <= 1; play_W(10, 227) <= 1; play_W(10, 228) <= 1; play_W(10, 229) <= 1; play_W(10, 230) <= 1; play_W(10, 231) <= 1; play_W(10, 232) <= 1; play_W(10, 233) <= 1; play_W(10, 234) <= 1; play_W(10, 235) <= 1; play_W(10, 236) <= 1; play_W(10, 237) <= 0; play_W(10, 238) <= 0; play_W(10, 239) <= 0; play_W(10, 240) <= 0; play_W(10, 241) <= 0; play_W(10, 242) <= 0; play_W(10, 243) <= 0; play_W(10, 244) <= 0; play_W(10, 245) <= 0; play_W(10, 246) <= 1; play_W(10, 247) <= 1; play_W(10, 248) <= 1; play_W(10, 249) <= 1; play_W(10, 250) <= 1; play_W(10, 251) <= 1; play_W(10, 252) <= 0; play_W(10, 253) <= 0; play_W(10, 254) <= 0; play_W(10, 255) <= 0; play_W(10, 256) <= 0; play_W(10, 257) <= 0; play_W(10, 258) <= 1; play_W(10, 259) <= 1; play_W(10, 260) <= 1; play_W(10, 261) <= 1; play_W(10, 262) <= 1; play_W(10, 263) <= 1; play_W(10, 264) <= 0; play_W(10, 265) <= 0; play_W(10, 266) <= 0; play_W(10, 267) <= 0; play_W(10, 268) <= 0; play_W(10, 269) <= 0; 
play_W(11, 0) <= 0; play_W(11, 1) <= 0; play_W(11, 2) <= 0; play_W(11, 3) <= 1; play_W(11, 4) <= 1; play_W(11, 5) <= 1; play_W(11, 6) <= 1; play_W(11, 7) <= 1; play_W(11, 8) <= 1; play_W(11, 9) <= 0; play_W(11, 10) <= 0; play_W(11, 11) <= 0; play_W(11, 12) <= 0; play_W(11, 13) <= 0; play_W(11, 14) <= 0; play_W(11, 15) <= 1; play_W(11, 16) <= 1; play_W(11, 17) <= 1; play_W(11, 18) <= 1; play_W(11, 19) <= 1; play_W(11, 20) <= 1; play_W(11, 21) <= 0; play_W(11, 22) <= 0; play_W(11, 23) <= 0; play_W(11, 24) <= 0; play_W(11, 25) <= 0; play_W(11, 26) <= 0; play_W(11, 27) <= 0; play_W(11, 28) <= 0; play_W(11, 29) <= 0; play_W(11, 30) <= 1; play_W(11, 31) <= 1; play_W(11, 32) <= 1; play_W(11, 33) <= 1; play_W(11, 34) <= 1; play_W(11, 35) <= 1; play_W(11, 36) <= 0; play_W(11, 37) <= 0; play_W(11, 38) <= 0; play_W(11, 39) <= 0; play_W(11, 40) <= 0; play_W(11, 41) <= 0; play_W(11, 42) <= 0; play_W(11, 43) <= 0; play_W(11, 44) <= 0; play_W(11, 45) <= 0; play_W(11, 46) <= 0; play_W(11, 47) <= 0; play_W(11, 48) <= 0; play_W(11, 49) <= 0; play_W(11, 50) <= 0; play_W(11, 51) <= 0; play_W(11, 52) <= 0; play_W(11, 53) <= 0; play_W(11, 54) <= 1; play_W(11, 55) <= 1; play_W(11, 56) <= 1; play_W(11, 57) <= 1; play_W(11, 58) <= 1; play_W(11, 59) <= 1; play_W(11, 60) <= 0; play_W(11, 61) <= 0; play_W(11, 62) <= 0; play_W(11, 63) <= 0; play_W(11, 64) <= 0; play_W(11, 65) <= 0; play_W(11, 66) <= 0; play_W(11, 67) <= 0; play_W(11, 68) <= 0; play_W(11, 69) <= 1; play_W(11, 70) <= 1; play_W(11, 71) <= 1; play_W(11, 72) <= 1; play_W(11, 73) <= 1; play_W(11, 74) <= 1; play_W(11, 75) <= 0; play_W(11, 76) <= 0; play_W(11, 77) <= 0; play_W(11, 78) <= 0; play_W(11, 79) <= 0; play_W(11, 80) <= 0; play_W(11, 81) <= 0; play_W(11, 82) <= 0; play_W(11, 83) <= 0; play_W(11, 84) <= 1; play_W(11, 85) <= 1; play_W(11, 86) <= 1; play_W(11, 87) <= 1; play_W(11, 88) <= 1; play_W(11, 89) <= 1; play_W(11, 90) <= 0; play_W(11, 91) <= 0; play_W(11, 92) <= 0; play_W(11, 93) <= 0; play_W(11, 94) <= 0; play_W(11, 95) <= 0; play_W(11, 96) <= 1; play_W(11, 97) <= 1; play_W(11, 98) <= 1; play_W(11, 99) <= 1; play_W(11, 100) <= 1; play_W(11, 101) <= 1; play_W(11, 102) <= 0; play_W(11, 103) <= 0; play_W(11, 104) <= 0; play_W(11, 105) <= 0; play_W(11, 106) <= 0; play_W(11, 107) <= 0; play_W(11, 108) <= 0; play_W(11, 109) <= 0; play_W(11, 110) <= 0; play_W(11, 111) <= 0; play_W(11, 112) <= 0; play_W(11, 113) <= 0; play_W(11, 114) <= 0; play_W(11, 115) <= 0; play_W(11, 116) <= 0; play_W(11, 117) <= 1; play_W(11, 118) <= 1; play_W(11, 119) <= 1; play_W(11, 120) <= 1; play_W(11, 121) <= 1; play_W(11, 122) <= 1; play_W(11, 123) <= 0; play_W(11, 124) <= 0; play_W(11, 125) <= 0; play_W(11, 126) <= 0; play_W(11, 127) <= 0; play_W(11, 128) <= 0; play_W(11, 129) <= 0; play_W(11, 130) <= 0; play_W(11, 131) <= 0; play_W(11, 132) <= 0; play_W(11, 133) <= 0; play_W(11, 134) <= 0; play_W(11, 135) <= 0; play_W(11, 136) <= 0; play_W(11, 137) <= 0; play_W(11, 138) <= 0; play_W(11, 139) <= 0; play_W(11, 140) <= 0; play_W(11, 141) <= 0; play_W(11, 142) <= 0; play_W(11, 143) <= 0; play_W(11, 144) <= 0; play_W(11, 145) <= 0; play_W(11, 146) <= 0; play_W(11, 147) <= 0; play_W(11, 148) <= 0; play_W(11, 149) <= 0; play_W(11, 150) <= 0; play_W(11, 151) <= 0; play_W(11, 152) <= 0; play_W(11, 153) <= 0; play_W(11, 154) <= 0; play_W(11, 155) <= 0; play_W(11, 156) <= 0; play_W(11, 157) <= 0; play_W(11, 158) <= 0; play_W(11, 159) <= 0; play_W(11, 160) <= 0; play_W(11, 161) <= 0; play_W(11, 162) <= 0; play_W(11, 163) <= 0; play_W(11, 164) <= 0; play_W(11, 165) <= 1; play_W(11, 166) <= 1; play_W(11, 167) <= 1; play_W(11, 168) <= 1; play_W(11, 169) <= 1; play_W(11, 170) <= 1; play_W(11, 171) <= 0; play_W(11, 172) <= 0; play_W(11, 173) <= 0; play_W(11, 174) <= 0; play_W(11, 175) <= 0; play_W(11, 176) <= 0; play_W(11, 177) <= 1; play_W(11, 178) <= 1; play_W(11, 179) <= 1; play_W(11, 180) <= 1; play_W(11, 181) <= 1; play_W(11, 182) <= 1; play_W(11, 183) <= 0; play_W(11, 184) <= 0; play_W(11, 185) <= 0; play_W(11, 186) <= 0; play_W(11, 187) <= 0; play_W(11, 188) <= 0; play_W(11, 189) <= 0; play_W(11, 190) <= 0; play_W(11, 191) <= 0; play_W(11, 192) <= 0; play_W(11, 193) <= 0; play_W(11, 194) <= 0; play_W(11, 195) <= 0; play_W(11, 196) <= 0; play_W(11, 197) <= 0; play_W(11, 198) <= 1; play_W(11, 199) <= 1; play_W(11, 200) <= 1; play_W(11, 201) <= 1; play_W(11, 202) <= 1; play_W(11, 203) <= 1; play_W(11, 204) <= 0; play_W(11, 205) <= 0; play_W(11, 206) <= 0; play_W(11, 207) <= 0; play_W(11, 208) <= 0; play_W(11, 209) <= 0; play_W(11, 210) <= 0; play_W(11, 211) <= 0; play_W(11, 212) <= 0; play_W(11, 213) <= 0; play_W(11, 214) <= 0; play_W(11, 215) <= 0; play_W(11, 216) <= 1; play_W(11, 217) <= 1; play_W(11, 218) <= 1; play_W(11, 219) <= 1; play_W(11, 220) <= 1; play_W(11, 221) <= 1; play_W(11, 222) <= 1; play_W(11, 223) <= 1; play_W(11, 224) <= 1; play_W(11, 225) <= 1; play_W(11, 226) <= 1; play_W(11, 227) <= 1; play_W(11, 228) <= 1; play_W(11, 229) <= 1; play_W(11, 230) <= 1; play_W(11, 231) <= 1; play_W(11, 232) <= 1; play_W(11, 233) <= 1; play_W(11, 234) <= 1; play_W(11, 235) <= 1; play_W(11, 236) <= 1; play_W(11, 237) <= 0; play_W(11, 238) <= 0; play_W(11, 239) <= 0; play_W(11, 240) <= 0; play_W(11, 241) <= 0; play_W(11, 242) <= 0; play_W(11, 243) <= 0; play_W(11, 244) <= 0; play_W(11, 245) <= 0; play_W(11, 246) <= 1; play_W(11, 247) <= 1; play_W(11, 248) <= 1; play_W(11, 249) <= 1; play_W(11, 250) <= 1; play_W(11, 251) <= 1; play_W(11, 252) <= 0; play_W(11, 253) <= 0; play_W(11, 254) <= 0; play_W(11, 255) <= 0; play_W(11, 256) <= 0; play_W(11, 257) <= 0; play_W(11, 258) <= 1; play_W(11, 259) <= 1; play_W(11, 260) <= 1; play_W(11, 261) <= 1; play_W(11, 262) <= 1; play_W(11, 263) <= 1; play_W(11, 264) <= 0; play_W(11, 265) <= 0; play_W(11, 266) <= 0; play_W(11, 267) <= 0; play_W(11, 268) <= 0; play_W(11, 269) <= 0; 
play_W(12, 0) <= 0; play_W(12, 1) <= 0; play_W(12, 2) <= 0; play_W(12, 3) <= 1; play_W(12, 4) <= 1; play_W(12, 5) <= 1; play_W(12, 6) <= 1; play_W(12, 7) <= 1; play_W(12, 8) <= 1; play_W(12, 9) <= 1; play_W(12, 10) <= 1; play_W(12, 11) <= 1; play_W(12, 12) <= 1; play_W(12, 13) <= 1; play_W(12, 14) <= 1; play_W(12, 15) <= 1; play_W(12, 16) <= 1; play_W(12, 17) <= 1; play_W(12, 18) <= 0; play_W(12, 19) <= 0; play_W(12, 20) <= 0; play_W(12, 21) <= 0; play_W(12, 22) <= 0; play_W(12, 23) <= 0; play_W(12, 24) <= 0; play_W(12, 25) <= 0; play_W(12, 26) <= 0; play_W(12, 27) <= 0; play_W(12, 28) <= 0; play_W(12, 29) <= 0; play_W(12, 30) <= 1; play_W(12, 31) <= 1; play_W(12, 32) <= 1; play_W(12, 33) <= 1; play_W(12, 34) <= 1; play_W(12, 35) <= 1; play_W(12, 36) <= 0; play_W(12, 37) <= 0; play_W(12, 38) <= 0; play_W(12, 39) <= 0; play_W(12, 40) <= 0; play_W(12, 41) <= 0; play_W(12, 42) <= 0; play_W(12, 43) <= 0; play_W(12, 44) <= 0; play_W(12, 45) <= 0; play_W(12, 46) <= 0; play_W(12, 47) <= 0; play_W(12, 48) <= 0; play_W(12, 49) <= 0; play_W(12, 50) <= 0; play_W(12, 51) <= 0; play_W(12, 52) <= 0; play_W(12, 53) <= 0; play_W(12, 54) <= 1; play_W(12, 55) <= 1; play_W(12, 56) <= 1; play_W(12, 57) <= 1; play_W(12, 58) <= 1; play_W(12, 59) <= 1; play_W(12, 60) <= 0; play_W(12, 61) <= 0; play_W(12, 62) <= 0; play_W(12, 63) <= 0; play_W(12, 64) <= 0; play_W(12, 65) <= 0; play_W(12, 66) <= 0; play_W(12, 67) <= 0; play_W(12, 68) <= 0; play_W(12, 69) <= 1; play_W(12, 70) <= 1; play_W(12, 71) <= 1; play_W(12, 72) <= 1; play_W(12, 73) <= 1; play_W(12, 74) <= 1; play_W(12, 75) <= 0; play_W(12, 76) <= 0; play_W(12, 77) <= 0; play_W(12, 78) <= 0; play_W(12, 79) <= 0; play_W(12, 80) <= 0; play_W(12, 81) <= 0; play_W(12, 82) <= 0; play_W(12, 83) <= 0; play_W(12, 84) <= 0; play_W(12, 85) <= 0; play_W(12, 86) <= 0; play_W(12, 87) <= 1; play_W(12, 88) <= 1; play_W(12, 89) <= 1; play_W(12, 90) <= 1; play_W(12, 91) <= 1; play_W(12, 92) <= 1; play_W(12, 93) <= 1; play_W(12, 94) <= 1; play_W(12, 95) <= 1; play_W(12, 96) <= 1; play_W(12, 97) <= 1; play_W(12, 98) <= 1; play_W(12, 99) <= 0; play_W(12, 100) <= 0; play_W(12, 101) <= 0; play_W(12, 102) <= 0; play_W(12, 103) <= 0; play_W(12, 104) <= 0; play_W(12, 105) <= 0; play_W(12, 106) <= 0; play_W(12, 107) <= 0; play_W(12, 108) <= 0; play_W(12, 109) <= 0; play_W(12, 110) <= 0; play_W(12, 111) <= 0; play_W(12, 112) <= 0; play_W(12, 113) <= 0; play_W(12, 114) <= 0; play_W(12, 115) <= 0; play_W(12, 116) <= 0; play_W(12, 117) <= 0; play_W(12, 118) <= 0; play_W(12, 119) <= 0; play_W(12, 120) <= 0; play_W(12, 121) <= 0; play_W(12, 122) <= 0; play_W(12, 123) <= 0; play_W(12, 124) <= 0; play_W(12, 125) <= 0; play_W(12, 126) <= 0; play_W(12, 127) <= 0; play_W(12, 128) <= 0; play_W(12, 129) <= 0; play_W(12, 130) <= 0; play_W(12, 131) <= 0; play_W(12, 132) <= 0; play_W(12, 133) <= 0; play_W(12, 134) <= 0; play_W(12, 135) <= 0; play_W(12, 136) <= 0; play_W(12, 137) <= 0; play_W(12, 138) <= 0; play_W(12, 139) <= 0; play_W(12, 140) <= 0; play_W(12, 141) <= 0; play_W(12, 142) <= 0; play_W(12, 143) <= 0; play_W(12, 144) <= 0; play_W(12, 145) <= 0; play_W(12, 146) <= 0; play_W(12, 147) <= 0; play_W(12, 148) <= 0; play_W(12, 149) <= 0; play_W(12, 150) <= 0; play_W(12, 151) <= 0; play_W(12, 152) <= 0; play_W(12, 153) <= 0; play_W(12, 154) <= 0; play_W(12, 155) <= 0; play_W(12, 156) <= 0; play_W(12, 157) <= 0; play_W(12, 158) <= 0; play_W(12, 159) <= 0; play_W(12, 160) <= 0; play_W(12, 161) <= 0; play_W(12, 162) <= 0; play_W(12, 163) <= 0; play_W(12, 164) <= 0; play_W(12, 165) <= 1; play_W(12, 166) <= 1; play_W(12, 167) <= 1; play_W(12, 168) <= 1; play_W(12, 169) <= 1; play_W(12, 170) <= 1; play_W(12, 171) <= 1; play_W(12, 172) <= 1; play_W(12, 173) <= 1; play_W(12, 174) <= 1; play_W(12, 175) <= 1; play_W(12, 176) <= 1; play_W(12, 177) <= 1; play_W(12, 178) <= 1; play_W(12, 179) <= 1; play_W(12, 180) <= 0; play_W(12, 181) <= 0; play_W(12, 182) <= 0; play_W(12, 183) <= 0; play_W(12, 184) <= 0; play_W(12, 185) <= 0; play_W(12, 186) <= 0; play_W(12, 187) <= 0; play_W(12, 188) <= 0; play_W(12, 189) <= 0; play_W(12, 190) <= 0; play_W(12, 191) <= 0; play_W(12, 192) <= 0; play_W(12, 193) <= 0; play_W(12, 194) <= 0; play_W(12, 195) <= 0; play_W(12, 196) <= 0; play_W(12, 197) <= 0; play_W(12, 198) <= 1; play_W(12, 199) <= 1; play_W(12, 200) <= 1; play_W(12, 201) <= 1; play_W(12, 202) <= 1; play_W(12, 203) <= 1; play_W(12, 204) <= 0; play_W(12, 205) <= 0; play_W(12, 206) <= 0; play_W(12, 207) <= 0; play_W(12, 208) <= 0; play_W(12, 209) <= 0; play_W(12, 210) <= 0; play_W(12, 211) <= 0; play_W(12, 212) <= 0; play_W(12, 213) <= 0; play_W(12, 214) <= 0; play_W(12, 215) <= 0; play_W(12, 216) <= 1; play_W(12, 217) <= 1; play_W(12, 218) <= 1; play_W(12, 219) <= 1; play_W(12, 220) <= 1; play_W(12, 221) <= 1; play_W(12, 222) <= 0; play_W(12, 223) <= 0; play_W(12, 224) <= 0; play_W(12, 225) <= 1; play_W(12, 226) <= 1; play_W(12, 227) <= 1; play_W(12, 228) <= 1; play_W(12, 229) <= 1; play_W(12, 230) <= 1; play_W(12, 231) <= 1; play_W(12, 232) <= 1; play_W(12, 233) <= 1; play_W(12, 234) <= 1; play_W(12, 235) <= 1; play_W(12, 236) <= 1; play_W(12, 237) <= 0; play_W(12, 238) <= 0; play_W(12, 239) <= 0; play_W(12, 240) <= 0; play_W(12, 241) <= 0; play_W(12, 242) <= 0; play_W(12, 243) <= 0; play_W(12, 244) <= 0; play_W(12, 245) <= 0; play_W(12, 246) <= 1; play_W(12, 247) <= 1; play_W(12, 248) <= 1; play_W(12, 249) <= 1; play_W(12, 250) <= 1; play_W(12, 251) <= 1; play_W(12, 252) <= 1; play_W(12, 253) <= 1; play_W(12, 254) <= 1; play_W(12, 255) <= 1; play_W(12, 256) <= 1; play_W(12, 257) <= 1; play_W(12, 258) <= 1; play_W(12, 259) <= 1; play_W(12, 260) <= 1; play_W(12, 261) <= 0; play_W(12, 262) <= 0; play_W(12, 263) <= 0; play_W(12, 264) <= 0; play_W(12, 265) <= 0; play_W(12, 266) <= 0; play_W(12, 267) <= 0; play_W(12, 268) <= 0; play_W(12, 269) <= 0; 
play_W(13, 0) <= 0; play_W(13, 1) <= 0; play_W(13, 2) <= 0; play_W(13, 3) <= 1; play_W(13, 4) <= 1; play_W(13, 5) <= 1; play_W(13, 6) <= 1; play_W(13, 7) <= 1; play_W(13, 8) <= 1; play_W(13, 9) <= 1; play_W(13, 10) <= 1; play_W(13, 11) <= 1; play_W(13, 12) <= 1; play_W(13, 13) <= 1; play_W(13, 14) <= 1; play_W(13, 15) <= 1; play_W(13, 16) <= 1; play_W(13, 17) <= 1; play_W(13, 18) <= 0; play_W(13, 19) <= 0; play_W(13, 20) <= 0; play_W(13, 21) <= 0; play_W(13, 22) <= 0; play_W(13, 23) <= 0; play_W(13, 24) <= 0; play_W(13, 25) <= 0; play_W(13, 26) <= 0; play_W(13, 27) <= 0; play_W(13, 28) <= 0; play_W(13, 29) <= 0; play_W(13, 30) <= 1; play_W(13, 31) <= 1; play_W(13, 32) <= 1; play_W(13, 33) <= 1; play_W(13, 34) <= 1; play_W(13, 35) <= 1; play_W(13, 36) <= 0; play_W(13, 37) <= 0; play_W(13, 38) <= 0; play_W(13, 39) <= 0; play_W(13, 40) <= 0; play_W(13, 41) <= 0; play_W(13, 42) <= 0; play_W(13, 43) <= 0; play_W(13, 44) <= 0; play_W(13, 45) <= 0; play_W(13, 46) <= 0; play_W(13, 47) <= 0; play_W(13, 48) <= 0; play_W(13, 49) <= 0; play_W(13, 50) <= 0; play_W(13, 51) <= 0; play_W(13, 52) <= 0; play_W(13, 53) <= 0; play_W(13, 54) <= 1; play_W(13, 55) <= 1; play_W(13, 56) <= 1; play_W(13, 57) <= 1; play_W(13, 58) <= 1; play_W(13, 59) <= 1; play_W(13, 60) <= 0; play_W(13, 61) <= 0; play_W(13, 62) <= 0; play_W(13, 63) <= 0; play_W(13, 64) <= 0; play_W(13, 65) <= 0; play_W(13, 66) <= 0; play_W(13, 67) <= 0; play_W(13, 68) <= 0; play_W(13, 69) <= 1; play_W(13, 70) <= 1; play_W(13, 71) <= 1; play_W(13, 72) <= 1; play_W(13, 73) <= 1; play_W(13, 74) <= 1; play_W(13, 75) <= 0; play_W(13, 76) <= 0; play_W(13, 77) <= 0; play_W(13, 78) <= 0; play_W(13, 79) <= 0; play_W(13, 80) <= 0; play_W(13, 81) <= 0; play_W(13, 82) <= 0; play_W(13, 83) <= 0; play_W(13, 84) <= 0; play_W(13, 85) <= 0; play_W(13, 86) <= 0; play_W(13, 87) <= 1; play_W(13, 88) <= 1; play_W(13, 89) <= 1; play_W(13, 90) <= 1; play_W(13, 91) <= 1; play_W(13, 92) <= 1; play_W(13, 93) <= 1; play_W(13, 94) <= 1; play_W(13, 95) <= 1; play_W(13, 96) <= 1; play_W(13, 97) <= 1; play_W(13, 98) <= 1; play_W(13, 99) <= 0; play_W(13, 100) <= 0; play_W(13, 101) <= 0; play_W(13, 102) <= 0; play_W(13, 103) <= 0; play_W(13, 104) <= 0; play_W(13, 105) <= 0; play_W(13, 106) <= 0; play_W(13, 107) <= 0; play_W(13, 108) <= 0; play_W(13, 109) <= 0; play_W(13, 110) <= 0; play_W(13, 111) <= 0; play_W(13, 112) <= 0; play_W(13, 113) <= 0; play_W(13, 114) <= 0; play_W(13, 115) <= 0; play_W(13, 116) <= 0; play_W(13, 117) <= 0; play_W(13, 118) <= 0; play_W(13, 119) <= 0; play_W(13, 120) <= 0; play_W(13, 121) <= 0; play_W(13, 122) <= 0; play_W(13, 123) <= 0; play_W(13, 124) <= 0; play_W(13, 125) <= 0; play_W(13, 126) <= 0; play_W(13, 127) <= 0; play_W(13, 128) <= 0; play_W(13, 129) <= 0; play_W(13, 130) <= 0; play_W(13, 131) <= 0; play_W(13, 132) <= 0; play_W(13, 133) <= 0; play_W(13, 134) <= 0; play_W(13, 135) <= 0; play_W(13, 136) <= 0; play_W(13, 137) <= 0; play_W(13, 138) <= 0; play_W(13, 139) <= 0; play_W(13, 140) <= 0; play_W(13, 141) <= 0; play_W(13, 142) <= 0; play_W(13, 143) <= 0; play_W(13, 144) <= 0; play_W(13, 145) <= 0; play_W(13, 146) <= 0; play_W(13, 147) <= 0; play_W(13, 148) <= 0; play_W(13, 149) <= 0; play_W(13, 150) <= 0; play_W(13, 151) <= 0; play_W(13, 152) <= 0; play_W(13, 153) <= 0; play_W(13, 154) <= 0; play_W(13, 155) <= 0; play_W(13, 156) <= 0; play_W(13, 157) <= 0; play_W(13, 158) <= 0; play_W(13, 159) <= 0; play_W(13, 160) <= 0; play_W(13, 161) <= 0; play_W(13, 162) <= 0; play_W(13, 163) <= 0; play_W(13, 164) <= 0; play_W(13, 165) <= 1; play_W(13, 166) <= 1; play_W(13, 167) <= 1; play_W(13, 168) <= 1; play_W(13, 169) <= 1; play_W(13, 170) <= 1; play_W(13, 171) <= 1; play_W(13, 172) <= 1; play_W(13, 173) <= 1; play_W(13, 174) <= 1; play_W(13, 175) <= 1; play_W(13, 176) <= 1; play_W(13, 177) <= 1; play_W(13, 178) <= 1; play_W(13, 179) <= 1; play_W(13, 180) <= 0; play_W(13, 181) <= 0; play_W(13, 182) <= 0; play_W(13, 183) <= 0; play_W(13, 184) <= 0; play_W(13, 185) <= 0; play_W(13, 186) <= 0; play_W(13, 187) <= 0; play_W(13, 188) <= 0; play_W(13, 189) <= 0; play_W(13, 190) <= 0; play_W(13, 191) <= 0; play_W(13, 192) <= 0; play_W(13, 193) <= 0; play_W(13, 194) <= 0; play_W(13, 195) <= 0; play_W(13, 196) <= 0; play_W(13, 197) <= 0; play_W(13, 198) <= 1; play_W(13, 199) <= 1; play_W(13, 200) <= 1; play_W(13, 201) <= 1; play_W(13, 202) <= 1; play_W(13, 203) <= 1; play_W(13, 204) <= 0; play_W(13, 205) <= 0; play_W(13, 206) <= 0; play_W(13, 207) <= 0; play_W(13, 208) <= 0; play_W(13, 209) <= 0; play_W(13, 210) <= 0; play_W(13, 211) <= 0; play_W(13, 212) <= 0; play_W(13, 213) <= 0; play_W(13, 214) <= 0; play_W(13, 215) <= 0; play_W(13, 216) <= 1; play_W(13, 217) <= 1; play_W(13, 218) <= 1; play_W(13, 219) <= 1; play_W(13, 220) <= 1; play_W(13, 221) <= 1; play_W(13, 222) <= 0; play_W(13, 223) <= 0; play_W(13, 224) <= 0; play_W(13, 225) <= 1; play_W(13, 226) <= 1; play_W(13, 227) <= 1; play_W(13, 228) <= 1; play_W(13, 229) <= 1; play_W(13, 230) <= 1; play_W(13, 231) <= 1; play_W(13, 232) <= 1; play_W(13, 233) <= 1; play_W(13, 234) <= 1; play_W(13, 235) <= 1; play_W(13, 236) <= 1; play_W(13, 237) <= 0; play_W(13, 238) <= 0; play_W(13, 239) <= 0; play_W(13, 240) <= 0; play_W(13, 241) <= 0; play_W(13, 242) <= 0; play_W(13, 243) <= 0; play_W(13, 244) <= 0; play_W(13, 245) <= 0; play_W(13, 246) <= 1; play_W(13, 247) <= 1; play_W(13, 248) <= 1; play_W(13, 249) <= 1; play_W(13, 250) <= 1; play_W(13, 251) <= 1; play_W(13, 252) <= 1; play_W(13, 253) <= 1; play_W(13, 254) <= 1; play_W(13, 255) <= 1; play_W(13, 256) <= 1; play_W(13, 257) <= 1; play_W(13, 258) <= 1; play_W(13, 259) <= 1; play_W(13, 260) <= 1; play_W(13, 261) <= 0; play_W(13, 262) <= 0; play_W(13, 263) <= 0; play_W(13, 264) <= 0; play_W(13, 265) <= 0; play_W(13, 266) <= 0; play_W(13, 267) <= 0; play_W(13, 268) <= 0; play_W(13, 269) <= 0; 
play_W(14, 0) <= 0; play_W(14, 1) <= 0; play_W(14, 2) <= 0; play_W(14, 3) <= 1; play_W(14, 4) <= 1; play_W(14, 5) <= 1; play_W(14, 6) <= 1; play_W(14, 7) <= 1; play_W(14, 8) <= 1; play_W(14, 9) <= 1; play_W(14, 10) <= 1; play_W(14, 11) <= 1; play_W(14, 12) <= 1; play_W(14, 13) <= 1; play_W(14, 14) <= 1; play_W(14, 15) <= 1; play_W(14, 16) <= 1; play_W(14, 17) <= 1; play_W(14, 18) <= 0; play_W(14, 19) <= 0; play_W(14, 20) <= 0; play_W(14, 21) <= 0; play_W(14, 22) <= 0; play_W(14, 23) <= 0; play_W(14, 24) <= 0; play_W(14, 25) <= 0; play_W(14, 26) <= 0; play_W(14, 27) <= 0; play_W(14, 28) <= 0; play_W(14, 29) <= 0; play_W(14, 30) <= 1; play_W(14, 31) <= 1; play_W(14, 32) <= 1; play_W(14, 33) <= 1; play_W(14, 34) <= 1; play_W(14, 35) <= 1; play_W(14, 36) <= 0; play_W(14, 37) <= 0; play_W(14, 38) <= 0; play_W(14, 39) <= 0; play_W(14, 40) <= 0; play_W(14, 41) <= 0; play_W(14, 42) <= 0; play_W(14, 43) <= 0; play_W(14, 44) <= 0; play_W(14, 45) <= 0; play_W(14, 46) <= 0; play_W(14, 47) <= 0; play_W(14, 48) <= 0; play_W(14, 49) <= 0; play_W(14, 50) <= 0; play_W(14, 51) <= 0; play_W(14, 52) <= 0; play_W(14, 53) <= 0; play_W(14, 54) <= 1; play_W(14, 55) <= 1; play_W(14, 56) <= 1; play_W(14, 57) <= 1; play_W(14, 58) <= 1; play_W(14, 59) <= 1; play_W(14, 60) <= 0; play_W(14, 61) <= 0; play_W(14, 62) <= 0; play_W(14, 63) <= 0; play_W(14, 64) <= 0; play_W(14, 65) <= 0; play_W(14, 66) <= 0; play_W(14, 67) <= 0; play_W(14, 68) <= 0; play_W(14, 69) <= 1; play_W(14, 70) <= 1; play_W(14, 71) <= 1; play_W(14, 72) <= 1; play_W(14, 73) <= 1; play_W(14, 74) <= 1; play_W(14, 75) <= 0; play_W(14, 76) <= 0; play_W(14, 77) <= 0; play_W(14, 78) <= 0; play_W(14, 79) <= 0; play_W(14, 80) <= 0; play_W(14, 81) <= 0; play_W(14, 82) <= 0; play_W(14, 83) <= 0; play_W(14, 84) <= 0; play_W(14, 85) <= 0; play_W(14, 86) <= 0; play_W(14, 87) <= 1; play_W(14, 88) <= 1; play_W(14, 89) <= 1; play_W(14, 90) <= 1; play_W(14, 91) <= 1; play_W(14, 92) <= 1; play_W(14, 93) <= 1; play_W(14, 94) <= 1; play_W(14, 95) <= 1; play_W(14, 96) <= 1; play_W(14, 97) <= 1; play_W(14, 98) <= 1; play_W(14, 99) <= 0; play_W(14, 100) <= 0; play_W(14, 101) <= 0; play_W(14, 102) <= 0; play_W(14, 103) <= 0; play_W(14, 104) <= 0; play_W(14, 105) <= 0; play_W(14, 106) <= 0; play_W(14, 107) <= 0; play_W(14, 108) <= 0; play_W(14, 109) <= 0; play_W(14, 110) <= 0; play_W(14, 111) <= 0; play_W(14, 112) <= 0; play_W(14, 113) <= 0; play_W(14, 114) <= 0; play_W(14, 115) <= 0; play_W(14, 116) <= 0; play_W(14, 117) <= 0; play_W(14, 118) <= 0; play_W(14, 119) <= 0; play_W(14, 120) <= 0; play_W(14, 121) <= 0; play_W(14, 122) <= 0; play_W(14, 123) <= 0; play_W(14, 124) <= 0; play_W(14, 125) <= 0; play_W(14, 126) <= 0; play_W(14, 127) <= 0; play_W(14, 128) <= 0; play_W(14, 129) <= 0; play_W(14, 130) <= 0; play_W(14, 131) <= 0; play_W(14, 132) <= 0; play_W(14, 133) <= 0; play_W(14, 134) <= 0; play_W(14, 135) <= 0; play_W(14, 136) <= 0; play_W(14, 137) <= 0; play_W(14, 138) <= 0; play_W(14, 139) <= 0; play_W(14, 140) <= 0; play_W(14, 141) <= 0; play_W(14, 142) <= 0; play_W(14, 143) <= 0; play_W(14, 144) <= 0; play_W(14, 145) <= 0; play_W(14, 146) <= 0; play_W(14, 147) <= 0; play_W(14, 148) <= 0; play_W(14, 149) <= 0; play_W(14, 150) <= 0; play_W(14, 151) <= 0; play_W(14, 152) <= 0; play_W(14, 153) <= 0; play_W(14, 154) <= 0; play_W(14, 155) <= 0; play_W(14, 156) <= 0; play_W(14, 157) <= 0; play_W(14, 158) <= 0; play_W(14, 159) <= 0; play_W(14, 160) <= 0; play_W(14, 161) <= 0; play_W(14, 162) <= 0; play_W(14, 163) <= 0; play_W(14, 164) <= 0; play_W(14, 165) <= 1; play_W(14, 166) <= 1; play_W(14, 167) <= 1; play_W(14, 168) <= 1; play_W(14, 169) <= 1; play_W(14, 170) <= 1; play_W(14, 171) <= 1; play_W(14, 172) <= 1; play_W(14, 173) <= 1; play_W(14, 174) <= 1; play_W(14, 175) <= 1; play_W(14, 176) <= 1; play_W(14, 177) <= 1; play_W(14, 178) <= 1; play_W(14, 179) <= 1; play_W(14, 180) <= 0; play_W(14, 181) <= 0; play_W(14, 182) <= 0; play_W(14, 183) <= 0; play_W(14, 184) <= 0; play_W(14, 185) <= 0; play_W(14, 186) <= 0; play_W(14, 187) <= 0; play_W(14, 188) <= 0; play_W(14, 189) <= 0; play_W(14, 190) <= 0; play_W(14, 191) <= 0; play_W(14, 192) <= 0; play_W(14, 193) <= 0; play_W(14, 194) <= 0; play_W(14, 195) <= 0; play_W(14, 196) <= 0; play_W(14, 197) <= 0; play_W(14, 198) <= 1; play_W(14, 199) <= 1; play_W(14, 200) <= 1; play_W(14, 201) <= 1; play_W(14, 202) <= 1; play_W(14, 203) <= 1; play_W(14, 204) <= 0; play_W(14, 205) <= 0; play_W(14, 206) <= 0; play_W(14, 207) <= 0; play_W(14, 208) <= 0; play_W(14, 209) <= 0; play_W(14, 210) <= 0; play_W(14, 211) <= 0; play_W(14, 212) <= 0; play_W(14, 213) <= 0; play_W(14, 214) <= 0; play_W(14, 215) <= 0; play_W(14, 216) <= 1; play_W(14, 217) <= 1; play_W(14, 218) <= 1; play_W(14, 219) <= 1; play_W(14, 220) <= 1; play_W(14, 221) <= 1; play_W(14, 222) <= 0; play_W(14, 223) <= 0; play_W(14, 224) <= 0; play_W(14, 225) <= 1; play_W(14, 226) <= 1; play_W(14, 227) <= 1; play_W(14, 228) <= 1; play_W(14, 229) <= 1; play_W(14, 230) <= 1; play_W(14, 231) <= 1; play_W(14, 232) <= 1; play_W(14, 233) <= 1; play_W(14, 234) <= 1; play_W(14, 235) <= 1; play_W(14, 236) <= 1; play_W(14, 237) <= 0; play_W(14, 238) <= 0; play_W(14, 239) <= 0; play_W(14, 240) <= 0; play_W(14, 241) <= 0; play_W(14, 242) <= 0; play_W(14, 243) <= 0; play_W(14, 244) <= 0; play_W(14, 245) <= 0; play_W(14, 246) <= 1; play_W(14, 247) <= 1; play_W(14, 248) <= 1; play_W(14, 249) <= 1; play_W(14, 250) <= 1; play_W(14, 251) <= 1; play_W(14, 252) <= 1; play_W(14, 253) <= 1; play_W(14, 254) <= 1; play_W(14, 255) <= 1; play_W(14, 256) <= 1; play_W(14, 257) <= 1; play_W(14, 258) <= 1; play_W(14, 259) <= 1; play_W(14, 260) <= 1; play_W(14, 261) <= 0; play_W(14, 262) <= 0; play_W(14, 263) <= 0; play_W(14, 264) <= 0; play_W(14, 265) <= 0; play_W(14, 266) <= 0; play_W(14, 267) <= 0; play_W(14, 268) <= 0; play_W(14, 269) <= 0; 
play_W(15, 0) <= 0; play_W(15, 1) <= 0; play_W(15, 2) <= 0; play_W(15, 3) <= 1; play_W(15, 4) <= 1; play_W(15, 5) <= 1; play_W(15, 6) <= 1; play_W(15, 7) <= 1; play_W(15, 8) <= 1; play_W(15, 9) <= 0; play_W(15, 10) <= 0; play_W(15, 11) <= 0; play_W(15, 12) <= 0; play_W(15, 13) <= 0; play_W(15, 14) <= 0; play_W(15, 15) <= 0; play_W(15, 16) <= 0; play_W(15, 17) <= 0; play_W(15, 18) <= 0; play_W(15, 19) <= 0; play_W(15, 20) <= 0; play_W(15, 21) <= 0; play_W(15, 22) <= 0; play_W(15, 23) <= 0; play_W(15, 24) <= 0; play_W(15, 25) <= 0; play_W(15, 26) <= 0; play_W(15, 27) <= 0; play_W(15, 28) <= 0; play_W(15, 29) <= 0; play_W(15, 30) <= 1; play_W(15, 31) <= 1; play_W(15, 32) <= 1; play_W(15, 33) <= 1; play_W(15, 34) <= 1; play_W(15, 35) <= 1; play_W(15, 36) <= 0; play_W(15, 37) <= 0; play_W(15, 38) <= 0; play_W(15, 39) <= 0; play_W(15, 40) <= 0; play_W(15, 41) <= 0; play_W(15, 42) <= 0; play_W(15, 43) <= 0; play_W(15, 44) <= 0; play_W(15, 45) <= 0; play_W(15, 46) <= 0; play_W(15, 47) <= 0; play_W(15, 48) <= 0; play_W(15, 49) <= 0; play_W(15, 50) <= 0; play_W(15, 51) <= 0; play_W(15, 52) <= 0; play_W(15, 53) <= 0; play_W(15, 54) <= 1; play_W(15, 55) <= 1; play_W(15, 56) <= 1; play_W(15, 57) <= 1; play_W(15, 58) <= 1; play_W(15, 59) <= 1; play_W(15, 60) <= 1; play_W(15, 61) <= 1; play_W(15, 62) <= 1; play_W(15, 63) <= 1; play_W(15, 64) <= 1; play_W(15, 65) <= 1; play_W(15, 66) <= 1; play_W(15, 67) <= 1; play_W(15, 68) <= 1; play_W(15, 69) <= 1; play_W(15, 70) <= 1; play_W(15, 71) <= 1; play_W(15, 72) <= 1; play_W(15, 73) <= 1; play_W(15, 74) <= 1; play_W(15, 75) <= 0; play_W(15, 76) <= 0; play_W(15, 77) <= 0; play_W(15, 78) <= 0; play_W(15, 79) <= 0; play_W(15, 80) <= 0; play_W(15, 81) <= 0; play_W(15, 82) <= 0; play_W(15, 83) <= 0; play_W(15, 84) <= 0; play_W(15, 85) <= 0; play_W(15, 86) <= 0; play_W(15, 87) <= 0; play_W(15, 88) <= 0; play_W(15, 89) <= 0; play_W(15, 90) <= 1; play_W(15, 91) <= 1; play_W(15, 92) <= 1; play_W(15, 93) <= 1; play_W(15, 94) <= 1; play_W(15, 95) <= 1; play_W(15, 96) <= 0; play_W(15, 97) <= 0; play_W(15, 98) <= 0; play_W(15, 99) <= 0; play_W(15, 100) <= 0; play_W(15, 101) <= 0; play_W(15, 102) <= 0; play_W(15, 103) <= 0; play_W(15, 104) <= 0; play_W(15, 105) <= 0; play_W(15, 106) <= 0; play_W(15, 107) <= 0; play_W(15, 108) <= 0; play_W(15, 109) <= 0; play_W(15, 110) <= 0; play_W(15, 111) <= 0; play_W(15, 112) <= 0; play_W(15, 113) <= 0; play_W(15, 114) <= 0; play_W(15, 115) <= 0; play_W(15, 116) <= 0; play_W(15, 117) <= 0; play_W(15, 118) <= 0; play_W(15, 119) <= 0; play_W(15, 120) <= 0; play_W(15, 121) <= 0; play_W(15, 122) <= 0; play_W(15, 123) <= 0; play_W(15, 124) <= 0; play_W(15, 125) <= 0; play_W(15, 126) <= 0; play_W(15, 127) <= 0; play_W(15, 128) <= 0; play_W(15, 129) <= 0; play_W(15, 130) <= 0; play_W(15, 131) <= 0; play_W(15, 132) <= 0; play_W(15, 133) <= 0; play_W(15, 134) <= 0; play_W(15, 135) <= 0; play_W(15, 136) <= 0; play_W(15, 137) <= 0; play_W(15, 138) <= 0; play_W(15, 139) <= 0; play_W(15, 140) <= 0; play_W(15, 141) <= 0; play_W(15, 142) <= 0; play_W(15, 143) <= 0; play_W(15, 144) <= 0; play_W(15, 145) <= 0; play_W(15, 146) <= 0; play_W(15, 147) <= 0; play_W(15, 148) <= 0; play_W(15, 149) <= 0; play_W(15, 150) <= 0; play_W(15, 151) <= 0; play_W(15, 152) <= 0; play_W(15, 153) <= 0; play_W(15, 154) <= 0; play_W(15, 155) <= 0; play_W(15, 156) <= 0; play_W(15, 157) <= 0; play_W(15, 158) <= 0; play_W(15, 159) <= 0; play_W(15, 160) <= 0; play_W(15, 161) <= 0; play_W(15, 162) <= 0; play_W(15, 163) <= 0; play_W(15, 164) <= 0; play_W(15, 165) <= 1; play_W(15, 166) <= 1; play_W(15, 167) <= 1; play_W(15, 168) <= 1; play_W(15, 169) <= 1; play_W(15, 170) <= 1; play_W(15, 171) <= 0; play_W(15, 172) <= 0; play_W(15, 173) <= 0; play_W(15, 174) <= 0; play_W(15, 175) <= 0; play_W(15, 176) <= 0; play_W(15, 177) <= 1; play_W(15, 178) <= 1; play_W(15, 179) <= 1; play_W(15, 180) <= 1; play_W(15, 181) <= 1; play_W(15, 182) <= 1; play_W(15, 183) <= 0; play_W(15, 184) <= 0; play_W(15, 185) <= 0; play_W(15, 186) <= 0; play_W(15, 187) <= 0; play_W(15, 188) <= 0; play_W(15, 189) <= 0; play_W(15, 190) <= 0; play_W(15, 191) <= 0; play_W(15, 192) <= 0; play_W(15, 193) <= 0; play_W(15, 194) <= 0; play_W(15, 195) <= 0; play_W(15, 196) <= 0; play_W(15, 197) <= 0; play_W(15, 198) <= 1; play_W(15, 199) <= 1; play_W(15, 200) <= 1; play_W(15, 201) <= 1; play_W(15, 202) <= 1; play_W(15, 203) <= 1; play_W(15, 204) <= 0; play_W(15, 205) <= 0; play_W(15, 206) <= 0; play_W(15, 207) <= 0; play_W(15, 208) <= 0; play_W(15, 209) <= 0; play_W(15, 210) <= 0; play_W(15, 211) <= 0; play_W(15, 212) <= 0; play_W(15, 213) <= 0; play_W(15, 214) <= 0; play_W(15, 215) <= 0; play_W(15, 216) <= 1; play_W(15, 217) <= 1; play_W(15, 218) <= 1; play_W(15, 219) <= 1; play_W(15, 220) <= 1; play_W(15, 221) <= 1; play_W(15, 222) <= 0; play_W(15, 223) <= 0; play_W(15, 224) <= 0; play_W(15, 225) <= 0; play_W(15, 226) <= 0; play_W(15, 227) <= 0; play_W(15, 228) <= 1; play_W(15, 229) <= 1; play_W(15, 230) <= 1; play_W(15, 231) <= 1; play_W(15, 232) <= 1; play_W(15, 233) <= 1; play_W(15, 234) <= 1; play_W(15, 235) <= 1; play_W(15, 236) <= 1; play_W(15, 237) <= 0; play_W(15, 238) <= 0; play_W(15, 239) <= 0; play_W(15, 240) <= 0; play_W(15, 241) <= 0; play_W(15, 242) <= 0; play_W(15, 243) <= 0; play_W(15, 244) <= 0; play_W(15, 245) <= 0; play_W(15, 246) <= 1; play_W(15, 247) <= 1; play_W(15, 248) <= 1; play_W(15, 249) <= 1; play_W(15, 250) <= 1; play_W(15, 251) <= 1; play_W(15, 252) <= 0; play_W(15, 253) <= 0; play_W(15, 254) <= 0; play_W(15, 255) <= 1; play_W(15, 256) <= 1; play_W(15, 257) <= 1; play_W(15, 258) <= 1; play_W(15, 259) <= 1; play_W(15, 260) <= 1; play_W(15, 261) <= 0; play_W(15, 262) <= 0; play_W(15, 263) <= 0; play_W(15, 264) <= 0; play_W(15, 265) <= 0; play_W(15, 266) <= 0; play_W(15, 267) <= 0; play_W(15, 268) <= 0; play_W(15, 269) <= 0; 
play_W(16, 0) <= 0; play_W(16, 1) <= 0; play_W(16, 2) <= 0; play_W(16, 3) <= 1; play_W(16, 4) <= 1; play_W(16, 5) <= 1; play_W(16, 6) <= 1; play_W(16, 7) <= 1; play_W(16, 8) <= 1; play_W(16, 9) <= 0; play_W(16, 10) <= 0; play_W(16, 11) <= 0; play_W(16, 12) <= 0; play_W(16, 13) <= 0; play_W(16, 14) <= 0; play_W(16, 15) <= 0; play_W(16, 16) <= 0; play_W(16, 17) <= 0; play_W(16, 18) <= 0; play_W(16, 19) <= 0; play_W(16, 20) <= 0; play_W(16, 21) <= 0; play_W(16, 22) <= 0; play_W(16, 23) <= 0; play_W(16, 24) <= 0; play_W(16, 25) <= 0; play_W(16, 26) <= 0; play_W(16, 27) <= 0; play_W(16, 28) <= 0; play_W(16, 29) <= 0; play_W(16, 30) <= 1; play_W(16, 31) <= 1; play_W(16, 32) <= 1; play_W(16, 33) <= 1; play_W(16, 34) <= 1; play_W(16, 35) <= 1; play_W(16, 36) <= 0; play_W(16, 37) <= 0; play_W(16, 38) <= 0; play_W(16, 39) <= 0; play_W(16, 40) <= 0; play_W(16, 41) <= 0; play_W(16, 42) <= 0; play_W(16, 43) <= 0; play_W(16, 44) <= 0; play_W(16, 45) <= 0; play_W(16, 46) <= 0; play_W(16, 47) <= 0; play_W(16, 48) <= 0; play_W(16, 49) <= 0; play_W(16, 50) <= 0; play_W(16, 51) <= 0; play_W(16, 52) <= 0; play_W(16, 53) <= 0; play_W(16, 54) <= 1; play_W(16, 55) <= 1; play_W(16, 56) <= 1; play_W(16, 57) <= 1; play_W(16, 58) <= 1; play_W(16, 59) <= 1; play_W(16, 60) <= 1; play_W(16, 61) <= 1; play_W(16, 62) <= 1; play_W(16, 63) <= 1; play_W(16, 64) <= 1; play_W(16, 65) <= 1; play_W(16, 66) <= 1; play_W(16, 67) <= 1; play_W(16, 68) <= 1; play_W(16, 69) <= 1; play_W(16, 70) <= 1; play_W(16, 71) <= 1; play_W(16, 72) <= 1; play_W(16, 73) <= 1; play_W(16, 74) <= 1; play_W(16, 75) <= 0; play_W(16, 76) <= 0; play_W(16, 77) <= 0; play_W(16, 78) <= 0; play_W(16, 79) <= 0; play_W(16, 80) <= 0; play_W(16, 81) <= 0; play_W(16, 82) <= 0; play_W(16, 83) <= 0; play_W(16, 84) <= 0; play_W(16, 85) <= 0; play_W(16, 86) <= 0; play_W(16, 87) <= 0; play_W(16, 88) <= 0; play_W(16, 89) <= 0; play_W(16, 90) <= 1; play_W(16, 91) <= 1; play_W(16, 92) <= 1; play_W(16, 93) <= 1; play_W(16, 94) <= 1; play_W(16, 95) <= 1; play_W(16, 96) <= 0; play_W(16, 97) <= 0; play_W(16, 98) <= 0; play_W(16, 99) <= 0; play_W(16, 100) <= 0; play_W(16, 101) <= 0; play_W(16, 102) <= 0; play_W(16, 103) <= 0; play_W(16, 104) <= 0; play_W(16, 105) <= 0; play_W(16, 106) <= 0; play_W(16, 107) <= 0; play_W(16, 108) <= 0; play_W(16, 109) <= 0; play_W(16, 110) <= 0; play_W(16, 111) <= 0; play_W(16, 112) <= 0; play_W(16, 113) <= 0; play_W(16, 114) <= 0; play_W(16, 115) <= 0; play_W(16, 116) <= 0; play_W(16, 117) <= 0; play_W(16, 118) <= 0; play_W(16, 119) <= 0; play_W(16, 120) <= 0; play_W(16, 121) <= 0; play_W(16, 122) <= 0; play_W(16, 123) <= 0; play_W(16, 124) <= 0; play_W(16, 125) <= 0; play_W(16, 126) <= 0; play_W(16, 127) <= 0; play_W(16, 128) <= 0; play_W(16, 129) <= 0; play_W(16, 130) <= 0; play_W(16, 131) <= 0; play_W(16, 132) <= 0; play_W(16, 133) <= 0; play_W(16, 134) <= 0; play_W(16, 135) <= 0; play_W(16, 136) <= 0; play_W(16, 137) <= 0; play_W(16, 138) <= 0; play_W(16, 139) <= 0; play_W(16, 140) <= 0; play_W(16, 141) <= 0; play_W(16, 142) <= 0; play_W(16, 143) <= 0; play_W(16, 144) <= 0; play_W(16, 145) <= 0; play_W(16, 146) <= 0; play_W(16, 147) <= 0; play_W(16, 148) <= 0; play_W(16, 149) <= 0; play_W(16, 150) <= 0; play_W(16, 151) <= 0; play_W(16, 152) <= 0; play_W(16, 153) <= 0; play_W(16, 154) <= 0; play_W(16, 155) <= 0; play_W(16, 156) <= 0; play_W(16, 157) <= 0; play_W(16, 158) <= 0; play_W(16, 159) <= 0; play_W(16, 160) <= 0; play_W(16, 161) <= 0; play_W(16, 162) <= 0; play_W(16, 163) <= 0; play_W(16, 164) <= 0; play_W(16, 165) <= 1; play_W(16, 166) <= 1; play_W(16, 167) <= 1; play_W(16, 168) <= 1; play_W(16, 169) <= 1; play_W(16, 170) <= 1; play_W(16, 171) <= 0; play_W(16, 172) <= 0; play_W(16, 173) <= 0; play_W(16, 174) <= 0; play_W(16, 175) <= 0; play_W(16, 176) <= 0; play_W(16, 177) <= 1; play_W(16, 178) <= 1; play_W(16, 179) <= 1; play_W(16, 180) <= 1; play_W(16, 181) <= 1; play_W(16, 182) <= 1; play_W(16, 183) <= 0; play_W(16, 184) <= 0; play_W(16, 185) <= 0; play_W(16, 186) <= 0; play_W(16, 187) <= 0; play_W(16, 188) <= 0; play_W(16, 189) <= 0; play_W(16, 190) <= 0; play_W(16, 191) <= 0; play_W(16, 192) <= 0; play_W(16, 193) <= 0; play_W(16, 194) <= 0; play_W(16, 195) <= 0; play_W(16, 196) <= 0; play_W(16, 197) <= 0; play_W(16, 198) <= 1; play_W(16, 199) <= 1; play_W(16, 200) <= 1; play_W(16, 201) <= 1; play_W(16, 202) <= 1; play_W(16, 203) <= 1; play_W(16, 204) <= 0; play_W(16, 205) <= 0; play_W(16, 206) <= 0; play_W(16, 207) <= 0; play_W(16, 208) <= 0; play_W(16, 209) <= 0; play_W(16, 210) <= 0; play_W(16, 211) <= 0; play_W(16, 212) <= 0; play_W(16, 213) <= 0; play_W(16, 214) <= 0; play_W(16, 215) <= 0; play_W(16, 216) <= 1; play_W(16, 217) <= 1; play_W(16, 218) <= 1; play_W(16, 219) <= 1; play_W(16, 220) <= 1; play_W(16, 221) <= 1; play_W(16, 222) <= 0; play_W(16, 223) <= 0; play_W(16, 224) <= 0; play_W(16, 225) <= 0; play_W(16, 226) <= 0; play_W(16, 227) <= 0; play_W(16, 228) <= 1; play_W(16, 229) <= 1; play_W(16, 230) <= 1; play_W(16, 231) <= 1; play_W(16, 232) <= 1; play_W(16, 233) <= 1; play_W(16, 234) <= 1; play_W(16, 235) <= 1; play_W(16, 236) <= 1; play_W(16, 237) <= 0; play_W(16, 238) <= 0; play_W(16, 239) <= 0; play_W(16, 240) <= 0; play_W(16, 241) <= 0; play_W(16, 242) <= 0; play_W(16, 243) <= 0; play_W(16, 244) <= 0; play_W(16, 245) <= 0; play_W(16, 246) <= 1; play_W(16, 247) <= 1; play_W(16, 248) <= 1; play_W(16, 249) <= 1; play_W(16, 250) <= 1; play_W(16, 251) <= 1; play_W(16, 252) <= 0; play_W(16, 253) <= 0; play_W(16, 254) <= 0; play_W(16, 255) <= 1; play_W(16, 256) <= 1; play_W(16, 257) <= 1; play_W(16, 258) <= 1; play_W(16, 259) <= 1; play_W(16, 260) <= 1; play_W(16, 261) <= 0; play_W(16, 262) <= 0; play_W(16, 263) <= 0; play_W(16, 264) <= 0; play_W(16, 265) <= 0; play_W(16, 266) <= 0; play_W(16, 267) <= 0; play_W(16, 268) <= 0; play_W(16, 269) <= 0; 
play_W(17, 0) <= 0; play_W(17, 1) <= 0; play_W(17, 2) <= 0; play_W(17, 3) <= 1; play_W(17, 4) <= 1; play_W(17, 5) <= 1; play_W(17, 6) <= 1; play_W(17, 7) <= 1; play_W(17, 8) <= 1; play_W(17, 9) <= 0; play_W(17, 10) <= 0; play_W(17, 11) <= 0; play_W(17, 12) <= 0; play_W(17, 13) <= 0; play_W(17, 14) <= 0; play_W(17, 15) <= 0; play_W(17, 16) <= 0; play_W(17, 17) <= 0; play_W(17, 18) <= 0; play_W(17, 19) <= 0; play_W(17, 20) <= 0; play_W(17, 21) <= 0; play_W(17, 22) <= 0; play_W(17, 23) <= 0; play_W(17, 24) <= 0; play_W(17, 25) <= 0; play_W(17, 26) <= 0; play_W(17, 27) <= 0; play_W(17, 28) <= 0; play_W(17, 29) <= 0; play_W(17, 30) <= 1; play_W(17, 31) <= 1; play_W(17, 32) <= 1; play_W(17, 33) <= 1; play_W(17, 34) <= 1; play_W(17, 35) <= 1; play_W(17, 36) <= 0; play_W(17, 37) <= 0; play_W(17, 38) <= 0; play_W(17, 39) <= 0; play_W(17, 40) <= 0; play_W(17, 41) <= 0; play_W(17, 42) <= 0; play_W(17, 43) <= 0; play_W(17, 44) <= 0; play_W(17, 45) <= 0; play_W(17, 46) <= 0; play_W(17, 47) <= 0; play_W(17, 48) <= 0; play_W(17, 49) <= 0; play_W(17, 50) <= 0; play_W(17, 51) <= 0; play_W(17, 52) <= 0; play_W(17, 53) <= 0; play_W(17, 54) <= 1; play_W(17, 55) <= 1; play_W(17, 56) <= 1; play_W(17, 57) <= 1; play_W(17, 58) <= 1; play_W(17, 59) <= 1; play_W(17, 60) <= 1; play_W(17, 61) <= 1; play_W(17, 62) <= 1; play_W(17, 63) <= 1; play_W(17, 64) <= 1; play_W(17, 65) <= 1; play_W(17, 66) <= 1; play_W(17, 67) <= 1; play_W(17, 68) <= 1; play_W(17, 69) <= 1; play_W(17, 70) <= 1; play_W(17, 71) <= 1; play_W(17, 72) <= 1; play_W(17, 73) <= 1; play_W(17, 74) <= 1; play_W(17, 75) <= 0; play_W(17, 76) <= 0; play_W(17, 77) <= 0; play_W(17, 78) <= 0; play_W(17, 79) <= 0; play_W(17, 80) <= 0; play_W(17, 81) <= 0; play_W(17, 82) <= 0; play_W(17, 83) <= 0; play_W(17, 84) <= 0; play_W(17, 85) <= 0; play_W(17, 86) <= 0; play_W(17, 87) <= 0; play_W(17, 88) <= 0; play_W(17, 89) <= 0; play_W(17, 90) <= 1; play_W(17, 91) <= 1; play_W(17, 92) <= 1; play_W(17, 93) <= 1; play_W(17, 94) <= 1; play_W(17, 95) <= 1; play_W(17, 96) <= 0; play_W(17, 97) <= 0; play_W(17, 98) <= 0; play_W(17, 99) <= 0; play_W(17, 100) <= 0; play_W(17, 101) <= 0; play_W(17, 102) <= 0; play_W(17, 103) <= 0; play_W(17, 104) <= 0; play_W(17, 105) <= 0; play_W(17, 106) <= 0; play_W(17, 107) <= 0; play_W(17, 108) <= 0; play_W(17, 109) <= 0; play_W(17, 110) <= 0; play_W(17, 111) <= 0; play_W(17, 112) <= 0; play_W(17, 113) <= 0; play_W(17, 114) <= 0; play_W(17, 115) <= 0; play_W(17, 116) <= 0; play_W(17, 117) <= 0; play_W(17, 118) <= 0; play_W(17, 119) <= 0; play_W(17, 120) <= 0; play_W(17, 121) <= 0; play_W(17, 122) <= 0; play_W(17, 123) <= 0; play_W(17, 124) <= 0; play_W(17, 125) <= 0; play_W(17, 126) <= 0; play_W(17, 127) <= 0; play_W(17, 128) <= 0; play_W(17, 129) <= 0; play_W(17, 130) <= 0; play_W(17, 131) <= 0; play_W(17, 132) <= 0; play_W(17, 133) <= 0; play_W(17, 134) <= 0; play_W(17, 135) <= 0; play_W(17, 136) <= 0; play_W(17, 137) <= 0; play_W(17, 138) <= 0; play_W(17, 139) <= 0; play_W(17, 140) <= 0; play_W(17, 141) <= 0; play_W(17, 142) <= 0; play_W(17, 143) <= 0; play_W(17, 144) <= 0; play_W(17, 145) <= 0; play_W(17, 146) <= 0; play_W(17, 147) <= 0; play_W(17, 148) <= 0; play_W(17, 149) <= 0; play_W(17, 150) <= 0; play_W(17, 151) <= 0; play_W(17, 152) <= 0; play_W(17, 153) <= 0; play_W(17, 154) <= 0; play_W(17, 155) <= 0; play_W(17, 156) <= 0; play_W(17, 157) <= 0; play_W(17, 158) <= 0; play_W(17, 159) <= 0; play_W(17, 160) <= 0; play_W(17, 161) <= 0; play_W(17, 162) <= 0; play_W(17, 163) <= 0; play_W(17, 164) <= 0; play_W(17, 165) <= 1; play_W(17, 166) <= 1; play_W(17, 167) <= 1; play_W(17, 168) <= 1; play_W(17, 169) <= 1; play_W(17, 170) <= 1; play_W(17, 171) <= 0; play_W(17, 172) <= 0; play_W(17, 173) <= 0; play_W(17, 174) <= 0; play_W(17, 175) <= 0; play_W(17, 176) <= 0; play_W(17, 177) <= 1; play_W(17, 178) <= 1; play_W(17, 179) <= 1; play_W(17, 180) <= 1; play_W(17, 181) <= 1; play_W(17, 182) <= 1; play_W(17, 183) <= 0; play_W(17, 184) <= 0; play_W(17, 185) <= 0; play_W(17, 186) <= 0; play_W(17, 187) <= 0; play_W(17, 188) <= 0; play_W(17, 189) <= 0; play_W(17, 190) <= 0; play_W(17, 191) <= 0; play_W(17, 192) <= 0; play_W(17, 193) <= 0; play_W(17, 194) <= 0; play_W(17, 195) <= 0; play_W(17, 196) <= 0; play_W(17, 197) <= 0; play_W(17, 198) <= 1; play_W(17, 199) <= 1; play_W(17, 200) <= 1; play_W(17, 201) <= 1; play_W(17, 202) <= 1; play_W(17, 203) <= 1; play_W(17, 204) <= 0; play_W(17, 205) <= 0; play_W(17, 206) <= 0; play_W(17, 207) <= 0; play_W(17, 208) <= 0; play_W(17, 209) <= 0; play_W(17, 210) <= 0; play_W(17, 211) <= 0; play_W(17, 212) <= 0; play_W(17, 213) <= 0; play_W(17, 214) <= 0; play_W(17, 215) <= 0; play_W(17, 216) <= 1; play_W(17, 217) <= 1; play_W(17, 218) <= 1; play_W(17, 219) <= 1; play_W(17, 220) <= 1; play_W(17, 221) <= 1; play_W(17, 222) <= 0; play_W(17, 223) <= 0; play_W(17, 224) <= 0; play_W(17, 225) <= 0; play_W(17, 226) <= 0; play_W(17, 227) <= 0; play_W(17, 228) <= 1; play_W(17, 229) <= 1; play_W(17, 230) <= 1; play_W(17, 231) <= 1; play_W(17, 232) <= 1; play_W(17, 233) <= 1; play_W(17, 234) <= 1; play_W(17, 235) <= 1; play_W(17, 236) <= 1; play_W(17, 237) <= 0; play_W(17, 238) <= 0; play_W(17, 239) <= 0; play_W(17, 240) <= 0; play_W(17, 241) <= 0; play_W(17, 242) <= 0; play_W(17, 243) <= 0; play_W(17, 244) <= 0; play_W(17, 245) <= 0; play_W(17, 246) <= 1; play_W(17, 247) <= 1; play_W(17, 248) <= 1; play_W(17, 249) <= 1; play_W(17, 250) <= 1; play_W(17, 251) <= 1; play_W(17, 252) <= 0; play_W(17, 253) <= 0; play_W(17, 254) <= 0; play_W(17, 255) <= 1; play_W(17, 256) <= 1; play_W(17, 257) <= 1; play_W(17, 258) <= 1; play_W(17, 259) <= 1; play_W(17, 260) <= 1; play_W(17, 261) <= 0; play_W(17, 262) <= 0; play_W(17, 263) <= 0; play_W(17, 264) <= 0; play_W(17, 265) <= 0; play_W(17, 266) <= 0; play_W(17, 267) <= 0; play_W(17, 268) <= 0; play_W(17, 269) <= 0; 
play_W(18, 0) <= 0; play_W(18, 1) <= 0; play_W(18, 2) <= 0; play_W(18, 3) <= 1; play_W(18, 4) <= 1; play_W(18, 5) <= 1; play_W(18, 6) <= 1; play_W(18, 7) <= 1; play_W(18, 8) <= 1; play_W(18, 9) <= 0; play_W(18, 10) <= 0; play_W(18, 11) <= 0; play_W(18, 12) <= 0; play_W(18, 13) <= 0; play_W(18, 14) <= 0; play_W(18, 15) <= 0; play_W(18, 16) <= 0; play_W(18, 17) <= 0; play_W(18, 18) <= 0; play_W(18, 19) <= 0; play_W(18, 20) <= 0; play_W(18, 21) <= 0; play_W(18, 22) <= 0; play_W(18, 23) <= 0; play_W(18, 24) <= 0; play_W(18, 25) <= 0; play_W(18, 26) <= 0; play_W(18, 27) <= 0; play_W(18, 28) <= 0; play_W(18, 29) <= 0; play_W(18, 30) <= 1; play_W(18, 31) <= 1; play_W(18, 32) <= 1; play_W(18, 33) <= 1; play_W(18, 34) <= 1; play_W(18, 35) <= 1; play_W(18, 36) <= 0; play_W(18, 37) <= 0; play_W(18, 38) <= 0; play_W(18, 39) <= 0; play_W(18, 40) <= 0; play_W(18, 41) <= 0; play_W(18, 42) <= 0; play_W(18, 43) <= 0; play_W(18, 44) <= 0; play_W(18, 45) <= 0; play_W(18, 46) <= 0; play_W(18, 47) <= 0; play_W(18, 48) <= 0; play_W(18, 49) <= 0; play_W(18, 50) <= 0; play_W(18, 51) <= 0; play_W(18, 52) <= 0; play_W(18, 53) <= 0; play_W(18, 54) <= 1; play_W(18, 55) <= 1; play_W(18, 56) <= 1; play_W(18, 57) <= 1; play_W(18, 58) <= 1; play_W(18, 59) <= 1; play_W(18, 60) <= 0; play_W(18, 61) <= 0; play_W(18, 62) <= 0; play_W(18, 63) <= 0; play_W(18, 64) <= 0; play_W(18, 65) <= 0; play_W(18, 66) <= 0; play_W(18, 67) <= 0; play_W(18, 68) <= 0; play_W(18, 69) <= 1; play_W(18, 70) <= 1; play_W(18, 71) <= 1; play_W(18, 72) <= 1; play_W(18, 73) <= 1; play_W(18, 74) <= 1; play_W(18, 75) <= 0; play_W(18, 76) <= 0; play_W(18, 77) <= 0; play_W(18, 78) <= 0; play_W(18, 79) <= 0; play_W(18, 80) <= 0; play_W(18, 81) <= 0; play_W(18, 82) <= 0; play_W(18, 83) <= 0; play_W(18, 84) <= 0; play_W(18, 85) <= 0; play_W(18, 86) <= 0; play_W(18, 87) <= 0; play_W(18, 88) <= 0; play_W(18, 89) <= 0; play_W(18, 90) <= 1; play_W(18, 91) <= 1; play_W(18, 92) <= 1; play_W(18, 93) <= 1; play_W(18, 94) <= 1; play_W(18, 95) <= 1; play_W(18, 96) <= 0; play_W(18, 97) <= 0; play_W(18, 98) <= 0; play_W(18, 99) <= 0; play_W(18, 100) <= 0; play_W(18, 101) <= 0; play_W(18, 102) <= 0; play_W(18, 103) <= 0; play_W(18, 104) <= 0; play_W(18, 105) <= 0; play_W(18, 106) <= 0; play_W(18, 107) <= 0; play_W(18, 108) <= 0; play_W(18, 109) <= 0; play_W(18, 110) <= 0; play_W(18, 111) <= 0; play_W(18, 112) <= 0; play_W(18, 113) <= 0; play_W(18, 114) <= 0; play_W(18, 115) <= 0; play_W(18, 116) <= 0; play_W(18, 117) <= 1; play_W(18, 118) <= 1; play_W(18, 119) <= 1; play_W(18, 120) <= 1; play_W(18, 121) <= 1; play_W(18, 122) <= 1; play_W(18, 123) <= 0; play_W(18, 124) <= 0; play_W(18, 125) <= 0; play_W(18, 126) <= 0; play_W(18, 127) <= 0; play_W(18, 128) <= 0; play_W(18, 129) <= 0; play_W(18, 130) <= 0; play_W(18, 131) <= 0; play_W(18, 132) <= 0; play_W(18, 133) <= 0; play_W(18, 134) <= 0; play_W(18, 135) <= 0; play_W(18, 136) <= 0; play_W(18, 137) <= 0; play_W(18, 138) <= 0; play_W(18, 139) <= 0; play_W(18, 140) <= 0; play_W(18, 141) <= 0; play_W(18, 142) <= 0; play_W(18, 143) <= 0; play_W(18, 144) <= 0; play_W(18, 145) <= 0; play_W(18, 146) <= 0; play_W(18, 147) <= 0; play_W(18, 148) <= 0; play_W(18, 149) <= 0; play_W(18, 150) <= 0; play_W(18, 151) <= 0; play_W(18, 152) <= 0; play_W(18, 153) <= 0; play_W(18, 154) <= 0; play_W(18, 155) <= 0; play_W(18, 156) <= 0; play_W(18, 157) <= 0; play_W(18, 158) <= 0; play_W(18, 159) <= 0; play_W(18, 160) <= 0; play_W(18, 161) <= 0; play_W(18, 162) <= 0; play_W(18, 163) <= 0; play_W(18, 164) <= 0; play_W(18, 165) <= 1; play_W(18, 166) <= 1; play_W(18, 167) <= 1; play_W(18, 168) <= 1; play_W(18, 169) <= 1; play_W(18, 170) <= 1; play_W(18, 171) <= 0; play_W(18, 172) <= 0; play_W(18, 173) <= 0; play_W(18, 174) <= 0; play_W(18, 175) <= 0; play_W(18, 176) <= 0; play_W(18, 177) <= 1; play_W(18, 178) <= 1; play_W(18, 179) <= 1; play_W(18, 180) <= 1; play_W(18, 181) <= 1; play_W(18, 182) <= 1; play_W(18, 183) <= 0; play_W(18, 184) <= 0; play_W(18, 185) <= 0; play_W(18, 186) <= 0; play_W(18, 187) <= 0; play_W(18, 188) <= 0; play_W(18, 189) <= 0; play_W(18, 190) <= 0; play_W(18, 191) <= 0; play_W(18, 192) <= 0; play_W(18, 193) <= 0; play_W(18, 194) <= 0; play_W(18, 195) <= 0; play_W(18, 196) <= 0; play_W(18, 197) <= 0; play_W(18, 198) <= 1; play_W(18, 199) <= 1; play_W(18, 200) <= 1; play_W(18, 201) <= 1; play_W(18, 202) <= 1; play_W(18, 203) <= 1; play_W(18, 204) <= 0; play_W(18, 205) <= 0; play_W(18, 206) <= 0; play_W(18, 207) <= 0; play_W(18, 208) <= 0; play_W(18, 209) <= 0; play_W(18, 210) <= 0; play_W(18, 211) <= 0; play_W(18, 212) <= 0; play_W(18, 213) <= 0; play_W(18, 214) <= 0; play_W(18, 215) <= 0; play_W(18, 216) <= 1; play_W(18, 217) <= 1; play_W(18, 218) <= 1; play_W(18, 219) <= 1; play_W(18, 220) <= 1; play_W(18, 221) <= 1; play_W(18, 222) <= 0; play_W(18, 223) <= 0; play_W(18, 224) <= 0; play_W(18, 225) <= 0; play_W(18, 226) <= 0; play_W(18, 227) <= 0; play_W(18, 228) <= 0; play_W(18, 229) <= 0; play_W(18, 230) <= 0; play_W(18, 231) <= 1; play_W(18, 232) <= 1; play_W(18, 233) <= 1; play_W(18, 234) <= 1; play_W(18, 235) <= 1; play_W(18, 236) <= 1; play_W(18, 237) <= 0; play_W(18, 238) <= 0; play_W(18, 239) <= 0; play_W(18, 240) <= 0; play_W(18, 241) <= 0; play_W(18, 242) <= 0; play_W(18, 243) <= 0; play_W(18, 244) <= 0; play_W(18, 245) <= 0; play_W(18, 246) <= 1; play_W(18, 247) <= 1; play_W(18, 248) <= 1; play_W(18, 249) <= 1; play_W(18, 250) <= 1; play_W(18, 251) <= 1; play_W(18, 252) <= 0; play_W(18, 253) <= 0; play_W(18, 254) <= 0; play_W(18, 255) <= 0; play_W(18, 256) <= 0; play_W(18, 257) <= 0; play_W(18, 258) <= 1; play_W(18, 259) <= 1; play_W(18, 260) <= 1; play_W(18, 261) <= 1; play_W(18, 262) <= 1; play_W(18, 263) <= 1; play_W(18, 264) <= 0; play_W(18, 265) <= 0; play_W(18, 266) <= 0; play_W(18, 267) <= 0; play_W(18, 268) <= 0; play_W(18, 269) <= 0; 
play_W(19, 0) <= 0; play_W(19, 1) <= 0; play_W(19, 2) <= 0; play_W(19, 3) <= 1; play_W(19, 4) <= 1; play_W(19, 5) <= 1; play_W(19, 6) <= 1; play_W(19, 7) <= 1; play_W(19, 8) <= 1; play_W(19, 9) <= 0; play_W(19, 10) <= 0; play_W(19, 11) <= 0; play_W(19, 12) <= 0; play_W(19, 13) <= 0; play_W(19, 14) <= 0; play_W(19, 15) <= 0; play_W(19, 16) <= 0; play_W(19, 17) <= 0; play_W(19, 18) <= 0; play_W(19, 19) <= 0; play_W(19, 20) <= 0; play_W(19, 21) <= 0; play_W(19, 22) <= 0; play_W(19, 23) <= 0; play_W(19, 24) <= 0; play_W(19, 25) <= 0; play_W(19, 26) <= 0; play_W(19, 27) <= 0; play_W(19, 28) <= 0; play_W(19, 29) <= 0; play_W(19, 30) <= 1; play_W(19, 31) <= 1; play_W(19, 32) <= 1; play_W(19, 33) <= 1; play_W(19, 34) <= 1; play_W(19, 35) <= 1; play_W(19, 36) <= 0; play_W(19, 37) <= 0; play_W(19, 38) <= 0; play_W(19, 39) <= 0; play_W(19, 40) <= 0; play_W(19, 41) <= 0; play_W(19, 42) <= 0; play_W(19, 43) <= 0; play_W(19, 44) <= 0; play_W(19, 45) <= 0; play_W(19, 46) <= 0; play_W(19, 47) <= 0; play_W(19, 48) <= 0; play_W(19, 49) <= 0; play_W(19, 50) <= 0; play_W(19, 51) <= 0; play_W(19, 52) <= 0; play_W(19, 53) <= 0; play_W(19, 54) <= 1; play_W(19, 55) <= 1; play_W(19, 56) <= 1; play_W(19, 57) <= 1; play_W(19, 58) <= 1; play_W(19, 59) <= 1; play_W(19, 60) <= 0; play_W(19, 61) <= 0; play_W(19, 62) <= 0; play_W(19, 63) <= 0; play_W(19, 64) <= 0; play_W(19, 65) <= 0; play_W(19, 66) <= 0; play_W(19, 67) <= 0; play_W(19, 68) <= 0; play_W(19, 69) <= 1; play_W(19, 70) <= 1; play_W(19, 71) <= 1; play_W(19, 72) <= 1; play_W(19, 73) <= 1; play_W(19, 74) <= 1; play_W(19, 75) <= 0; play_W(19, 76) <= 0; play_W(19, 77) <= 0; play_W(19, 78) <= 0; play_W(19, 79) <= 0; play_W(19, 80) <= 0; play_W(19, 81) <= 0; play_W(19, 82) <= 0; play_W(19, 83) <= 0; play_W(19, 84) <= 0; play_W(19, 85) <= 0; play_W(19, 86) <= 0; play_W(19, 87) <= 0; play_W(19, 88) <= 0; play_W(19, 89) <= 0; play_W(19, 90) <= 1; play_W(19, 91) <= 1; play_W(19, 92) <= 1; play_W(19, 93) <= 1; play_W(19, 94) <= 1; play_W(19, 95) <= 1; play_W(19, 96) <= 0; play_W(19, 97) <= 0; play_W(19, 98) <= 0; play_W(19, 99) <= 0; play_W(19, 100) <= 0; play_W(19, 101) <= 0; play_W(19, 102) <= 0; play_W(19, 103) <= 0; play_W(19, 104) <= 0; play_W(19, 105) <= 0; play_W(19, 106) <= 0; play_W(19, 107) <= 0; play_W(19, 108) <= 0; play_W(19, 109) <= 0; play_W(19, 110) <= 0; play_W(19, 111) <= 0; play_W(19, 112) <= 0; play_W(19, 113) <= 0; play_W(19, 114) <= 0; play_W(19, 115) <= 0; play_W(19, 116) <= 0; play_W(19, 117) <= 1; play_W(19, 118) <= 1; play_W(19, 119) <= 1; play_W(19, 120) <= 1; play_W(19, 121) <= 1; play_W(19, 122) <= 1; play_W(19, 123) <= 0; play_W(19, 124) <= 0; play_W(19, 125) <= 0; play_W(19, 126) <= 0; play_W(19, 127) <= 0; play_W(19, 128) <= 0; play_W(19, 129) <= 0; play_W(19, 130) <= 0; play_W(19, 131) <= 0; play_W(19, 132) <= 0; play_W(19, 133) <= 0; play_W(19, 134) <= 0; play_W(19, 135) <= 0; play_W(19, 136) <= 0; play_W(19, 137) <= 0; play_W(19, 138) <= 0; play_W(19, 139) <= 0; play_W(19, 140) <= 0; play_W(19, 141) <= 0; play_W(19, 142) <= 0; play_W(19, 143) <= 0; play_W(19, 144) <= 0; play_W(19, 145) <= 0; play_W(19, 146) <= 0; play_W(19, 147) <= 0; play_W(19, 148) <= 0; play_W(19, 149) <= 0; play_W(19, 150) <= 0; play_W(19, 151) <= 0; play_W(19, 152) <= 0; play_W(19, 153) <= 0; play_W(19, 154) <= 0; play_W(19, 155) <= 0; play_W(19, 156) <= 0; play_W(19, 157) <= 0; play_W(19, 158) <= 0; play_W(19, 159) <= 0; play_W(19, 160) <= 0; play_W(19, 161) <= 0; play_W(19, 162) <= 0; play_W(19, 163) <= 0; play_W(19, 164) <= 0; play_W(19, 165) <= 1; play_W(19, 166) <= 1; play_W(19, 167) <= 1; play_W(19, 168) <= 1; play_W(19, 169) <= 1; play_W(19, 170) <= 1; play_W(19, 171) <= 0; play_W(19, 172) <= 0; play_W(19, 173) <= 0; play_W(19, 174) <= 0; play_W(19, 175) <= 0; play_W(19, 176) <= 0; play_W(19, 177) <= 1; play_W(19, 178) <= 1; play_W(19, 179) <= 1; play_W(19, 180) <= 1; play_W(19, 181) <= 1; play_W(19, 182) <= 1; play_W(19, 183) <= 0; play_W(19, 184) <= 0; play_W(19, 185) <= 0; play_W(19, 186) <= 0; play_W(19, 187) <= 0; play_W(19, 188) <= 0; play_W(19, 189) <= 0; play_W(19, 190) <= 0; play_W(19, 191) <= 0; play_W(19, 192) <= 0; play_W(19, 193) <= 0; play_W(19, 194) <= 0; play_W(19, 195) <= 0; play_W(19, 196) <= 0; play_W(19, 197) <= 0; play_W(19, 198) <= 1; play_W(19, 199) <= 1; play_W(19, 200) <= 1; play_W(19, 201) <= 1; play_W(19, 202) <= 1; play_W(19, 203) <= 1; play_W(19, 204) <= 0; play_W(19, 205) <= 0; play_W(19, 206) <= 0; play_W(19, 207) <= 0; play_W(19, 208) <= 0; play_W(19, 209) <= 0; play_W(19, 210) <= 0; play_W(19, 211) <= 0; play_W(19, 212) <= 0; play_W(19, 213) <= 0; play_W(19, 214) <= 0; play_W(19, 215) <= 0; play_W(19, 216) <= 1; play_W(19, 217) <= 1; play_W(19, 218) <= 1; play_W(19, 219) <= 1; play_W(19, 220) <= 1; play_W(19, 221) <= 1; play_W(19, 222) <= 0; play_W(19, 223) <= 0; play_W(19, 224) <= 0; play_W(19, 225) <= 0; play_W(19, 226) <= 0; play_W(19, 227) <= 0; play_W(19, 228) <= 0; play_W(19, 229) <= 0; play_W(19, 230) <= 0; play_W(19, 231) <= 1; play_W(19, 232) <= 1; play_W(19, 233) <= 1; play_W(19, 234) <= 1; play_W(19, 235) <= 1; play_W(19, 236) <= 1; play_W(19, 237) <= 0; play_W(19, 238) <= 0; play_W(19, 239) <= 0; play_W(19, 240) <= 0; play_W(19, 241) <= 0; play_W(19, 242) <= 0; play_W(19, 243) <= 0; play_W(19, 244) <= 0; play_W(19, 245) <= 0; play_W(19, 246) <= 1; play_W(19, 247) <= 1; play_W(19, 248) <= 1; play_W(19, 249) <= 1; play_W(19, 250) <= 1; play_W(19, 251) <= 1; play_W(19, 252) <= 0; play_W(19, 253) <= 0; play_W(19, 254) <= 0; play_W(19, 255) <= 0; play_W(19, 256) <= 0; play_W(19, 257) <= 0; play_W(19, 258) <= 1; play_W(19, 259) <= 1; play_W(19, 260) <= 1; play_W(19, 261) <= 1; play_W(19, 262) <= 1; play_W(19, 263) <= 1; play_W(19, 264) <= 0; play_W(19, 265) <= 0; play_W(19, 266) <= 0; play_W(19, 267) <= 0; play_W(19, 268) <= 0; play_W(19, 269) <= 0; 
play_W(20, 0) <= 0; play_W(20, 1) <= 0; play_W(20, 2) <= 0; play_W(20, 3) <= 1; play_W(20, 4) <= 1; play_W(20, 5) <= 1; play_W(20, 6) <= 1; play_W(20, 7) <= 1; play_W(20, 8) <= 1; play_W(20, 9) <= 0; play_W(20, 10) <= 0; play_W(20, 11) <= 0; play_W(20, 12) <= 0; play_W(20, 13) <= 0; play_W(20, 14) <= 0; play_W(20, 15) <= 0; play_W(20, 16) <= 0; play_W(20, 17) <= 0; play_W(20, 18) <= 0; play_W(20, 19) <= 0; play_W(20, 20) <= 0; play_W(20, 21) <= 0; play_W(20, 22) <= 0; play_W(20, 23) <= 0; play_W(20, 24) <= 0; play_W(20, 25) <= 0; play_W(20, 26) <= 0; play_W(20, 27) <= 0; play_W(20, 28) <= 0; play_W(20, 29) <= 0; play_W(20, 30) <= 1; play_W(20, 31) <= 1; play_W(20, 32) <= 1; play_W(20, 33) <= 1; play_W(20, 34) <= 1; play_W(20, 35) <= 1; play_W(20, 36) <= 0; play_W(20, 37) <= 0; play_W(20, 38) <= 0; play_W(20, 39) <= 0; play_W(20, 40) <= 0; play_W(20, 41) <= 0; play_W(20, 42) <= 0; play_W(20, 43) <= 0; play_W(20, 44) <= 0; play_W(20, 45) <= 0; play_W(20, 46) <= 0; play_W(20, 47) <= 0; play_W(20, 48) <= 0; play_W(20, 49) <= 0; play_W(20, 50) <= 0; play_W(20, 51) <= 0; play_W(20, 52) <= 0; play_W(20, 53) <= 0; play_W(20, 54) <= 1; play_W(20, 55) <= 1; play_W(20, 56) <= 1; play_W(20, 57) <= 1; play_W(20, 58) <= 1; play_W(20, 59) <= 1; play_W(20, 60) <= 0; play_W(20, 61) <= 0; play_W(20, 62) <= 0; play_W(20, 63) <= 0; play_W(20, 64) <= 0; play_W(20, 65) <= 0; play_W(20, 66) <= 0; play_W(20, 67) <= 0; play_W(20, 68) <= 0; play_W(20, 69) <= 1; play_W(20, 70) <= 1; play_W(20, 71) <= 1; play_W(20, 72) <= 1; play_W(20, 73) <= 1; play_W(20, 74) <= 1; play_W(20, 75) <= 0; play_W(20, 76) <= 0; play_W(20, 77) <= 0; play_W(20, 78) <= 0; play_W(20, 79) <= 0; play_W(20, 80) <= 0; play_W(20, 81) <= 0; play_W(20, 82) <= 0; play_W(20, 83) <= 0; play_W(20, 84) <= 0; play_W(20, 85) <= 0; play_W(20, 86) <= 0; play_W(20, 87) <= 0; play_W(20, 88) <= 0; play_W(20, 89) <= 0; play_W(20, 90) <= 1; play_W(20, 91) <= 1; play_W(20, 92) <= 1; play_W(20, 93) <= 1; play_W(20, 94) <= 1; play_W(20, 95) <= 1; play_W(20, 96) <= 0; play_W(20, 97) <= 0; play_W(20, 98) <= 0; play_W(20, 99) <= 0; play_W(20, 100) <= 0; play_W(20, 101) <= 0; play_W(20, 102) <= 0; play_W(20, 103) <= 0; play_W(20, 104) <= 0; play_W(20, 105) <= 0; play_W(20, 106) <= 0; play_W(20, 107) <= 0; play_W(20, 108) <= 0; play_W(20, 109) <= 0; play_W(20, 110) <= 0; play_W(20, 111) <= 0; play_W(20, 112) <= 0; play_W(20, 113) <= 0; play_W(20, 114) <= 0; play_W(20, 115) <= 0; play_W(20, 116) <= 0; play_W(20, 117) <= 1; play_W(20, 118) <= 1; play_W(20, 119) <= 1; play_W(20, 120) <= 1; play_W(20, 121) <= 1; play_W(20, 122) <= 1; play_W(20, 123) <= 0; play_W(20, 124) <= 0; play_W(20, 125) <= 0; play_W(20, 126) <= 0; play_W(20, 127) <= 0; play_W(20, 128) <= 0; play_W(20, 129) <= 0; play_W(20, 130) <= 0; play_W(20, 131) <= 0; play_W(20, 132) <= 0; play_W(20, 133) <= 0; play_W(20, 134) <= 0; play_W(20, 135) <= 0; play_W(20, 136) <= 0; play_W(20, 137) <= 0; play_W(20, 138) <= 0; play_W(20, 139) <= 0; play_W(20, 140) <= 0; play_W(20, 141) <= 0; play_W(20, 142) <= 0; play_W(20, 143) <= 0; play_W(20, 144) <= 0; play_W(20, 145) <= 0; play_W(20, 146) <= 0; play_W(20, 147) <= 0; play_W(20, 148) <= 0; play_W(20, 149) <= 0; play_W(20, 150) <= 0; play_W(20, 151) <= 0; play_W(20, 152) <= 0; play_W(20, 153) <= 0; play_W(20, 154) <= 0; play_W(20, 155) <= 0; play_W(20, 156) <= 0; play_W(20, 157) <= 0; play_W(20, 158) <= 0; play_W(20, 159) <= 0; play_W(20, 160) <= 0; play_W(20, 161) <= 0; play_W(20, 162) <= 0; play_W(20, 163) <= 0; play_W(20, 164) <= 0; play_W(20, 165) <= 1; play_W(20, 166) <= 1; play_W(20, 167) <= 1; play_W(20, 168) <= 1; play_W(20, 169) <= 1; play_W(20, 170) <= 1; play_W(20, 171) <= 0; play_W(20, 172) <= 0; play_W(20, 173) <= 0; play_W(20, 174) <= 0; play_W(20, 175) <= 0; play_W(20, 176) <= 0; play_W(20, 177) <= 1; play_W(20, 178) <= 1; play_W(20, 179) <= 1; play_W(20, 180) <= 1; play_W(20, 181) <= 1; play_W(20, 182) <= 1; play_W(20, 183) <= 0; play_W(20, 184) <= 0; play_W(20, 185) <= 0; play_W(20, 186) <= 0; play_W(20, 187) <= 0; play_W(20, 188) <= 0; play_W(20, 189) <= 0; play_W(20, 190) <= 0; play_W(20, 191) <= 0; play_W(20, 192) <= 0; play_W(20, 193) <= 0; play_W(20, 194) <= 0; play_W(20, 195) <= 0; play_W(20, 196) <= 0; play_W(20, 197) <= 0; play_W(20, 198) <= 1; play_W(20, 199) <= 1; play_W(20, 200) <= 1; play_W(20, 201) <= 1; play_W(20, 202) <= 1; play_W(20, 203) <= 1; play_W(20, 204) <= 0; play_W(20, 205) <= 0; play_W(20, 206) <= 0; play_W(20, 207) <= 0; play_W(20, 208) <= 0; play_W(20, 209) <= 0; play_W(20, 210) <= 0; play_W(20, 211) <= 0; play_W(20, 212) <= 0; play_W(20, 213) <= 0; play_W(20, 214) <= 0; play_W(20, 215) <= 0; play_W(20, 216) <= 1; play_W(20, 217) <= 1; play_W(20, 218) <= 1; play_W(20, 219) <= 1; play_W(20, 220) <= 1; play_W(20, 221) <= 1; play_W(20, 222) <= 0; play_W(20, 223) <= 0; play_W(20, 224) <= 0; play_W(20, 225) <= 0; play_W(20, 226) <= 0; play_W(20, 227) <= 0; play_W(20, 228) <= 0; play_W(20, 229) <= 0; play_W(20, 230) <= 0; play_W(20, 231) <= 1; play_W(20, 232) <= 1; play_W(20, 233) <= 1; play_W(20, 234) <= 1; play_W(20, 235) <= 1; play_W(20, 236) <= 1; play_W(20, 237) <= 0; play_W(20, 238) <= 0; play_W(20, 239) <= 0; play_W(20, 240) <= 0; play_W(20, 241) <= 0; play_W(20, 242) <= 0; play_W(20, 243) <= 0; play_W(20, 244) <= 0; play_W(20, 245) <= 0; play_W(20, 246) <= 1; play_W(20, 247) <= 1; play_W(20, 248) <= 1; play_W(20, 249) <= 1; play_W(20, 250) <= 1; play_W(20, 251) <= 1; play_W(20, 252) <= 0; play_W(20, 253) <= 0; play_W(20, 254) <= 0; play_W(20, 255) <= 0; play_W(20, 256) <= 0; play_W(20, 257) <= 0; play_W(20, 258) <= 1; play_W(20, 259) <= 1; play_W(20, 260) <= 1; play_W(20, 261) <= 1; play_W(20, 262) <= 1; play_W(20, 263) <= 1; play_W(20, 264) <= 0; play_W(20, 265) <= 0; play_W(20, 266) <= 0; play_W(20, 267) <= 0; play_W(20, 268) <= 0; play_W(20, 269) <= 0; 
play_W(21, 0) <= 0; play_W(21, 1) <= 0; play_W(21, 2) <= 0; play_W(21, 3) <= 1; play_W(21, 4) <= 1; play_W(21, 5) <= 1; play_W(21, 6) <= 1; play_W(21, 7) <= 1; play_W(21, 8) <= 1; play_W(21, 9) <= 0; play_W(21, 10) <= 0; play_W(21, 11) <= 0; play_W(21, 12) <= 0; play_W(21, 13) <= 0; play_W(21, 14) <= 0; play_W(21, 15) <= 0; play_W(21, 16) <= 0; play_W(21, 17) <= 0; play_W(21, 18) <= 0; play_W(21, 19) <= 0; play_W(21, 20) <= 0; play_W(21, 21) <= 0; play_W(21, 22) <= 0; play_W(21, 23) <= 0; play_W(21, 24) <= 0; play_W(21, 25) <= 0; play_W(21, 26) <= 0; play_W(21, 27) <= 0; play_W(21, 28) <= 0; play_W(21, 29) <= 0; play_W(21, 30) <= 1; play_W(21, 31) <= 1; play_W(21, 32) <= 1; play_W(21, 33) <= 1; play_W(21, 34) <= 1; play_W(21, 35) <= 1; play_W(21, 36) <= 0; play_W(21, 37) <= 0; play_W(21, 38) <= 0; play_W(21, 39) <= 0; play_W(21, 40) <= 0; play_W(21, 41) <= 0; play_W(21, 42) <= 0; play_W(21, 43) <= 0; play_W(21, 44) <= 0; play_W(21, 45) <= 1; play_W(21, 46) <= 1; play_W(21, 47) <= 1; play_W(21, 48) <= 0; play_W(21, 49) <= 0; play_W(21, 50) <= 0; play_W(21, 51) <= 0; play_W(21, 52) <= 0; play_W(21, 53) <= 0; play_W(21, 54) <= 1; play_W(21, 55) <= 1; play_W(21, 56) <= 1; play_W(21, 57) <= 1; play_W(21, 58) <= 1; play_W(21, 59) <= 1; play_W(21, 60) <= 0; play_W(21, 61) <= 0; play_W(21, 62) <= 0; play_W(21, 63) <= 0; play_W(21, 64) <= 0; play_W(21, 65) <= 0; play_W(21, 66) <= 0; play_W(21, 67) <= 0; play_W(21, 68) <= 0; play_W(21, 69) <= 1; play_W(21, 70) <= 1; play_W(21, 71) <= 1; play_W(21, 72) <= 1; play_W(21, 73) <= 1; play_W(21, 74) <= 1; play_W(21, 75) <= 0; play_W(21, 76) <= 0; play_W(21, 77) <= 0; play_W(21, 78) <= 0; play_W(21, 79) <= 0; play_W(21, 80) <= 0; play_W(21, 81) <= 0; play_W(21, 82) <= 0; play_W(21, 83) <= 0; play_W(21, 84) <= 0; play_W(21, 85) <= 0; play_W(21, 86) <= 0; play_W(21, 87) <= 0; play_W(21, 88) <= 0; play_W(21, 89) <= 0; play_W(21, 90) <= 1; play_W(21, 91) <= 1; play_W(21, 92) <= 1; play_W(21, 93) <= 1; play_W(21, 94) <= 1; play_W(21, 95) <= 1; play_W(21, 96) <= 0; play_W(21, 97) <= 0; play_W(21, 98) <= 0; play_W(21, 99) <= 0; play_W(21, 100) <= 0; play_W(21, 101) <= 0; play_W(21, 102) <= 0; play_W(21, 103) <= 0; play_W(21, 104) <= 0; play_W(21, 105) <= 0; play_W(21, 106) <= 0; play_W(21, 107) <= 0; play_W(21, 108) <= 0; play_W(21, 109) <= 0; play_W(21, 110) <= 0; play_W(21, 111) <= 0; play_W(21, 112) <= 0; play_W(21, 113) <= 0; play_W(21, 114) <= 0; play_W(21, 115) <= 0; play_W(21, 116) <= 0; play_W(21, 117) <= 1; play_W(21, 118) <= 1; play_W(21, 119) <= 1; play_W(21, 120) <= 1; play_W(21, 121) <= 1; play_W(21, 122) <= 1; play_W(21, 123) <= 0; play_W(21, 124) <= 0; play_W(21, 125) <= 0; play_W(21, 126) <= 0; play_W(21, 127) <= 0; play_W(21, 128) <= 0; play_W(21, 129) <= 0; play_W(21, 130) <= 0; play_W(21, 131) <= 0; play_W(21, 132) <= 0; play_W(21, 133) <= 0; play_W(21, 134) <= 0; play_W(21, 135) <= 0; play_W(21, 136) <= 0; play_W(21, 137) <= 0; play_W(21, 138) <= 0; play_W(21, 139) <= 0; play_W(21, 140) <= 0; play_W(21, 141) <= 0; play_W(21, 142) <= 0; play_W(21, 143) <= 0; play_W(21, 144) <= 0; play_W(21, 145) <= 0; play_W(21, 146) <= 0; play_W(21, 147) <= 0; play_W(21, 148) <= 0; play_W(21, 149) <= 0; play_W(21, 150) <= 0; play_W(21, 151) <= 0; play_W(21, 152) <= 0; play_W(21, 153) <= 0; play_W(21, 154) <= 0; play_W(21, 155) <= 0; play_W(21, 156) <= 0; play_W(21, 157) <= 0; play_W(21, 158) <= 0; play_W(21, 159) <= 0; play_W(21, 160) <= 0; play_W(21, 161) <= 0; play_W(21, 162) <= 0; play_W(21, 163) <= 0; play_W(21, 164) <= 0; play_W(21, 165) <= 1; play_W(21, 166) <= 1; play_W(21, 167) <= 1; play_W(21, 168) <= 1; play_W(21, 169) <= 1; play_W(21, 170) <= 1; play_W(21, 171) <= 0; play_W(21, 172) <= 0; play_W(21, 173) <= 0; play_W(21, 174) <= 0; play_W(21, 175) <= 0; play_W(21, 176) <= 0; play_W(21, 177) <= 1; play_W(21, 178) <= 1; play_W(21, 179) <= 1; play_W(21, 180) <= 1; play_W(21, 181) <= 1; play_W(21, 182) <= 1; play_W(21, 183) <= 0; play_W(21, 184) <= 0; play_W(21, 185) <= 0; play_W(21, 186) <= 0; play_W(21, 187) <= 0; play_W(21, 188) <= 0; play_W(21, 189) <= 0; play_W(21, 190) <= 0; play_W(21, 191) <= 0; play_W(21, 192) <= 0; play_W(21, 193) <= 0; play_W(21, 194) <= 0; play_W(21, 195) <= 0; play_W(21, 196) <= 0; play_W(21, 197) <= 0; play_W(21, 198) <= 1; play_W(21, 199) <= 1; play_W(21, 200) <= 1; play_W(21, 201) <= 1; play_W(21, 202) <= 1; play_W(21, 203) <= 1; play_W(21, 204) <= 0; play_W(21, 205) <= 0; play_W(21, 206) <= 0; play_W(21, 207) <= 0; play_W(21, 208) <= 0; play_W(21, 209) <= 0; play_W(21, 210) <= 0; play_W(21, 211) <= 0; play_W(21, 212) <= 0; play_W(21, 213) <= 0; play_W(21, 214) <= 0; play_W(21, 215) <= 0; play_W(21, 216) <= 1; play_W(21, 217) <= 1; play_W(21, 218) <= 1; play_W(21, 219) <= 1; play_W(21, 220) <= 1; play_W(21, 221) <= 1; play_W(21, 222) <= 0; play_W(21, 223) <= 0; play_W(21, 224) <= 0; play_W(21, 225) <= 0; play_W(21, 226) <= 0; play_W(21, 227) <= 0; play_W(21, 228) <= 0; play_W(21, 229) <= 0; play_W(21, 230) <= 0; play_W(21, 231) <= 1; play_W(21, 232) <= 1; play_W(21, 233) <= 1; play_W(21, 234) <= 1; play_W(21, 235) <= 1; play_W(21, 236) <= 1; play_W(21, 237) <= 0; play_W(21, 238) <= 0; play_W(21, 239) <= 0; play_W(21, 240) <= 0; play_W(21, 241) <= 0; play_W(21, 242) <= 0; play_W(21, 243) <= 0; play_W(21, 244) <= 0; play_W(21, 245) <= 0; play_W(21, 246) <= 1; play_W(21, 247) <= 1; play_W(21, 248) <= 1; play_W(21, 249) <= 1; play_W(21, 250) <= 1; play_W(21, 251) <= 1; play_W(21, 252) <= 0; play_W(21, 253) <= 0; play_W(21, 254) <= 0; play_W(21, 255) <= 0; play_W(21, 256) <= 0; play_W(21, 257) <= 0; play_W(21, 258) <= 1; play_W(21, 259) <= 1; play_W(21, 260) <= 1; play_W(21, 261) <= 1; play_W(21, 262) <= 1; play_W(21, 263) <= 1; play_W(21, 264) <= 0; play_W(21, 265) <= 0; play_W(21, 266) <= 0; play_W(21, 267) <= 0; play_W(21, 268) <= 0; play_W(21, 269) <= 0; 
play_W(22, 0) <= 0; play_W(22, 1) <= 0; play_W(22, 2) <= 0; play_W(22, 3) <= 1; play_W(22, 4) <= 1; play_W(22, 5) <= 1; play_W(22, 6) <= 1; play_W(22, 7) <= 1; play_W(22, 8) <= 1; play_W(22, 9) <= 0; play_W(22, 10) <= 0; play_W(22, 11) <= 0; play_W(22, 12) <= 0; play_W(22, 13) <= 0; play_W(22, 14) <= 0; play_W(22, 15) <= 0; play_W(22, 16) <= 0; play_W(22, 17) <= 0; play_W(22, 18) <= 0; play_W(22, 19) <= 0; play_W(22, 20) <= 0; play_W(22, 21) <= 0; play_W(22, 22) <= 0; play_W(22, 23) <= 0; play_W(22, 24) <= 0; play_W(22, 25) <= 0; play_W(22, 26) <= 0; play_W(22, 27) <= 0; play_W(22, 28) <= 0; play_W(22, 29) <= 0; play_W(22, 30) <= 1; play_W(22, 31) <= 1; play_W(22, 32) <= 1; play_W(22, 33) <= 1; play_W(22, 34) <= 1; play_W(22, 35) <= 1; play_W(22, 36) <= 0; play_W(22, 37) <= 0; play_W(22, 38) <= 0; play_W(22, 39) <= 0; play_W(22, 40) <= 0; play_W(22, 41) <= 0; play_W(22, 42) <= 0; play_W(22, 43) <= 0; play_W(22, 44) <= 0; play_W(22, 45) <= 1; play_W(22, 46) <= 1; play_W(22, 47) <= 1; play_W(22, 48) <= 0; play_W(22, 49) <= 0; play_W(22, 50) <= 0; play_W(22, 51) <= 0; play_W(22, 52) <= 0; play_W(22, 53) <= 0; play_W(22, 54) <= 1; play_W(22, 55) <= 1; play_W(22, 56) <= 1; play_W(22, 57) <= 1; play_W(22, 58) <= 1; play_W(22, 59) <= 1; play_W(22, 60) <= 0; play_W(22, 61) <= 0; play_W(22, 62) <= 0; play_W(22, 63) <= 0; play_W(22, 64) <= 0; play_W(22, 65) <= 0; play_W(22, 66) <= 0; play_W(22, 67) <= 0; play_W(22, 68) <= 0; play_W(22, 69) <= 1; play_W(22, 70) <= 1; play_W(22, 71) <= 1; play_W(22, 72) <= 1; play_W(22, 73) <= 1; play_W(22, 74) <= 1; play_W(22, 75) <= 0; play_W(22, 76) <= 0; play_W(22, 77) <= 0; play_W(22, 78) <= 0; play_W(22, 79) <= 0; play_W(22, 80) <= 0; play_W(22, 81) <= 0; play_W(22, 82) <= 0; play_W(22, 83) <= 0; play_W(22, 84) <= 0; play_W(22, 85) <= 0; play_W(22, 86) <= 0; play_W(22, 87) <= 0; play_W(22, 88) <= 0; play_W(22, 89) <= 0; play_W(22, 90) <= 1; play_W(22, 91) <= 1; play_W(22, 92) <= 1; play_W(22, 93) <= 1; play_W(22, 94) <= 1; play_W(22, 95) <= 1; play_W(22, 96) <= 0; play_W(22, 97) <= 0; play_W(22, 98) <= 0; play_W(22, 99) <= 0; play_W(22, 100) <= 0; play_W(22, 101) <= 0; play_W(22, 102) <= 0; play_W(22, 103) <= 0; play_W(22, 104) <= 0; play_W(22, 105) <= 0; play_W(22, 106) <= 0; play_W(22, 107) <= 0; play_W(22, 108) <= 0; play_W(22, 109) <= 0; play_W(22, 110) <= 0; play_W(22, 111) <= 0; play_W(22, 112) <= 0; play_W(22, 113) <= 0; play_W(22, 114) <= 0; play_W(22, 115) <= 0; play_W(22, 116) <= 0; play_W(22, 117) <= 1; play_W(22, 118) <= 1; play_W(22, 119) <= 1; play_W(22, 120) <= 1; play_W(22, 121) <= 1; play_W(22, 122) <= 1; play_W(22, 123) <= 0; play_W(22, 124) <= 0; play_W(22, 125) <= 0; play_W(22, 126) <= 0; play_W(22, 127) <= 0; play_W(22, 128) <= 0; play_W(22, 129) <= 0; play_W(22, 130) <= 0; play_W(22, 131) <= 0; play_W(22, 132) <= 0; play_W(22, 133) <= 0; play_W(22, 134) <= 0; play_W(22, 135) <= 0; play_W(22, 136) <= 0; play_W(22, 137) <= 0; play_W(22, 138) <= 0; play_W(22, 139) <= 0; play_W(22, 140) <= 0; play_W(22, 141) <= 0; play_W(22, 142) <= 0; play_W(22, 143) <= 0; play_W(22, 144) <= 0; play_W(22, 145) <= 0; play_W(22, 146) <= 0; play_W(22, 147) <= 0; play_W(22, 148) <= 0; play_W(22, 149) <= 0; play_W(22, 150) <= 0; play_W(22, 151) <= 0; play_W(22, 152) <= 0; play_W(22, 153) <= 0; play_W(22, 154) <= 0; play_W(22, 155) <= 0; play_W(22, 156) <= 0; play_W(22, 157) <= 0; play_W(22, 158) <= 0; play_W(22, 159) <= 0; play_W(22, 160) <= 0; play_W(22, 161) <= 0; play_W(22, 162) <= 0; play_W(22, 163) <= 0; play_W(22, 164) <= 0; play_W(22, 165) <= 1; play_W(22, 166) <= 1; play_W(22, 167) <= 1; play_W(22, 168) <= 1; play_W(22, 169) <= 1; play_W(22, 170) <= 1; play_W(22, 171) <= 0; play_W(22, 172) <= 0; play_W(22, 173) <= 0; play_W(22, 174) <= 0; play_W(22, 175) <= 0; play_W(22, 176) <= 0; play_W(22, 177) <= 1; play_W(22, 178) <= 1; play_W(22, 179) <= 1; play_W(22, 180) <= 1; play_W(22, 181) <= 1; play_W(22, 182) <= 1; play_W(22, 183) <= 0; play_W(22, 184) <= 0; play_W(22, 185) <= 0; play_W(22, 186) <= 0; play_W(22, 187) <= 0; play_W(22, 188) <= 0; play_W(22, 189) <= 0; play_W(22, 190) <= 0; play_W(22, 191) <= 0; play_W(22, 192) <= 0; play_W(22, 193) <= 0; play_W(22, 194) <= 0; play_W(22, 195) <= 0; play_W(22, 196) <= 0; play_W(22, 197) <= 0; play_W(22, 198) <= 1; play_W(22, 199) <= 1; play_W(22, 200) <= 1; play_W(22, 201) <= 1; play_W(22, 202) <= 1; play_W(22, 203) <= 1; play_W(22, 204) <= 0; play_W(22, 205) <= 0; play_W(22, 206) <= 0; play_W(22, 207) <= 0; play_W(22, 208) <= 0; play_W(22, 209) <= 0; play_W(22, 210) <= 0; play_W(22, 211) <= 0; play_W(22, 212) <= 0; play_W(22, 213) <= 0; play_W(22, 214) <= 0; play_W(22, 215) <= 0; play_W(22, 216) <= 1; play_W(22, 217) <= 1; play_W(22, 218) <= 1; play_W(22, 219) <= 1; play_W(22, 220) <= 1; play_W(22, 221) <= 1; play_W(22, 222) <= 0; play_W(22, 223) <= 0; play_W(22, 224) <= 0; play_W(22, 225) <= 0; play_W(22, 226) <= 0; play_W(22, 227) <= 0; play_W(22, 228) <= 0; play_W(22, 229) <= 0; play_W(22, 230) <= 0; play_W(22, 231) <= 1; play_W(22, 232) <= 1; play_W(22, 233) <= 1; play_W(22, 234) <= 1; play_W(22, 235) <= 1; play_W(22, 236) <= 1; play_W(22, 237) <= 0; play_W(22, 238) <= 0; play_W(22, 239) <= 0; play_W(22, 240) <= 0; play_W(22, 241) <= 0; play_W(22, 242) <= 0; play_W(22, 243) <= 0; play_W(22, 244) <= 0; play_W(22, 245) <= 0; play_W(22, 246) <= 1; play_W(22, 247) <= 1; play_W(22, 248) <= 1; play_W(22, 249) <= 1; play_W(22, 250) <= 1; play_W(22, 251) <= 1; play_W(22, 252) <= 0; play_W(22, 253) <= 0; play_W(22, 254) <= 0; play_W(22, 255) <= 0; play_W(22, 256) <= 0; play_W(22, 257) <= 0; play_W(22, 258) <= 1; play_W(22, 259) <= 1; play_W(22, 260) <= 1; play_W(22, 261) <= 1; play_W(22, 262) <= 1; play_W(22, 263) <= 1; play_W(22, 264) <= 0; play_W(22, 265) <= 0; play_W(22, 266) <= 0; play_W(22, 267) <= 0; play_W(22, 268) <= 0; play_W(22, 269) <= 0; 
play_W(23, 0) <= 0; play_W(23, 1) <= 0; play_W(23, 2) <= 0; play_W(23, 3) <= 1; play_W(23, 4) <= 1; play_W(23, 5) <= 1; play_W(23, 6) <= 1; play_W(23, 7) <= 1; play_W(23, 8) <= 1; play_W(23, 9) <= 0; play_W(23, 10) <= 0; play_W(23, 11) <= 0; play_W(23, 12) <= 0; play_W(23, 13) <= 0; play_W(23, 14) <= 0; play_W(23, 15) <= 0; play_W(23, 16) <= 0; play_W(23, 17) <= 0; play_W(23, 18) <= 0; play_W(23, 19) <= 0; play_W(23, 20) <= 0; play_W(23, 21) <= 0; play_W(23, 22) <= 0; play_W(23, 23) <= 0; play_W(23, 24) <= 0; play_W(23, 25) <= 0; play_W(23, 26) <= 0; play_W(23, 27) <= 0; play_W(23, 28) <= 0; play_W(23, 29) <= 0; play_W(23, 30) <= 1; play_W(23, 31) <= 1; play_W(23, 32) <= 1; play_W(23, 33) <= 1; play_W(23, 34) <= 1; play_W(23, 35) <= 1; play_W(23, 36) <= 0; play_W(23, 37) <= 0; play_W(23, 38) <= 0; play_W(23, 39) <= 0; play_W(23, 40) <= 0; play_W(23, 41) <= 0; play_W(23, 42) <= 0; play_W(23, 43) <= 0; play_W(23, 44) <= 0; play_W(23, 45) <= 1; play_W(23, 46) <= 1; play_W(23, 47) <= 1; play_W(23, 48) <= 0; play_W(23, 49) <= 0; play_W(23, 50) <= 0; play_W(23, 51) <= 0; play_W(23, 52) <= 0; play_W(23, 53) <= 0; play_W(23, 54) <= 1; play_W(23, 55) <= 1; play_W(23, 56) <= 1; play_W(23, 57) <= 1; play_W(23, 58) <= 1; play_W(23, 59) <= 1; play_W(23, 60) <= 0; play_W(23, 61) <= 0; play_W(23, 62) <= 0; play_W(23, 63) <= 0; play_W(23, 64) <= 0; play_W(23, 65) <= 0; play_W(23, 66) <= 0; play_W(23, 67) <= 0; play_W(23, 68) <= 0; play_W(23, 69) <= 1; play_W(23, 70) <= 1; play_W(23, 71) <= 1; play_W(23, 72) <= 1; play_W(23, 73) <= 1; play_W(23, 74) <= 1; play_W(23, 75) <= 0; play_W(23, 76) <= 0; play_W(23, 77) <= 0; play_W(23, 78) <= 0; play_W(23, 79) <= 0; play_W(23, 80) <= 0; play_W(23, 81) <= 0; play_W(23, 82) <= 0; play_W(23, 83) <= 0; play_W(23, 84) <= 0; play_W(23, 85) <= 0; play_W(23, 86) <= 0; play_W(23, 87) <= 0; play_W(23, 88) <= 0; play_W(23, 89) <= 0; play_W(23, 90) <= 1; play_W(23, 91) <= 1; play_W(23, 92) <= 1; play_W(23, 93) <= 1; play_W(23, 94) <= 1; play_W(23, 95) <= 1; play_W(23, 96) <= 0; play_W(23, 97) <= 0; play_W(23, 98) <= 0; play_W(23, 99) <= 0; play_W(23, 100) <= 0; play_W(23, 101) <= 0; play_W(23, 102) <= 0; play_W(23, 103) <= 0; play_W(23, 104) <= 0; play_W(23, 105) <= 0; play_W(23, 106) <= 0; play_W(23, 107) <= 0; play_W(23, 108) <= 0; play_W(23, 109) <= 0; play_W(23, 110) <= 0; play_W(23, 111) <= 0; play_W(23, 112) <= 0; play_W(23, 113) <= 0; play_W(23, 114) <= 0; play_W(23, 115) <= 0; play_W(23, 116) <= 0; play_W(23, 117) <= 1; play_W(23, 118) <= 1; play_W(23, 119) <= 1; play_W(23, 120) <= 1; play_W(23, 121) <= 1; play_W(23, 122) <= 1; play_W(23, 123) <= 0; play_W(23, 124) <= 0; play_W(23, 125) <= 0; play_W(23, 126) <= 0; play_W(23, 127) <= 0; play_W(23, 128) <= 0; play_W(23, 129) <= 0; play_W(23, 130) <= 0; play_W(23, 131) <= 0; play_W(23, 132) <= 0; play_W(23, 133) <= 0; play_W(23, 134) <= 0; play_W(23, 135) <= 0; play_W(23, 136) <= 0; play_W(23, 137) <= 0; play_W(23, 138) <= 0; play_W(23, 139) <= 0; play_W(23, 140) <= 0; play_W(23, 141) <= 0; play_W(23, 142) <= 0; play_W(23, 143) <= 0; play_W(23, 144) <= 0; play_W(23, 145) <= 0; play_W(23, 146) <= 0; play_W(23, 147) <= 0; play_W(23, 148) <= 0; play_W(23, 149) <= 0; play_W(23, 150) <= 0; play_W(23, 151) <= 0; play_W(23, 152) <= 0; play_W(23, 153) <= 0; play_W(23, 154) <= 0; play_W(23, 155) <= 0; play_W(23, 156) <= 0; play_W(23, 157) <= 0; play_W(23, 158) <= 0; play_W(23, 159) <= 0; play_W(23, 160) <= 0; play_W(23, 161) <= 0; play_W(23, 162) <= 0; play_W(23, 163) <= 0; play_W(23, 164) <= 0; play_W(23, 165) <= 1; play_W(23, 166) <= 1; play_W(23, 167) <= 1; play_W(23, 168) <= 1; play_W(23, 169) <= 1; play_W(23, 170) <= 1; play_W(23, 171) <= 0; play_W(23, 172) <= 0; play_W(23, 173) <= 0; play_W(23, 174) <= 0; play_W(23, 175) <= 0; play_W(23, 176) <= 0; play_W(23, 177) <= 1; play_W(23, 178) <= 1; play_W(23, 179) <= 1; play_W(23, 180) <= 1; play_W(23, 181) <= 1; play_W(23, 182) <= 1; play_W(23, 183) <= 0; play_W(23, 184) <= 0; play_W(23, 185) <= 0; play_W(23, 186) <= 0; play_W(23, 187) <= 0; play_W(23, 188) <= 0; play_W(23, 189) <= 0; play_W(23, 190) <= 0; play_W(23, 191) <= 0; play_W(23, 192) <= 0; play_W(23, 193) <= 0; play_W(23, 194) <= 0; play_W(23, 195) <= 0; play_W(23, 196) <= 0; play_W(23, 197) <= 0; play_W(23, 198) <= 1; play_W(23, 199) <= 1; play_W(23, 200) <= 1; play_W(23, 201) <= 1; play_W(23, 202) <= 1; play_W(23, 203) <= 1; play_W(23, 204) <= 0; play_W(23, 205) <= 0; play_W(23, 206) <= 0; play_W(23, 207) <= 0; play_W(23, 208) <= 0; play_W(23, 209) <= 0; play_W(23, 210) <= 0; play_W(23, 211) <= 0; play_W(23, 212) <= 0; play_W(23, 213) <= 0; play_W(23, 214) <= 0; play_W(23, 215) <= 0; play_W(23, 216) <= 1; play_W(23, 217) <= 1; play_W(23, 218) <= 1; play_W(23, 219) <= 1; play_W(23, 220) <= 1; play_W(23, 221) <= 1; play_W(23, 222) <= 0; play_W(23, 223) <= 0; play_W(23, 224) <= 0; play_W(23, 225) <= 0; play_W(23, 226) <= 0; play_W(23, 227) <= 0; play_W(23, 228) <= 0; play_W(23, 229) <= 0; play_W(23, 230) <= 0; play_W(23, 231) <= 1; play_W(23, 232) <= 1; play_W(23, 233) <= 1; play_W(23, 234) <= 1; play_W(23, 235) <= 1; play_W(23, 236) <= 1; play_W(23, 237) <= 0; play_W(23, 238) <= 0; play_W(23, 239) <= 0; play_W(23, 240) <= 0; play_W(23, 241) <= 0; play_W(23, 242) <= 0; play_W(23, 243) <= 0; play_W(23, 244) <= 0; play_W(23, 245) <= 0; play_W(23, 246) <= 1; play_W(23, 247) <= 1; play_W(23, 248) <= 1; play_W(23, 249) <= 1; play_W(23, 250) <= 1; play_W(23, 251) <= 1; play_W(23, 252) <= 0; play_W(23, 253) <= 0; play_W(23, 254) <= 0; play_W(23, 255) <= 0; play_W(23, 256) <= 0; play_W(23, 257) <= 0; play_W(23, 258) <= 1; play_W(23, 259) <= 1; play_W(23, 260) <= 1; play_W(23, 261) <= 1; play_W(23, 262) <= 1; play_W(23, 263) <= 1; play_W(23, 264) <= 0; play_W(23, 265) <= 0; play_W(23, 266) <= 0; play_W(23, 267) <= 0; play_W(23, 268) <= 0; play_W(23, 269) <= 0; 
play_W(24, 0) <= 0; play_W(24, 1) <= 0; play_W(24, 2) <= 0; play_W(24, 3) <= 1; play_W(24, 4) <= 1; play_W(24, 5) <= 1; play_W(24, 6) <= 1; play_W(24, 7) <= 1; play_W(24, 8) <= 1; play_W(24, 9) <= 0; play_W(24, 10) <= 0; play_W(24, 11) <= 0; play_W(24, 12) <= 0; play_W(24, 13) <= 0; play_W(24, 14) <= 0; play_W(24, 15) <= 0; play_W(24, 16) <= 0; play_W(24, 17) <= 0; play_W(24, 18) <= 0; play_W(24, 19) <= 0; play_W(24, 20) <= 0; play_W(24, 21) <= 0; play_W(24, 22) <= 0; play_W(24, 23) <= 0; play_W(24, 24) <= 0; play_W(24, 25) <= 0; play_W(24, 26) <= 0; play_W(24, 27) <= 0; play_W(24, 28) <= 0; play_W(24, 29) <= 0; play_W(24, 30) <= 1; play_W(24, 31) <= 1; play_W(24, 32) <= 1; play_W(24, 33) <= 1; play_W(24, 34) <= 1; play_W(24, 35) <= 1; play_W(24, 36) <= 0; play_W(24, 37) <= 0; play_W(24, 38) <= 0; play_W(24, 39) <= 0; play_W(24, 40) <= 0; play_W(24, 41) <= 0; play_W(24, 42) <= 1; play_W(24, 43) <= 1; play_W(24, 44) <= 1; play_W(24, 45) <= 1; play_W(24, 46) <= 1; play_W(24, 47) <= 1; play_W(24, 48) <= 0; play_W(24, 49) <= 0; play_W(24, 50) <= 0; play_W(24, 51) <= 0; play_W(24, 52) <= 0; play_W(24, 53) <= 0; play_W(24, 54) <= 1; play_W(24, 55) <= 1; play_W(24, 56) <= 1; play_W(24, 57) <= 1; play_W(24, 58) <= 1; play_W(24, 59) <= 1; play_W(24, 60) <= 0; play_W(24, 61) <= 0; play_W(24, 62) <= 0; play_W(24, 63) <= 0; play_W(24, 64) <= 0; play_W(24, 65) <= 0; play_W(24, 66) <= 0; play_W(24, 67) <= 0; play_W(24, 68) <= 0; play_W(24, 69) <= 1; play_W(24, 70) <= 1; play_W(24, 71) <= 1; play_W(24, 72) <= 1; play_W(24, 73) <= 1; play_W(24, 74) <= 1; play_W(24, 75) <= 0; play_W(24, 76) <= 0; play_W(24, 77) <= 0; play_W(24, 78) <= 0; play_W(24, 79) <= 0; play_W(24, 80) <= 0; play_W(24, 81) <= 0; play_W(24, 82) <= 0; play_W(24, 83) <= 0; play_W(24, 84) <= 0; play_W(24, 85) <= 0; play_W(24, 86) <= 0; play_W(24, 87) <= 0; play_W(24, 88) <= 0; play_W(24, 89) <= 0; play_W(24, 90) <= 1; play_W(24, 91) <= 1; play_W(24, 92) <= 1; play_W(24, 93) <= 1; play_W(24, 94) <= 1; play_W(24, 95) <= 1; play_W(24, 96) <= 0; play_W(24, 97) <= 0; play_W(24, 98) <= 0; play_W(24, 99) <= 0; play_W(24, 100) <= 0; play_W(24, 101) <= 0; play_W(24, 102) <= 0; play_W(24, 103) <= 0; play_W(24, 104) <= 0; play_W(24, 105) <= 0; play_W(24, 106) <= 0; play_W(24, 107) <= 0; play_W(24, 108) <= 0; play_W(24, 109) <= 0; play_W(24, 110) <= 0; play_W(24, 111) <= 0; play_W(24, 112) <= 0; play_W(24, 113) <= 0; play_W(24, 114) <= 0; play_W(24, 115) <= 0; play_W(24, 116) <= 0; play_W(24, 117) <= 0; play_W(24, 118) <= 0; play_W(24, 119) <= 0; play_W(24, 120) <= 0; play_W(24, 121) <= 0; play_W(24, 122) <= 0; play_W(24, 123) <= 0; play_W(24, 124) <= 0; play_W(24, 125) <= 0; play_W(24, 126) <= 0; play_W(24, 127) <= 0; play_W(24, 128) <= 0; play_W(24, 129) <= 0; play_W(24, 130) <= 0; play_W(24, 131) <= 0; play_W(24, 132) <= 0; play_W(24, 133) <= 0; play_W(24, 134) <= 0; play_W(24, 135) <= 0; play_W(24, 136) <= 0; play_W(24, 137) <= 0; play_W(24, 138) <= 0; play_W(24, 139) <= 0; play_W(24, 140) <= 0; play_W(24, 141) <= 0; play_W(24, 142) <= 0; play_W(24, 143) <= 0; play_W(24, 144) <= 0; play_W(24, 145) <= 0; play_W(24, 146) <= 0; play_W(24, 147) <= 0; play_W(24, 148) <= 0; play_W(24, 149) <= 0; play_W(24, 150) <= 0; play_W(24, 151) <= 0; play_W(24, 152) <= 0; play_W(24, 153) <= 0; play_W(24, 154) <= 0; play_W(24, 155) <= 0; play_W(24, 156) <= 0; play_W(24, 157) <= 0; play_W(24, 158) <= 0; play_W(24, 159) <= 0; play_W(24, 160) <= 0; play_W(24, 161) <= 0; play_W(24, 162) <= 0; play_W(24, 163) <= 0; play_W(24, 164) <= 0; play_W(24, 165) <= 1; play_W(24, 166) <= 1; play_W(24, 167) <= 1; play_W(24, 168) <= 1; play_W(24, 169) <= 1; play_W(24, 170) <= 1; play_W(24, 171) <= 0; play_W(24, 172) <= 0; play_W(24, 173) <= 0; play_W(24, 174) <= 0; play_W(24, 175) <= 0; play_W(24, 176) <= 0; play_W(24, 177) <= 1; play_W(24, 178) <= 1; play_W(24, 179) <= 1; play_W(24, 180) <= 1; play_W(24, 181) <= 1; play_W(24, 182) <= 1; play_W(24, 183) <= 0; play_W(24, 184) <= 0; play_W(24, 185) <= 0; play_W(24, 186) <= 0; play_W(24, 187) <= 0; play_W(24, 188) <= 0; play_W(24, 189) <= 0; play_W(24, 190) <= 0; play_W(24, 191) <= 0; play_W(24, 192) <= 0; play_W(24, 193) <= 0; play_W(24, 194) <= 0; play_W(24, 195) <= 0; play_W(24, 196) <= 0; play_W(24, 197) <= 0; play_W(24, 198) <= 1; play_W(24, 199) <= 1; play_W(24, 200) <= 1; play_W(24, 201) <= 1; play_W(24, 202) <= 1; play_W(24, 203) <= 1; play_W(24, 204) <= 0; play_W(24, 205) <= 0; play_W(24, 206) <= 0; play_W(24, 207) <= 0; play_W(24, 208) <= 0; play_W(24, 209) <= 0; play_W(24, 210) <= 0; play_W(24, 211) <= 0; play_W(24, 212) <= 0; play_W(24, 213) <= 0; play_W(24, 214) <= 0; play_W(24, 215) <= 0; play_W(24, 216) <= 1; play_W(24, 217) <= 1; play_W(24, 218) <= 1; play_W(24, 219) <= 1; play_W(24, 220) <= 1; play_W(24, 221) <= 1; play_W(24, 222) <= 0; play_W(24, 223) <= 0; play_W(24, 224) <= 0; play_W(24, 225) <= 0; play_W(24, 226) <= 0; play_W(24, 227) <= 0; play_W(24, 228) <= 0; play_W(24, 229) <= 0; play_W(24, 230) <= 0; play_W(24, 231) <= 1; play_W(24, 232) <= 1; play_W(24, 233) <= 1; play_W(24, 234) <= 1; play_W(24, 235) <= 1; play_W(24, 236) <= 1; play_W(24, 237) <= 0; play_W(24, 238) <= 0; play_W(24, 239) <= 0; play_W(24, 240) <= 0; play_W(24, 241) <= 0; play_W(24, 242) <= 0; play_W(24, 243) <= 0; play_W(24, 244) <= 0; play_W(24, 245) <= 0; play_W(24, 246) <= 1; play_W(24, 247) <= 1; play_W(24, 248) <= 1; play_W(24, 249) <= 1; play_W(24, 250) <= 1; play_W(24, 251) <= 1; play_W(24, 252) <= 0; play_W(24, 253) <= 0; play_W(24, 254) <= 0; play_W(24, 255) <= 0; play_W(24, 256) <= 0; play_W(24, 257) <= 0; play_W(24, 258) <= 1; play_W(24, 259) <= 1; play_W(24, 260) <= 1; play_W(24, 261) <= 1; play_W(24, 262) <= 1; play_W(24, 263) <= 1; play_W(24, 264) <= 0; play_W(24, 265) <= 0; play_W(24, 266) <= 0; play_W(24, 267) <= 0; play_W(24, 268) <= 0; play_W(24, 269) <= 0; 
play_W(25, 0) <= 0; play_W(25, 1) <= 0; play_W(25, 2) <= 0; play_W(25, 3) <= 1; play_W(25, 4) <= 1; play_W(25, 5) <= 1; play_W(25, 6) <= 1; play_W(25, 7) <= 1; play_W(25, 8) <= 1; play_W(25, 9) <= 0; play_W(25, 10) <= 0; play_W(25, 11) <= 0; play_W(25, 12) <= 0; play_W(25, 13) <= 0; play_W(25, 14) <= 0; play_W(25, 15) <= 0; play_W(25, 16) <= 0; play_W(25, 17) <= 0; play_W(25, 18) <= 0; play_W(25, 19) <= 0; play_W(25, 20) <= 0; play_W(25, 21) <= 0; play_W(25, 22) <= 0; play_W(25, 23) <= 0; play_W(25, 24) <= 0; play_W(25, 25) <= 0; play_W(25, 26) <= 0; play_W(25, 27) <= 0; play_W(25, 28) <= 0; play_W(25, 29) <= 0; play_W(25, 30) <= 1; play_W(25, 31) <= 1; play_W(25, 32) <= 1; play_W(25, 33) <= 1; play_W(25, 34) <= 1; play_W(25, 35) <= 1; play_W(25, 36) <= 0; play_W(25, 37) <= 0; play_W(25, 38) <= 0; play_W(25, 39) <= 0; play_W(25, 40) <= 0; play_W(25, 41) <= 0; play_W(25, 42) <= 1; play_W(25, 43) <= 1; play_W(25, 44) <= 1; play_W(25, 45) <= 1; play_W(25, 46) <= 1; play_W(25, 47) <= 1; play_W(25, 48) <= 0; play_W(25, 49) <= 0; play_W(25, 50) <= 0; play_W(25, 51) <= 0; play_W(25, 52) <= 0; play_W(25, 53) <= 0; play_W(25, 54) <= 1; play_W(25, 55) <= 1; play_W(25, 56) <= 1; play_W(25, 57) <= 1; play_W(25, 58) <= 1; play_W(25, 59) <= 1; play_W(25, 60) <= 0; play_W(25, 61) <= 0; play_W(25, 62) <= 0; play_W(25, 63) <= 0; play_W(25, 64) <= 0; play_W(25, 65) <= 0; play_W(25, 66) <= 0; play_W(25, 67) <= 0; play_W(25, 68) <= 0; play_W(25, 69) <= 1; play_W(25, 70) <= 1; play_W(25, 71) <= 1; play_W(25, 72) <= 1; play_W(25, 73) <= 1; play_W(25, 74) <= 1; play_W(25, 75) <= 0; play_W(25, 76) <= 0; play_W(25, 77) <= 0; play_W(25, 78) <= 0; play_W(25, 79) <= 0; play_W(25, 80) <= 0; play_W(25, 81) <= 0; play_W(25, 82) <= 0; play_W(25, 83) <= 0; play_W(25, 84) <= 0; play_W(25, 85) <= 0; play_W(25, 86) <= 0; play_W(25, 87) <= 0; play_W(25, 88) <= 0; play_W(25, 89) <= 0; play_W(25, 90) <= 1; play_W(25, 91) <= 1; play_W(25, 92) <= 1; play_W(25, 93) <= 1; play_W(25, 94) <= 1; play_W(25, 95) <= 1; play_W(25, 96) <= 0; play_W(25, 97) <= 0; play_W(25, 98) <= 0; play_W(25, 99) <= 0; play_W(25, 100) <= 0; play_W(25, 101) <= 0; play_W(25, 102) <= 0; play_W(25, 103) <= 0; play_W(25, 104) <= 0; play_W(25, 105) <= 0; play_W(25, 106) <= 0; play_W(25, 107) <= 0; play_W(25, 108) <= 0; play_W(25, 109) <= 0; play_W(25, 110) <= 0; play_W(25, 111) <= 0; play_W(25, 112) <= 0; play_W(25, 113) <= 0; play_W(25, 114) <= 0; play_W(25, 115) <= 0; play_W(25, 116) <= 0; play_W(25, 117) <= 0; play_W(25, 118) <= 0; play_W(25, 119) <= 0; play_W(25, 120) <= 0; play_W(25, 121) <= 0; play_W(25, 122) <= 0; play_W(25, 123) <= 0; play_W(25, 124) <= 0; play_W(25, 125) <= 0; play_W(25, 126) <= 0; play_W(25, 127) <= 0; play_W(25, 128) <= 0; play_W(25, 129) <= 0; play_W(25, 130) <= 0; play_W(25, 131) <= 0; play_W(25, 132) <= 0; play_W(25, 133) <= 0; play_W(25, 134) <= 0; play_W(25, 135) <= 0; play_W(25, 136) <= 0; play_W(25, 137) <= 0; play_W(25, 138) <= 0; play_W(25, 139) <= 0; play_W(25, 140) <= 0; play_W(25, 141) <= 0; play_W(25, 142) <= 0; play_W(25, 143) <= 0; play_W(25, 144) <= 0; play_W(25, 145) <= 0; play_W(25, 146) <= 0; play_W(25, 147) <= 0; play_W(25, 148) <= 0; play_W(25, 149) <= 0; play_W(25, 150) <= 0; play_W(25, 151) <= 0; play_W(25, 152) <= 0; play_W(25, 153) <= 0; play_W(25, 154) <= 0; play_W(25, 155) <= 0; play_W(25, 156) <= 0; play_W(25, 157) <= 0; play_W(25, 158) <= 0; play_W(25, 159) <= 0; play_W(25, 160) <= 0; play_W(25, 161) <= 0; play_W(25, 162) <= 0; play_W(25, 163) <= 0; play_W(25, 164) <= 0; play_W(25, 165) <= 1; play_W(25, 166) <= 1; play_W(25, 167) <= 1; play_W(25, 168) <= 1; play_W(25, 169) <= 1; play_W(25, 170) <= 1; play_W(25, 171) <= 0; play_W(25, 172) <= 0; play_W(25, 173) <= 0; play_W(25, 174) <= 0; play_W(25, 175) <= 0; play_W(25, 176) <= 0; play_W(25, 177) <= 1; play_W(25, 178) <= 1; play_W(25, 179) <= 1; play_W(25, 180) <= 1; play_W(25, 181) <= 1; play_W(25, 182) <= 1; play_W(25, 183) <= 0; play_W(25, 184) <= 0; play_W(25, 185) <= 0; play_W(25, 186) <= 0; play_W(25, 187) <= 0; play_W(25, 188) <= 0; play_W(25, 189) <= 0; play_W(25, 190) <= 0; play_W(25, 191) <= 0; play_W(25, 192) <= 0; play_W(25, 193) <= 0; play_W(25, 194) <= 0; play_W(25, 195) <= 0; play_W(25, 196) <= 0; play_W(25, 197) <= 0; play_W(25, 198) <= 1; play_W(25, 199) <= 1; play_W(25, 200) <= 1; play_W(25, 201) <= 1; play_W(25, 202) <= 1; play_W(25, 203) <= 1; play_W(25, 204) <= 0; play_W(25, 205) <= 0; play_W(25, 206) <= 0; play_W(25, 207) <= 0; play_W(25, 208) <= 0; play_W(25, 209) <= 0; play_W(25, 210) <= 0; play_W(25, 211) <= 0; play_W(25, 212) <= 0; play_W(25, 213) <= 0; play_W(25, 214) <= 0; play_W(25, 215) <= 0; play_W(25, 216) <= 1; play_W(25, 217) <= 1; play_W(25, 218) <= 1; play_W(25, 219) <= 1; play_W(25, 220) <= 1; play_W(25, 221) <= 1; play_W(25, 222) <= 0; play_W(25, 223) <= 0; play_W(25, 224) <= 0; play_W(25, 225) <= 0; play_W(25, 226) <= 0; play_W(25, 227) <= 0; play_W(25, 228) <= 0; play_W(25, 229) <= 0; play_W(25, 230) <= 0; play_W(25, 231) <= 1; play_W(25, 232) <= 1; play_W(25, 233) <= 1; play_W(25, 234) <= 1; play_W(25, 235) <= 1; play_W(25, 236) <= 1; play_W(25, 237) <= 0; play_W(25, 238) <= 0; play_W(25, 239) <= 0; play_W(25, 240) <= 0; play_W(25, 241) <= 0; play_W(25, 242) <= 0; play_W(25, 243) <= 0; play_W(25, 244) <= 0; play_W(25, 245) <= 0; play_W(25, 246) <= 1; play_W(25, 247) <= 1; play_W(25, 248) <= 1; play_W(25, 249) <= 1; play_W(25, 250) <= 1; play_W(25, 251) <= 1; play_W(25, 252) <= 0; play_W(25, 253) <= 0; play_W(25, 254) <= 0; play_W(25, 255) <= 0; play_W(25, 256) <= 0; play_W(25, 257) <= 0; play_W(25, 258) <= 1; play_W(25, 259) <= 1; play_W(25, 260) <= 1; play_W(25, 261) <= 1; play_W(25, 262) <= 1; play_W(25, 263) <= 1; play_W(25, 264) <= 0; play_W(25, 265) <= 0; play_W(25, 266) <= 0; play_W(25, 267) <= 0; play_W(25, 268) <= 0; play_W(25, 269) <= 0; 
play_W(26, 0) <= 0; play_W(26, 1) <= 0; play_W(26, 2) <= 0; play_W(26, 3) <= 1; play_W(26, 4) <= 1; play_W(26, 5) <= 1; play_W(26, 6) <= 1; play_W(26, 7) <= 1; play_W(26, 8) <= 1; play_W(26, 9) <= 0; play_W(26, 10) <= 0; play_W(26, 11) <= 0; play_W(26, 12) <= 0; play_W(26, 13) <= 0; play_W(26, 14) <= 0; play_W(26, 15) <= 0; play_W(26, 16) <= 0; play_W(26, 17) <= 0; play_W(26, 18) <= 0; play_W(26, 19) <= 0; play_W(26, 20) <= 0; play_W(26, 21) <= 0; play_W(26, 22) <= 0; play_W(26, 23) <= 0; play_W(26, 24) <= 0; play_W(26, 25) <= 0; play_W(26, 26) <= 0; play_W(26, 27) <= 0; play_W(26, 28) <= 0; play_W(26, 29) <= 0; play_W(26, 30) <= 1; play_W(26, 31) <= 1; play_W(26, 32) <= 1; play_W(26, 33) <= 1; play_W(26, 34) <= 1; play_W(26, 35) <= 1; play_W(26, 36) <= 0; play_W(26, 37) <= 0; play_W(26, 38) <= 0; play_W(26, 39) <= 0; play_W(26, 40) <= 0; play_W(26, 41) <= 0; play_W(26, 42) <= 1; play_W(26, 43) <= 1; play_W(26, 44) <= 1; play_W(26, 45) <= 1; play_W(26, 46) <= 1; play_W(26, 47) <= 1; play_W(26, 48) <= 0; play_W(26, 49) <= 0; play_W(26, 50) <= 0; play_W(26, 51) <= 0; play_W(26, 52) <= 0; play_W(26, 53) <= 0; play_W(26, 54) <= 1; play_W(26, 55) <= 1; play_W(26, 56) <= 1; play_W(26, 57) <= 1; play_W(26, 58) <= 1; play_W(26, 59) <= 1; play_W(26, 60) <= 0; play_W(26, 61) <= 0; play_W(26, 62) <= 0; play_W(26, 63) <= 0; play_W(26, 64) <= 0; play_W(26, 65) <= 0; play_W(26, 66) <= 0; play_W(26, 67) <= 0; play_W(26, 68) <= 0; play_W(26, 69) <= 1; play_W(26, 70) <= 1; play_W(26, 71) <= 1; play_W(26, 72) <= 1; play_W(26, 73) <= 1; play_W(26, 74) <= 1; play_W(26, 75) <= 0; play_W(26, 76) <= 0; play_W(26, 77) <= 0; play_W(26, 78) <= 0; play_W(26, 79) <= 0; play_W(26, 80) <= 0; play_W(26, 81) <= 0; play_W(26, 82) <= 0; play_W(26, 83) <= 0; play_W(26, 84) <= 0; play_W(26, 85) <= 0; play_W(26, 86) <= 0; play_W(26, 87) <= 0; play_W(26, 88) <= 0; play_W(26, 89) <= 0; play_W(26, 90) <= 1; play_W(26, 91) <= 1; play_W(26, 92) <= 1; play_W(26, 93) <= 1; play_W(26, 94) <= 1; play_W(26, 95) <= 1; play_W(26, 96) <= 0; play_W(26, 97) <= 0; play_W(26, 98) <= 0; play_W(26, 99) <= 0; play_W(26, 100) <= 0; play_W(26, 101) <= 0; play_W(26, 102) <= 0; play_W(26, 103) <= 0; play_W(26, 104) <= 0; play_W(26, 105) <= 0; play_W(26, 106) <= 0; play_W(26, 107) <= 0; play_W(26, 108) <= 0; play_W(26, 109) <= 0; play_W(26, 110) <= 0; play_W(26, 111) <= 0; play_W(26, 112) <= 0; play_W(26, 113) <= 0; play_W(26, 114) <= 0; play_W(26, 115) <= 0; play_W(26, 116) <= 0; play_W(26, 117) <= 0; play_W(26, 118) <= 0; play_W(26, 119) <= 0; play_W(26, 120) <= 0; play_W(26, 121) <= 0; play_W(26, 122) <= 0; play_W(26, 123) <= 0; play_W(26, 124) <= 0; play_W(26, 125) <= 0; play_W(26, 126) <= 0; play_W(26, 127) <= 0; play_W(26, 128) <= 0; play_W(26, 129) <= 0; play_W(26, 130) <= 0; play_W(26, 131) <= 0; play_W(26, 132) <= 0; play_W(26, 133) <= 0; play_W(26, 134) <= 0; play_W(26, 135) <= 0; play_W(26, 136) <= 0; play_W(26, 137) <= 0; play_W(26, 138) <= 0; play_W(26, 139) <= 0; play_W(26, 140) <= 0; play_W(26, 141) <= 0; play_W(26, 142) <= 0; play_W(26, 143) <= 0; play_W(26, 144) <= 0; play_W(26, 145) <= 0; play_W(26, 146) <= 0; play_W(26, 147) <= 0; play_W(26, 148) <= 0; play_W(26, 149) <= 0; play_W(26, 150) <= 0; play_W(26, 151) <= 0; play_W(26, 152) <= 0; play_W(26, 153) <= 0; play_W(26, 154) <= 0; play_W(26, 155) <= 0; play_W(26, 156) <= 0; play_W(26, 157) <= 0; play_W(26, 158) <= 0; play_W(26, 159) <= 0; play_W(26, 160) <= 0; play_W(26, 161) <= 0; play_W(26, 162) <= 0; play_W(26, 163) <= 0; play_W(26, 164) <= 0; play_W(26, 165) <= 1; play_W(26, 166) <= 1; play_W(26, 167) <= 1; play_W(26, 168) <= 1; play_W(26, 169) <= 1; play_W(26, 170) <= 1; play_W(26, 171) <= 0; play_W(26, 172) <= 0; play_W(26, 173) <= 0; play_W(26, 174) <= 0; play_W(26, 175) <= 0; play_W(26, 176) <= 0; play_W(26, 177) <= 1; play_W(26, 178) <= 1; play_W(26, 179) <= 1; play_W(26, 180) <= 1; play_W(26, 181) <= 1; play_W(26, 182) <= 1; play_W(26, 183) <= 0; play_W(26, 184) <= 0; play_W(26, 185) <= 0; play_W(26, 186) <= 0; play_W(26, 187) <= 0; play_W(26, 188) <= 0; play_W(26, 189) <= 0; play_W(26, 190) <= 0; play_W(26, 191) <= 0; play_W(26, 192) <= 0; play_W(26, 193) <= 0; play_W(26, 194) <= 0; play_W(26, 195) <= 0; play_W(26, 196) <= 0; play_W(26, 197) <= 0; play_W(26, 198) <= 1; play_W(26, 199) <= 1; play_W(26, 200) <= 1; play_W(26, 201) <= 1; play_W(26, 202) <= 1; play_W(26, 203) <= 1; play_W(26, 204) <= 0; play_W(26, 205) <= 0; play_W(26, 206) <= 0; play_W(26, 207) <= 0; play_W(26, 208) <= 0; play_W(26, 209) <= 0; play_W(26, 210) <= 0; play_W(26, 211) <= 0; play_W(26, 212) <= 0; play_W(26, 213) <= 0; play_W(26, 214) <= 0; play_W(26, 215) <= 0; play_W(26, 216) <= 1; play_W(26, 217) <= 1; play_W(26, 218) <= 1; play_W(26, 219) <= 1; play_W(26, 220) <= 1; play_W(26, 221) <= 1; play_W(26, 222) <= 0; play_W(26, 223) <= 0; play_W(26, 224) <= 0; play_W(26, 225) <= 0; play_W(26, 226) <= 0; play_W(26, 227) <= 0; play_W(26, 228) <= 0; play_W(26, 229) <= 0; play_W(26, 230) <= 0; play_W(26, 231) <= 1; play_W(26, 232) <= 1; play_W(26, 233) <= 1; play_W(26, 234) <= 1; play_W(26, 235) <= 1; play_W(26, 236) <= 1; play_W(26, 237) <= 0; play_W(26, 238) <= 0; play_W(26, 239) <= 0; play_W(26, 240) <= 0; play_W(26, 241) <= 0; play_W(26, 242) <= 0; play_W(26, 243) <= 0; play_W(26, 244) <= 0; play_W(26, 245) <= 0; play_W(26, 246) <= 1; play_W(26, 247) <= 1; play_W(26, 248) <= 1; play_W(26, 249) <= 1; play_W(26, 250) <= 1; play_W(26, 251) <= 1; play_W(26, 252) <= 0; play_W(26, 253) <= 0; play_W(26, 254) <= 0; play_W(26, 255) <= 0; play_W(26, 256) <= 0; play_W(26, 257) <= 0; play_W(26, 258) <= 1; play_W(26, 259) <= 1; play_W(26, 260) <= 1; play_W(26, 261) <= 1; play_W(26, 262) <= 1; play_W(26, 263) <= 1; play_W(26, 264) <= 0; play_W(26, 265) <= 0; play_W(26, 266) <= 0; play_W(26, 267) <= 0; play_W(26, 268) <= 0; play_W(26, 269) <= 0; 
play_W(27, 0) <= 1; play_W(27, 1) <= 1; play_W(27, 2) <= 1; play_W(27, 3) <= 1; play_W(27, 4) <= 1; play_W(27, 5) <= 1; play_W(27, 6) <= 1; play_W(27, 7) <= 1; play_W(27, 8) <= 1; play_W(27, 9) <= 1; play_W(27, 10) <= 1; play_W(27, 11) <= 1; play_W(27, 12) <= 0; play_W(27, 13) <= 0; play_W(27, 14) <= 0; play_W(27, 15) <= 0; play_W(27, 16) <= 0; play_W(27, 17) <= 0; play_W(27, 18) <= 0; play_W(27, 19) <= 0; play_W(27, 20) <= 0; play_W(27, 21) <= 0; play_W(27, 22) <= 0; play_W(27, 23) <= 0; play_W(27, 24) <= 0; play_W(27, 25) <= 0; play_W(27, 26) <= 0; play_W(27, 27) <= 1; play_W(27, 28) <= 1; play_W(27, 29) <= 1; play_W(27, 30) <= 1; play_W(27, 31) <= 1; play_W(27, 32) <= 1; play_W(27, 33) <= 1; play_W(27, 34) <= 1; play_W(27, 35) <= 1; play_W(27, 36) <= 1; play_W(27, 37) <= 1; play_W(27, 38) <= 1; play_W(27, 39) <= 1; play_W(27, 40) <= 1; play_W(27, 41) <= 1; play_W(27, 42) <= 1; play_W(27, 43) <= 1; play_W(27, 44) <= 1; play_W(27, 45) <= 1; play_W(27, 46) <= 1; play_W(27, 47) <= 1; play_W(27, 48) <= 0; play_W(27, 49) <= 0; play_W(27, 50) <= 0; play_W(27, 51) <= 0; play_W(27, 52) <= 0; play_W(27, 53) <= 0; play_W(27, 54) <= 1; play_W(27, 55) <= 1; play_W(27, 56) <= 1; play_W(27, 57) <= 1; play_W(27, 58) <= 1; play_W(27, 59) <= 1; play_W(27, 60) <= 0; play_W(27, 61) <= 0; play_W(27, 62) <= 0; play_W(27, 63) <= 0; play_W(27, 64) <= 0; play_W(27, 65) <= 0; play_W(27, 66) <= 0; play_W(27, 67) <= 0; play_W(27, 68) <= 0; play_W(27, 69) <= 1; play_W(27, 70) <= 1; play_W(27, 71) <= 1; play_W(27, 72) <= 1; play_W(27, 73) <= 1; play_W(27, 74) <= 1; play_W(27, 75) <= 0; play_W(27, 76) <= 0; play_W(27, 77) <= 0; play_W(27, 78) <= 0; play_W(27, 79) <= 0; play_W(27, 80) <= 0; play_W(27, 81) <= 0; play_W(27, 82) <= 0; play_W(27, 83) <= 0; play_W(27, 84) <= 0; play_W(27, 85) <= 0; play_W(27, 86) <= 0; play_W(27, 87) <= 1; play_W(27, 88) <= 1; play_W(27, 89) <= 1; play_W(27, 90) <= 1; play_W(27, 91) <= 1; play_W(27, 92) <= 1; play_W(27, 93) <= 1; play_W(27, 94) <= 1; play_W(27, 95) <= 1; play_W(27, 96) <= 1; play_W(27, 97) <= 1; play_W(27, 98) <= 1; play_W(27, 99) <= 0; play_W(27, 100) <= 0; play_W(27, 101) <= 0; play_W(27, 102) <= 0; play_W(27, 103) <= 0; play_W(27, 104) <= 0; play_W(27, 105) <= 0; play_W(27, 106) <= 0; play_W(27, 107) <= 0; play_W(27, 108) <= 0; play_W(27, 109) <= 0; play_W(27, 110) <= 0; play_W(27, 111) <= 0; play_W(27, 112) <= 0; play_W(27, 113) <= 0; play_W(27, 114) <= 0; play_W(27, 115) <= 0; play_W(27, 116) <= 0; play_W(27, 117) <= 0; play_W(27, 118) <= 0; play_W(27, 119) <= 0; play_W(27, 120) <= 0; play_W(27, 121) <= 0; play_W(27, 122) <= 0; play_W(27, 123) <= 0; play_W(27, 124) <= 0; play_W(27, 125) <= 0; play_W(27, 126) <= 0; play_W(27, 127) <= 0; play_W(27, 128) <= 0; play_W(27, 129) <= 0; play_W(27, 130) <= 0; play_W(27, 131) <= 0; play_W(27, 132) <= 0; play_W(27, 133) <= 0; play_W(27, 134) <= 0; play_W(27, 135) <= 0; play_W(27, 136) <= 0; play_W(27, 137) <= 0; play_W(27, 138) <= 0; play_W(27, 139) <= 0; play_W(27, 140) <= 0; play_W(27, 141) <= 0; play_W(27, 142) <= 0; play_W(27, 143) <= 0; play_W(27, 144) <= 0; play_W(27, 145) <= 0; play_W(27, 146) <= 0; play_W(27, 147) <= 0; play_W(27, 148) <= 0; play_W(27, 149) <= 0; play_W(27, 150) <= 0; play_W(27, 151) <= 0; play_W(27, 152) <= 0; play_W(27, 153) <= 0; play_W(27, 154) <= 0; play_W(27, 155) <= 0; play_W(27, 156) <= 0; play_W(27, 157) <= 0; play_W(27, 158) <= 0; play_W(27, 159) <= 0; play_W(27, 160) <= 0; play_W(27, 161) <= 0; play_W(27, 162) <= 1; play_W(27, 163) <= 1; play_W(27, 164) <= 1; play_W(27, 165) <= 1; play_W(27, 166) <= 1; play_W(27, 167) <= 1; play_W(27, 168) <= 1; play_W(27, 169) <= 1; play_W(27, 170) <= 1; play_W(27, 171) <= 1; play_W(27, 172) <= 1; play_W(27, 173) <= 1; play_W(27, 174) <= 1; play_W(27, 175) <= 1; play_W(27, 176) <= 1; play_W(27, 177) <= 1; play_W(27, 178) <= 1; play_W(27, 179) <= 1; play_W(27, 180) <= 0; play_W(27, 181) <= 0; play_W(27, 182) <= 0; play_W(27, 183) <= 0; play_W(27, 184) <= 0; play_W(27, 185) <= 0; play_W(27, 186) <= 0; play_W(27, 187) <= 0; play_W(27, 188) <= 0; play_W(27, 189) <= 0; play_W(27, 190) <= 0; play_W(27, 191) <= 0; play_W(27, 192) <= 0; play_W(27, 193) <= 0; play_W(27, 194) <= 0; play_W(27, 195) <= 1; play_W(27, 196) <= 1; play_W(27, 197) <= 1; play_W(27, 198) <= 1; play_W(27, 199) <= 1; play_W(27, 200) <= 1; play_W(27, 201) <= 1; play_W(27, 202) <= 1; play_W(27, 203) <= 1; play_W(27, 204) <= 1; play_W(27, 205) <= 1; play_W(27, 206) <= 1; play_W(27, 207) <= 0; play_W(27, 208) <= 0; play_W(27, 209) <= 0; play_W(27, 210) <= 0; play_W(27, 211) <= 0; play_W(27, 212) <= 0; play_W(27, 213) <= 0; play_W(27, 214) <= 0; play_W(27, 215) <= 0; play_W(27, 216) <= 1; play_W(27, 217) <= 1; play_W(27, 218) <= 1; play_W(27, 219) <= 1; play_W(27, 220) <= 1; play_W(27, 221) <= 1; play_W(27, 222) <= 0; play_W(27, 223) <= 0; play_W(27, 224) <= 0; play_W(27, 225) <= 0; play_W(27, 226) <= 0; play_W(27, 227) <= 0; play_W(27, 228) <= 0; play_W(27, 229) <= 0; play_W(27, 230) <= 0; play_W(27, 231) <= 1; play_W(27, 232) <= 1; play_W(27, 233) <= 1; play_W(27, 234) <= 1; play_W(27, 235) <= 1; play_W(27, 236) <= 1; play_W(27, 237) <= 0; play_W(27, 238) <= 0; play_W(27, 239) <= 0; play_W(27, 240) <= 0; play_W(27, 241) <= 0; play_W(27, 242) <= 0; play_W(27, 243) <= 1; play_W(27, 244) <= 1; play_W(27, 245) <= 1; play_W(27, 246) <= 1; play_W(27, 247) <= 1; play_W(27, 248) <= 1; play_W(27, 249) <= 1; play_W(27, 250) <= 1; play_W(27, 251) <= 1; play_W(27, 252) <= 0; play_W(27, 253) <= 0; play_W(27, 254) <= 0; play_W(27, 255) <= 0; play_W(27, 256) <= 0; play_W(27, 257) <= 0; play_W(27, 258) <= 1; play_W(27, 259) <= 1; play_W(27, 260) <= 1; play_W(27, 261) <= 1; play_W(27, 262) <= 1; play_W(27, 263) <= 1; play_W(27, 264) <= 0; play_W(27, 265) <= 0; play_W(27, 266) <= 0; play_W(27, 267) <= 0; play_W(27, 268) <= 0; play_W(27, 269) <= 0; 
play_W(28, 0) <= 1; play_W(28, 1) <= 1; play_W(28, 2) <= 1; play_W(28, 3) <= 1; play_W(28, 4) <= 1; play_W(28, 5) <= 1; play_W(28, 6) <= 1; play_W(28, 7) <= 1; play_W(28, 8) <= 1; play_W(28, 9) <= 1; play_W(28, 10) <= 1; play_W(28, 11) <= 1; play_W(28, 12) <= 0; play_W(28, 13) <= 0; play_W(28, 14) <= 0; play_W(28, 15) <= 0; play_W(28, 16) <= 0; play_W(28, 17) <= 0; play_W(28, 18) <= 0; play_W(28, 19) <= 0; play_W(28, 20) <= 0; play_W(28, 21) <= 0; play_W(28, 22) <= 0; play_W(28, 23) <= 0; play_W(28, 24) <= 0; play_W(28, 25) <= 0; play_W(28, 26) <= 0; play_W(28, 27) <= 1; play_W(28, 28) <= 1; play_W(28, 29) <= 1; play_W(28, 30) <= 1; play_W(28, 31) <= 1; play_W(28, 32) <= 1; play_W(28, 33) <= 1; play_W(28, 34) <= 1; play_W(28, 35) <= 1; play_W(28, 36) <= 1; play_W(28, 37) <= 1; play_W(28, 38) <= 1; play_W(28, 39) <= 1; play_W(28, 40) <= 1; play_W(28, 41) <= 1; play_W(28, 42) <= 1; play_W(28, 43) <= 1; play_W(28, 44) <= 1; play_W(28, 45) <= 1; play_W(28, 46) <= 1; play_W(28, 47) <= 1; play_W(28, 48) <= 0; play_W(28, 49) <= 0; play_W(28, 50) <= 0; play_W(28, 51) <= 0; play_W(28, 52) <= 0; play_W(28, 53) <= 0; play_W(28, 54) <= 1; play_W(28, 55) <= 1; play_W(28, 56) <= 1; play_W(28, 57) <= 1; play_W(28, 58) <= 1; play_W(28, 59) <= 1; play_W(28, 60) <= 0; play_W(28, 61) <= 0; play_W(28, 62) <= 0; play_W(28, 63) <= 0; play_W(28, 64) <= 0; play_W(28, 65) <= 0; play_W(28, 66) <= 0; play_W(28, 67) <= 0; play_W(28, 68) <= 0; play_W(28, 69) <= 1; play_W(28, 70) <= 1; play_W(28, 71) <= 1; play_W(28, 72) <= 1; play_W(28, 73) <= 1; play_W(28, 74) <= 1; play_W(28, 75) <= 0; play_W(28, 76) <= 0; play_W(28, 77) <= 0; play_W(28, 78) <= 0; play_W(28, 79) <= 0; play_W(28, 80) <= 0; play_W(28, 81) <= 0; play_W(28, 82) <= 0; play_W(28, 83) <= 0; play_W(28, 84) <= 0; play_W(28, 85) <= 0; play_W(28, 86) <= 0; play_W(28, 87) <= 1; play_W(28, 88) <= 1; play_W(28, 89) <= 1; play_W(28, 90) <= 1; play_W(28, 91) <= 1; play_W(28, 92) <= 1; play_W(28, 93) <= 1; play_W(28, 94) <= 1; play_W(28, 95) <= 1; play_W(28, 96) <= 1; play_W(28, 97) <= 1; play_W(28, 98) <= 1; play_W(28, 99) <= 0; play_W(28, 100) <= 0; play_W(28, 101) <= 0; play_W(28, 102) <= 0; play_W(28, 103) <= 0; play_W(28, 104) <= 0; play_W(28, 105) <= 0; play_W(28, 106) <= 0; play_W(28, 107) <= 0; play_W(28, 108) <= 0; play_W(28, 109) <= 0; play_W(28, 110) <= 0; play_W(28, 111) <= 0; play_W(28, 112) <= 0; play_W(28, 113) <= 0; play_W(28, 114) <= 0; play_W(28, 115) <= 0; play_W(28, 116) <= 0; play_W(28, 117) <= 0; play_W(28, 118) <= 0; play_W(28, 119) <= 0; play_W(28, 120) <= 0; play_W(28, 121) <= 0; play_W(28, 122) <= 0; play_W(28, 123) <= 0; play_W(28, 124) <= 0; play_W(28, 125) <= 0; play_W(28, 126) <= 0; play_W(28, 127) <= 0; play_W(28, 128) <= 0; play_W(28, 129) <= 0; play_W(28, 130) <= 0; play_W(28, 131) <= 0; play_W(28, 132) <= 0; play_W(28, 133) <= 0; play_W(28, 134) <= 0; play_W(28, 135) <= 0; play_W(28, 136) <= 0; play_W(28, 137) <= 0; play_W(28, 138) <= 0; play_W(28, 139) <= 0; play_W(28, 140) <= 0; play_W(28, 141) <= 0; play_W(28, 142) <= 0; play_W(28, 143) <= 0; play_W(28, 144) <= 0; play_W(28, 145) <= 0; play_W(28, 146) <= 0; play_W(28, 147) <= 0; play_W(28, 148) <= 0; play_W(28, 149) <= 0; play_W(28, 150) <= 0; play_W(28, 151) <= 0; play_W(28, 152) <= 0; play_W(28, 153) <= 0; play_W(28, 154) <= 0; play_W(28, 155) <= 0; play_W(28, 156) <= 0; play_W(28, 157) <= 0; play_W(28, 158) <= 0; play_W(28, 159) <= 0; play_W(28, 160) <= 0; play_W(28, 161) <= 0; play_W(28, 162) <= 1; play_W(28, 163) <= 1; play_W(28, 164) <= 1; play_W(28, 165) <= 1; play_W(28, 166) <= 1; play_W(28, 167) <= 1; play_W(28, 168) <= 1; play_W(28, 169) <= 1; play_W(28, 170) <= 1; play_W(28, 171) <= 1; play_W(28, 172) <= 1; play_W(28, 173) <= 1; play_W(28, 174) <= 1; play_W(28, 175) <= 1; play_W(28, 176) <= 1; play_W(28, 177) <= 1; play_W(28, 178) <= 1; play_W(28, 179) <= 1; play_W(28, 180) <= 0; play_W(28, 181) <= 0; play_W(28, 182) <= 0; play_W(28, 183) <= 0; play_W(28, 184) <= 0; play_W(28, 185) <= 0; play_W(28, 186) <= 0; play_W(28, 187) <= 0; play_W(28, 188) <= 0; play_W(28, 189) <= 0; play_W(28, 190) <= 0; play_W(28, 191) <= 0; play_W(28, 192) <= 0; play_W(28, 193) <= 0; play_W(28, 194) <= 0; play_W(28, 195) <= 1; play_W(28, 196) <= 1; play_W(28, 197) <= 1; play_W(28, 198) <= 1; play_W(28, 199) <= 1; play_W(28, 200) <= 1; play_W(28, 201) <= 1; play_W(28, 202) <= 1; play_W(28, 203) <= 1; play_W(28, 204) <= 1; play_W(28, 205) <= 1; play_W(28, 206) <= 1; play_W(28, 207) <= 0; play_W(28, 208) <= 0; play_W(28, 209) <= 0; play_W(28, 210) <= 0; play_W(28, 211) <= 0; play_W(28, 212) <= 0; play_W(28, 213) <= 0; play_W(28, 214) <= 0; play_W(28, 215) <= 0; play_W(28, 216) <= 1; play_W(28, 217) <= 1; play_W(28, 218) <= 1; play_W(28, 219) <= 1; play_W(28, 220) <= 1; play_W(28, 221) <= 1; play_W(28, 222) <= 0; play_W(28, 223) <= 0; play_W(28, 224) <= 0; play_W(28, 225) <= 0; play_W(28, 226) <= 0; play_W(28, 227) <= 0; play_W(28, 228) <= 0; play_W(28, 229) <= 0; play_W(28, 230) <= 0; play_W(28, 231) <= 1; play_W(28, 232) <= 1; play_W(28, 233) <= 1; play_W(28, 234) <= 1; play_W(28, 235) <= 1; play_W(28, 236) <= 1; play_W(28, 237) <= 0; play_W(28, 238) <= 0; play_W(28, 239) <= 0; play_W(28, 240) <= 0; play_W(28, 241) <= 0; play_W(28, 242) <= 0; play_W(28, 243) <= 1; play_W(28, 244) <= 1; play_W(28, 245) <= 1; play_W(28, 246) <= 1; play_W(28, 247) <= 1; play_W(28, 248) <= 1; play_W(28, 249) <= 1; play_W(28, 250) <= 1; play_W(28, 251) <= 1; play_W(28, 252) <= 0; play_W(28, 253) <= 0; play_W(28, 254) <= 0; play_W(28, 255) <= 0; play_W(28, 256) <= 0; play_W(28, 257) <= 0; play_W(28, 258) <= 1; play_W(28, 259) <= 1; play_W(28, 260) <= 1; play_W(28, 261) <= 1; play_W(28, 262) <= 1; play_W(28, 263) <= 1; play_W(28, 264) <= 0; play_W(28, 265) <= 0; play_W(28, 266) <= 0; play_W(28, 267) <= 0; play_W(28, 268) <= 0; play_W(28, 269) <= 0; 
play_W(29, 0) <= 1; play_W(29, 1) <= 1; play_W(29, 2) <= 1; play_W(29, 3) <= 1; play_W(29, 4) <= 1; play_W(29, 5) <= 1; play_W(29, 6) <= 1; play_W(29, 7) <= 1; play_W(29, 8) <= 1; play_W(29, 9) <= 1; play_W(29, 10) <= 1; play_W(29, 11) <= 1; play_W(29, 12) <= 0; play_W(29, 13) <= 0; play_W(29, 14) <= 0; play_W(29, 15) <= 0; play_W(29, 16) <= 0; play_W(29, 17) <= 0; play_W(29, 18) <= 0; play_W(29, 19) <= 0; play_W(29, 20) <= 0; play_W(29, 21) <= 0; play_W(29, 22) <= 0; play_W(29, 23) <= 0; play_W(29, 24) <= 0; play_W(29, 25) <= 0; play_W(29, 26) <= 0; play_W(29, 27) <= 1; play_W(29, 28) <= 1; play_W(29, 29) <= 1; play_W(29, 30) <= 1; play_W(29, 31) <= 1; play_W(29, 32) <= 1; play_W(29, 33) <= 1; play_W(29, 34) <= 1; play_W(29, 35) <= 1; play_W(29, 36) <= 1; play_W(29, 37) <= 1; play_W(29, 38) <= 1; play_W(29, 39) <= 1; play_W(29, 40) <= 1; play_W(29, 41) <= 1; play_W(29, 42) <= 1; play_W(29, 43) <= 1; play_W(29, 44) <= 1; play_W(29, 45) <= 1; play_W(29, 46) <= 1; play_W(29, 47) <= 1; play_W(29, 48) <= 0; play_W(29, 49) <= 0; play_W(29, 50) <= 0; play_W(29, 51) <= 0; play_W(29, 52) <= 0; play_W(29, 53) <= 0; play_W(29, 54) <= 1; play_W(29, 55) <= 1; play_W(29, 56) <= 1; play_W(29, 57) <= 1; play_W(29, 58) <= 1; play_W(29, 59) <= 1; play_W(29, 60) <= 0; play_W(29, 61) <= 0; play_W(29, 62) <= 0; play_W(29, 63) <= 0; play_W(29, 64) <= 0; play_W(29, 65) <= 0; play_W(29, 66) <= 0; play_W(29, 67) <= 0; play_W(29, 68) <= 0; play_W(29, 69) <= 1; play_W(29, 70) <= 1; play_W(29, 71) <= 1; play_W(29, 72) <= 1; play_W(29, 73) <= 1; play_W(29, 74) <= 1; play_W(29, 75) <= 0; play_W(29, 76) <= 0; play_W(29, 77) <= 0; play_W(29, 78) <= 0; play_W(29, 79) <= 0; play_W(29, 80) <= 0; play_W(29, 81) <= 0; play_W(29, 82) <= 0; play_W(29, 83) <= 0; play_W(29, 84) <= 0; play_W(29, 85) <= 0; play_W(29, 86) <= 0; play_W(29, 87) <= 1; play_W(29, 88) <= 1; play_W(29, 89) <= 1; play_W(29, 90) <= 1; play_W(29, 91) <= 1; play_W(29, 92) <= 1; play_W(29, 93) <= 1; play_W(29, 94) <= 1; play_W(29, 95) <= 1; play_W(29, 96) <= 1; play_W(29, 97) <= 1; play_W(29, 98) <= 1; play_W(29, 99) <= 0; play_W(29, 100) <= 0; play_W(29, 101) <= 0; play_W(29, 102) <= 0; play_W(29, 103) <= 0; play_W(29, 104) <= 0; play_W(29, 105) <= 0; play_W(29, 106) <= 0; play_W(29, 107) <= 0; play_W(29, 108) <= 0; play_W(29, 109) <= 0; play_W(29, 110) <= 0; play_W(29, 111) <= 0; play_W(29, 112) <= 0; play_W(29, 113) <= 0; play_W(29, 114) <= 0; play_W(29, 115) <= 0; play_W(29, 116) <= 0; play_W(29, 117) <= 0; play_W(29, 118) <= 0; play_W(29, 119) <= 0; play_W(29, 120) <= 0; play_W(29, 121) <= 0; play_W(29, 122) <= 0; play_W(29, 123) <= 0; play_W(29, 124) <= 0; play_W(29, 125) <= 0; play_W(29, 126) <= 0; play_W(29, 127) <= 0; play_W(29, 128) <= 0; play_W(29, 129) <= 0; play_W(29, 130) <= 0; play_W(29, 131) <= 0; play_W(29, 132) <= 0; play_W(29, 133) <= 0; play_W(29, 134) <= 0; play_W(29, 135) <= 0; play_W(29, 136) <= 0; play_W(29, 137) <= 0; play_W(29, 138) <= 0; play_W(29, 139) <= 0; play_W(29, 140) <= 0; play_W(29, 141) <= 0; play_W(29, 142) <= 0; play_W(29, 143) <= 0; play_W(29, 144) <= 0; play_W(29, 145) <= 0; play_W(29, 146) <= 0; play_W(29, 147) <= 0; play_W(29, 148) <= 0; play_W(29, 149) <= 0; play_W(29, 150) <= 0; play_W(29, 151) <= 0; play_W(29, 152) <= 0; play_W(29, 153) <= 0; play_W(29, 154) <= 0; play_W(29, 155) <= 0; play_W(29, 156) <= 0; play_W(29, 157) <= 0; play_W(29, 158) <= 0; play_W(29, 159) <= 0; play_W(29, 160) <= 0; play_W(29, 161) <= 0; play_W(29, 162) <= 1; play_W(29, 163) <= 1; play_W(29, 164) <= 1; play_W(29, 165) <= 1; play_W(29, 166) <= 1; play_W(29, 167) <= 1; play_W(29, 168) <= 1; play_W(29, 169) <= 1; play_W(29, 170) <= 1; play_W(29, 171) <= 1; play_W(29, 172) <= 1; play_W(29, 173) <= 1; play_W(29, 174) <= 1; play_W(29, 175) <= 1; play_W(29, 176) <= 1; play_W(29, 177) <= 1; play_W(29, 178) <= 1; play_W(29, 179) <= 1; play_W(29, 180) <= 0; play_W(29, 181) <= 0; play_W(29, 182) <= 0; play_W(29, 183) <= 0; play_W(29, 184) <= 0; play_W(29, 185) <= 0; play_W(29, 186) <= 0; play_W(29, 187) <= 0; play_W(29, 188) <= 0; play_W(29, 189) <= 0; play_W(29, 190) <= 0; play_W(29, 191) <= 0; play_W(29, 192) <= 0; play_W(29, 193) <= 0; play_W(29, 194) <= 0; play_W(29, 195) <= 1; play_W(29, 196) <= 1; play_W(29, 197) <= 1; play_W(29, 198) <= 1; play_W(29, 199) <= 1; play_W(29, 200) <= 1; play_W(29, 201) <= 1; play_W(29, 202) <= 1; play_W(29, 203) <= 1; play_W(29, 204) <= 1; play_W(29, 205) <= 1; play_W(29, 206) <= 1; play_W(29, 207) <= 0; play_W(29, 208) <= 0; play_W(29, 209) <= 0; play_W(29, 210) <= 0; play_W(29, 211) <= 0; play_W(29, 212) <= 0; play_W(29, 213) <= 0; play_W(29, 214) <= 0; play_W(29, 215) <= 0; play_W(29, 216) <= 1; play_W(29, 217) <= 1; play_W(29, 218) <= 1; play_W(29, 219) <= 1; play_W(29, 220) <= 1; play_W(29, 221) <= 1; play_W(29, 222) <= 0; play_W(29, 223) <= 0; play_W(29, 224) <= 0; play_W(29, 225) <= 0; play_W(29, 226) <= 0; play_W(29, 227) <= 0; play_W(29, 228) <= 0; play_W(29, 229) <= 0; play_W(29, 230) <= 0; play_W(29, 231) <= 1; play_W(29, 232) <= 1; play_W(29, 233) <= 1; play_W(29, 234) <= 1; play_W(29, 235) <= 1; play_W(29, 236) <= 1; play_W(29, 237) <= 0; play_W(29, 238) <= 0; play_W(29, 239) <= 0; play_W(29, 240) <= 0; play_W(29, 241) <= 0; play_W(29, 242) <= 0; play_W(29, 243) <= 1; play_W(29, 244) <= 1; play_W(29, 245) <= 1; play_W(29, 246) <= 1; play_W(29, 247) <= 1; play_W(29, 248) <= 1; play_W(29, 249) <= 1; play_W(29, 250) <= 1; play_W(29, 251) <= 1; play_W(29, 252) <= 0; play_W(29, 253) <= 0; play_W(29, 254) <= 0; play_W(29, 255) <= 0; play_W(29, 256) <= 0; play_W(29, 257) <= 0; play_W(29, 258) <= 1; play_W(29, 259) <= 1; play_W(29, 260) <= 1; play_W(29, 261) <= 1; play_W(29, 262) <= 1; play_W(29, 263) <= 1; play_W(29, 264) <= 0; play_W(29, 265) <= 0; play_W(29, 266) <= 0; play_W(29, 267) <= 0; play_W(29, 268) <= 0; play_W(29, 269) <= 0; 
end Behavioral;
